magic
tech sky130A
magscale 1 2
timestamp 1647448289
<< viali >>
rect 2237 41157 2271 41191
rect 7941 41157 7975 41191
rect 24869 41157 24903 41191
rect 34897 41157 34931 41191
rect 41889 41157 41923 41191
rect 1869 41089 1903 41123
rect 2881 41089 2915 41123
rect 3801 41021 3835 41055
rect 3985 41021 4019 41055
rect 4813 41021 4847 41055
rect 12909 41021 12943 41055
rect 13369 41021 13403 41055
rect 13553 41021 13587 41055
rect 21833 41021 21867 41055
rect 22017 41021 22051 41055
rect 22293 41021 22327 41055
rect 33885 41021 33919 41055
rect 34713 41021 34747 41055
rect 35173 41021 35207 41055
rect 40049 41021 40083 41055
rect 40233 41021 40267 41055
rect 2789 40885 2823 40919
rect 8033 40885 8067 40919
rect 10977 40885 11011 40919
rect 14105 40885 14139 40919
rect 14749 40885 14783 40919
rect 20177 40885 20211 40919
rect 24961 40885 24995 40919
rect 26065 40885 26099 40919
rect 26985 40885 27019 40919
rect 29561 40885 29595 40919
rect 31585 40885 31619 40919
rect 32597 40885 32631 40919
rect 38485 40885 38519 40919
rect 39313 40885 39347 40919
rect 22477 40681 22511 40715
rect 9873 40613 9907 40647
rect 2053 40545 2087 40579
rect 5181 40545 5215 40579
rect 10977 40545 11011 40579
rect 11621 40545 11655 40579
rect 14105 40545 14139 40579
rect 14565 40545 14599 40579
rect 20177 40545 20211 40579
rect 20729 40545 20763 40579
rect 24869 40545 24903 40579
rect 26709 40545 26743 40579
rect 27169 40545 27203 40579
rect 29561 40545 29595 40579
rect 30021 40545 30055 40579
rect 32321 40545 32355 40579
rect 32873 40545 32907 40579
rect 36093 40545 36127 40579
rect 37473 40545 37507 40579
rect 39313 40545 39347 40579
rect 41889 40545 41923 40579
rect 3249 40477 3283 40511
rect 4261 40477 4295 40511
rect 4721 40477 4755 40511
rect 9229 40477 9263 40511
rect 10333 40477 10367 40511
rect 13369 40477 13403 40511
rect 23305 40477 23339 40511
rect 24409 40477 24443 40511
rect 37013 40477 37047 40511
rect 40325 40477 40359 40511
rect 3065 40409 3099 40443
rect 4905 40409 4939 40443
rect 10425 40409 10459 40443
rect 11161 40409 11195 40443
rect 14289 40409 14323 40443
rect 20361 40409 20395 40443
rect 24593 40409 24627 40443
rect 26893 40409 26927 40443
rect 29745 40409 29779 40443
rect 32505 40409 32539 40443
rect 36829 40409 36863 40443
rect 37657 40409 37691 40443
rect 40509 40409 40543 40443
rect 13461 40341 13495 40375
rect 4077 40137 4111 40171
rect 20361 40137 20395 40171
rect 21925 40137 21959 40171
rect 29377 40137 29411 40171
rect 38301 40137 38335 40171
rect 1869 40069 1903 40103
rect 3525 40069 3559 40103
rect 14289 40069 14323 40103
rect 32321 40069 32355 40103
rect 35081 40069 35115 40103
rect 36737 40069 36771 40103
rect 41889 40069 41923 40103
rect 4169 40001 4203 40035
rect 4721 40001 4755 40035
rect 4813 40001 4847 40035
rect 5641 40001 5675 40035
rect 5733 40001 5767 40035
rect 9137 40001 9171 40035
rect 20269 40001 20303 40035
rect 21833 40001 21867 40035
rect 25973 40001 26007 40035
rect 26065 40001 26099 40035
rect 26985 40001 27019 40035
rect 29285 40001 29319 40035
rect 31401 40001 31435 40035
rect 31493 40001 31527 40035
rect 32137 40001 32171 40035
rect 38209 40001 38243 40035
rect 40049 40001 40083 40035
rect 1685 39933 1719 39967
rect 9321 39933 9355 39967
rect 9689 39933 9723 39967
rect 12265 39933 12299 39967
rect 13277 39933 13311 39967
rect 13461 39933 13495 39967
rect 14105 39933 14139 39967
rect 15945 39933 15979 39967
rect 23305 39933 23339 39967
rect 23489 39933 23523 39967
rect 23857 39933 23891 39967
rect 27169 39933 27203 39967
rect 27445 39933 27479 39967
rect 32597 39933 32631 39967
rect 34897 39933 34931 39967
rect 40233 39933 40267 39967
rect 6377 39797 6411 39831
rect 39589 39797 39623 39831
rect 3801 39593 3835 39627
rect 9321 39593 9355 39627
rect 12541 39593 12575 39627
rect 13185 39593 13219 39627
rect 14197 39593 14231 39627
rect 23397 39593 23431 39627
rect 26709 39593 26743 39627
rect 32781 39593 32815 39627
rect 33977 39593 34011 39627
rect 34805 39593 34839 39627
rect 35817 39593 35851 39627
rect 36553 39593 36587 39627
rect 40049 39593 40083 39627
rect 41337 39593 41371 39627
rect 41981 39593 42015 39627
rect 39313 39525 39347 39559
rect 2881 39457 2915 39491
rect 5273 39457 5307 39491
rect 6469 39457 6503 39491
rect 1409 39389 1443 39423
rect 9229 39389 9263 39423
rect 10241 39389 10275 39423
rect 11621 39389 11655 39423
rect 12449 39389 12483 39423
rect 13093 39389 13127 39423
rect 14105 39389 14139 39423
rect 22753 39389 22787 39423
rect 22845 39389 22879 39423
rect 26617 39389 26651 39423
rect 32873 39389 32907 39423
rect 33885 39389 33919 39423
rect 34713 39389 34747 39423
rect 35909 39389 35943 39423
rect 39957 39389 39991 39423
rect 40785 39389 40819 39423
rect 41429 39389 41463 39423
rect 41889 39389 41923 39423
rect 1593 39321 1627 39355
rect 6285 39321 6319 39355
rect 11069 39321 11103 39355
rect 10425 39253 10459 39287
rect 40693 39253 40727 39287
rect 2145 39049 2179 39083
rect 4813 39049 4847 39083
rect 23397 39049 23431 39083
rect 40233 38981 40267 39015
rect 41889 38981 41923 39015
rect 1593 38913 1627 38947
rect 2237 38913 2271 38947
rect 3801 38913 3835 38947
rect 4721 38913 4755 38947
rect 8861 38913 8895 38947
rect 9597 38913 9631 38947
rect 10885 38913 10919 38947
rect 11529 38913 11563 38947
rect 13185 38913 13219 38947
rect 23305 38913 23339 38947
rect 32689 38913 32723 38947
rect 32873 38913 32907 38947
rect 33517 38913 33551 38947
rect 35265 38913 35299 38947
rect 36001 38913 36035 38947
rect 36185 38913 36219 38947
rect 36277 38913 36311 38947
rect 37933 38913 37967 38947
rect 38117 38913 38151 38947
rect 10333 38845 10367 38879
rect 12357 38845 12391 38879
rect 39589 38845 39623 38879
rect 40049 38845 40083 38879
rect 33057 38709 33091 38743
rect 33701 38709 33735 38743
rect 36001 38709 36035 38743
rect 38117 38709 38151 38743
rect 1685 38505 1719 38539
rect 30941 38505 30975 38539
rect 36921 38505 36955 38539
rect 31125 38437 31159 38471
rect 9229 38369 9263 38403
rect 25237 38369 25271 38403
rect 31585 38369 31619 38403
rect 41337 38369 41371 38403
rect 2789 38301 2823 38335
rect 3985 38301 4019 38335
rect 8953 38301 8987 38335
rect 10885 38301 10919 38335
rect 24961 38301 24995 38335
rect 25145 38301 25179 38335
rect 25881 38301 25915 38335
rect 26065 38301 26099 38335
rect 30205 38301 30239 38335
rect 31861 38301 31895 38335
rect 33802 38301 33836 38335
rect 34069 38301 34103 38335
rect 35541 38301 35575 38335
rect 38678 38301 38712 38335
rect 38945 38301 38979 38335
rect 42165 38301 42199 38335
rect 11713 38233 11747 38267
rect 30757 38233 30791 38267
rect 30973 38233 31007 38267
rect 31953 38233 31987 38267
rect 35808 38233 35842 38267
rect 41981 38233 42015 38267
rect 3893 38165 3927 38199
rect 24777 38165 24811 38199
rect 26249 38165 26283 38199
rect 30021 38165 30055 38199
rect 31769 38165 31803 38199
rect 32137 38165 32171 38199
rect 32689 38165 32723 38199
rect 37565 38165 37599 38199
rect 23949 37961 23983 37995
rect 29377 37961 29411 37995
rect 31217 37961 31251 37995
rect 32689 37961 32723 37995
rect 36277 37961 36311 37995
rect 38117 37961 38151 37995
rect 38945 37961 38979 37995
rect 41153 37961 41187 37995
rect 41705 37961 41739 37995
rect 4261 37893 4295 37927
rect 11989 37893 12023 37927
rect 32505 37893 32539 37927
rect 4445 37825 4479 37859
rect 11621 37825 11655 37859
rect 17500 37825 17534 37859
rect 21833 37825 21867 37859
rect 22089 37825 22123 37859
rect 23857 37825 23891 37859
rect 24133 37825 24167 37859
rect 25053 37825 25087 37859
rect 25309 37825 25343 37859
rect 27997 37825 28031 37859
rect 28264 37825 28298 37859
rect 29837 37825 29871 37859
rect 30104 37825 30138 37859
rect 32137 37825 32171 37859
rect 34538 37825 34572 37859
rect 36553 37825 36587 37859
rect 38393 37825 38427 37859
rect 38853 37825 38887 37859
rect 39129 37825 39163 37859
rect 40040 37825 40074 37859
rect 41613 37825 41647 37859
rect 2789 37757 2823 37791
rect 17233 37757 17267 37791
rect 34805 37757 34839 37791
rect 36277 37757 36311 37791
rect 36461 37757 36495 37791
rect 38117 37757 38151 37791
rect 39773 37757 39807 37791
rect 1685 37621 1719 37655
rect 18613 37621 18647 37655
rect 23213 37621 23247 37655
rect 24317 37621 24351 37655
rect 26433 37621 26467 37655
rect 32505 37621 32539 37655
rect 33425 37621 33459 37655
rect 38301 37621 38335 37655
rect 39313 37621 39347 37655
rect 17417 37417 17451 37451
rect 22937 37417 22971 37451
rect 25145 37417 25179 37451
rect 28825 37417 28859 37451
rect 30113 37417 30147 37451
rect 31125 37417 31159 37451
rect 31677 37417 31711 37451
rect 33333 37417 33367 37451
rect 39129 37417 39163 37451
rect 40049 37417 40083 37451
rect 41797 37417 41831 37451
rect 29929 37349 29963 37383
rect 38761 37349 38795 37383
rect 1409 37281 1443 37315
rect 17693 37281 17727 37315
rect 23121 37281 23155 37315
rect 37565 37281 37599 37315
rect 3249 37213 3283 37247
rect 4997 37213 5031 37247
rect 15485 37213 15519 37247
rect 17601 37213 17635 37247
rect 18521 37213 18555 37247
rect 20637 37213 20671 37247
rect 21097 37213 21131 37247
rect 23213 37213 23247 37247
rect 24409 37213 24443 37247
rect 25329 37213 25363 37247
rect 25421 37213 25455 37247
rect 26341 37213 26375 37247
rect 29653 37213 29687 37247
rect 30665 37213 30699 37247
rect 30941 37213 30975 37247
rect 31861 37213 31895 37247
rect 32045 37213 32079 37247
rect 32965 37213 32999 37247
rect 33977 37213 34011 37247
rect 36093 37213 36127 37247
rect 36369 37213 36403 37247
rect 37197 37213 37231 37247
rect 37682 37213 37716 37247
rect 39865 37213 39899 37247
rect 1593 37145 1627 37179
rect 4353 37145 4387 37179
rect 15730 37145 15764 37179
rect 20370 37145 20404 37179
rect 21342 37145 21376 37179
rect 24501 37145 24535 37179
rect 26608 37145 26642 37179
rect 29009 37145 29043 37179
rect 31585 37145 31619 37179
rect 33333 37145 33367 37179
rect 39129 37145 39163 37179
rect 16865 37077 16899 37111
rect 18061 37077 18095 37111
rect 18705 37077 18739 37111
rect 19257 37077 19291 37111
rect 22477 37077 22511 37111
rect 23581 37077 23615 37111
rect 25789 37077 25823 37111
rect 27721 37077 27755 37111
rect 28641 37077 28675 37111
rect 28809 37077 28843 37111
rect 30757 37077 30791 37111
rect 32229 37077 32263 37111
rect 33517 37077 33551 37111
rect 34161 37077 34195 37111
rect 35909 37077 35943 37111
rect 36277 37077 36311 37111
rect 37473 37077 37507 37111
rect 37841 37077 37875 37111
rect 39313 37077 39347 37111
rect 2053 36873 2087 36907
rect 15577 36873 15611 36907
rect 18613 36873 18647 36907
rect 20361 36873 20395 36907
rect 21097 36873 21131 36907
rect 23213 36873 23247 36907
rect 25789 36873 25823 36907
rect 28273 36873 28307 36907
rect 28917 36873 28951 36907
rect 29561 36873 29595 36907
rect 31309 36873 31343 36907
rect 36553 36873 36587 36907
rect 38577 36873 38611 36907
rect 39221 36873 39255 36907
rect 23673 36805 23707 36839
rect 29929 36805 29963 36839
rect 38209 36805 38243 36839
rect 39389 36805 39423 36839
rect 39589 36805 39623 36839
rect 2145 36737 2179 36771
rect 3525 36737 3559 36771
rect 4261 36737 4295 36771
rect 5825 36737 5859 36771
rect 14197 36737 14231 36771
rect 14289 36737 14323 36771
rect 14473 36737 14507 36771
rect 15853 36737 15887 36771
rect 17509 36737 17543 36771
rect 17693 36737 17727 36771
rect 18429 36737 18463 36771
rect 20269 36737 20303 36771
rect 20453 36737 20487 36771
rect 20913 36737 20947 36771
rect 22753 36737 22787 36771
rect 23397 36737 23431 36771
rect 25421 36737 25455 36771
rect 26433 36737 26467 36771
rect 28457 36737 28491 36771
rect 28917 36737 28951 36771
rect 29101 36737 29135 36771
rect 29745 36737 29779 36771
rect 31493 36737 31527 36771
rect 32413 36737 32447 36771
rect 35440 36737 35474 36771
rect 38393 36737 38427 36771
rect 38485 36737 38519 36771
rect 41613 36737 41647 36771
rect 3249 36669 3283 36703
rect 4905 36669 4939 36703
rect 15577 36669 15611 36703
rect 17233 36669 17267 36703
rect 18245 36669 18279 36703
rect 22477 36669 22511 36703
rect 23489 36669 23523 36703
rect 24133 36669 24167 36703
rect 24409 36669 24443 36703
rect 25513 36669 25547 36703
rect 32689 36669 32723 36703
rect 35173 36669 35207 36703
rect 38761 36601 38795 36635
rect 5641 36533 5675 36567
rect 14381 36533 14415 36567
rect 15761 36533 15795 36567
rect 17325 36533 17359 36567
rect 22569 36533 22603 36567
rect 22661 36533 22695 36567
rect 23489 36533 23523 36567
rect 25421 36533 25455 36567
rect 26341 36533 26375 36567
rect 39405 36533 39439 36567
rect 41705 36533 41739 36567
rect 15945 36329 15979 36363
rect 16957 36329 16991 36363
rect 17233 36329 17267 36363
rect 17693 36329 17727 36363
rect 21925 36329 21959 36363
rect 23765 36329 23799 36363
rect 24501 36329 24535 36363
rect 24869 36329 24903 36363
rect 26617 36329 26651 36363
rect 35909 36329 35943 36363
rect 39037 36329 39071 36363
rect 33885 36261 33919 36295
rect 38393 36261 38427 36295
rect 16957 36193 16991 36227
rect 18153 36193 18187 36227
rect 24409 36193 24443 36227
rect 25973 36193 26007 36227
rect 33241 36193 33275 36227
rect 33425 36193 33459 36227
rect 38853 36193 38887 36227
rect 41337 36193 41371 36227
rect 41981 36193 42015 36227
rect 2053 36125 2087 36159
rect 2881 36125 2915 36159
rect 4353 36125 4387 36159
rect 14105 36125 14139 36159
rect 14372 36125 14406 36159
rect 16129 36125 16163 36159
rect 16221 36125 16255 36159
rect 16865 36125 16899 36159
rect 17877 36125 17911 36159
rect 18061 36125 18095 36159
rect 19257 36125 19291 36159
rect 21925 36125 21959 36159
rect 22017 36125 22051 36159
rect 22201 36125 22235 36159
rect 23581 36125 23615 36159
rect 24685 36125 24719 36159
rect 25697 36125 25731 36159
rect 25789 36125 25823 36159
rect 26433 36125 26467 36159
rect 29745 36125 29779 36159
rect 30665 36125 30699 36159
rect 30757 36125 30791 36159
rect 33149 36125 33183 36159
rect 34161 36125 34195 36159
rect 36553 36125 36587 36159
rect 36645 36125 36679 36159
rect 36829 36125 36863 36159
rect 37473 36125 37507 36159
rect 38117 36125 38151 36159
rect 39129 36125 39163 36159
rect 42165 36125 42199 36159
rect 4997 36057 5031 36091
rect 23397 36057 23431 36091
rect 33425 36057 33459 36091
rect 33885 36057 33919 36091
rect 36093 36057 36127 36091
rect 38393 36057 38427 36091
rect 38853 36057 38887 36091
rect 2789 35989 2823 36023
rect 15485 35989 15519 36023
rect 19349 35989 19383 36023
rect 25697 35989 25731 36023
rect 29561 35989 29595 36023
rect 30941 35989 30975 36023
rect 34069 35989 34103 36023
rect 35725 35989 35759 36023
rect 35893 35989 35927 36023
rect 36553 35989 36587 36023
rect 37657 35989 37691 36023
rect 38209 35989 38243 36023
rect 14565 35785 14599 35819
rect 17141 35785 17175 35819
rect 24409 35785 24443 35819
rect 30297 35785 30331 35819
rect 32321 35785 32355 35819
rect 32413 35785 32447 35819
rect 35633 35785 35667 35819
rect 2145 35717 2179 35751
rect 15945 35717 15979 35751
rect 28724 35717 28758 35751
rect 30481 35717 30515 35751
rect 34538 35717 34572 35751
rect 40110 35717 40144 35751
rect 1961 35649 1995 35683
rect 5089 35649 5123 35683
rect 14841 35649 14875 35683
rect 16129 35649 16163 35683
rect 16681 35649 16715 35683
rect 16773 35649 16807 35683
rect 16957 35649 16991 35683
rect 17601 35649 17635 35683
rect 19625 35649 19659 35683
rect 19717 35649 19751 35683
rect 19809 35649 19843 35683
rect 19993 35649 20027 35683
rect 22937 35649 22971 35683
rect 23949 35649 23983 35683
rect 24409 35649 24443 35683
rect 24593 35649 24627 35683
rect 25237 35649 25271 35683
rect 25421 35649 25455 35683
rect 25513 35649 25547 35683
rect 25789 35649 25823 35683
rect 27353 35649 27387 35683
rect 28457 35649 28491 35683
rect 32505 35649 32539 35683
rect 35817 35649 35851 35683
rect 41889 35649 41923 35683
rect 2881 35581 2915 35615
rect 4813 35581 4847 35615
rect 14565 35581 14599 35615
rect 15761 35581 15795 35615
rect 22661 35581 22695 35615
rect 27261 35581 27295 35615
rect 34805 35581 34839 35615
rect 38577 35581 38611 35615
rect 38853 35581 38887 35615
rect 39865 35581 39899 35615
rect 22845 35513 22879 35547
rect 25605 35513 25639 35547
rect 29837 35513 29871 35547
rect 30849 35513 30883 35547
rect 32137 35513 32171 35547
rect 32689 35513 32723 35547
rect 33425 35513 33459 35547
rect 14749 35445 14783 35479
rect 17693 35445 17727 35479
rect 19349 35445 19383 35479
rect 22753 35445 22787 35479
rect 23857 35445 23891 35479
rect 25697 35445 25731 35479
rect 26985 35445 27019 35479
rect 30481 35445 30515 35479
rect 41245 35445 41279 35479
rect 15577 35241 15611 35275
rect 19901 35241 19935 35275
rect 23213 35241 23247 35275
rect 24777 35241 24811 35275
rect 24869 35241 24903 35275
rect 30941 35241 30975 35275
rect 38669 35173 38703 35207
rect 40049 35173 40083 35207
rect 15761 35105 15795 35139
rect 16957 35105 16991 35139
rect 18429 35105 18463 35139
rect 18705 35105 18739 35139
rect 21833 35105 21867 35139
rect 24685 35105 24719 35139
rect 29561 35105 29595 35139
rect 32781 35105 32815 35139
rect 38485 35105 38519 35139
rect 15577 35037 15611 35071
rect 15853 35037 15887 35071
rect 17233 35037 17267 35071
rect 18337 35037 18371 35071
rect 19257 35037 19291 35071
rect 19405 35037 19439 35071
rect 19722 35037 19756 35071
rect 24961 35037 24995 35071
rect 25651 35037 25685 35071
rect 25881 35037 25915 35071
rect 26009 35037 26043 35071
rect 26157 35037 26191 35071
rect 26617 35037 26651 35071
rect 26710 35037 26744 35071
rect 27082 35037 27116 35071
rect 32045 35037 32079 35071
rect 32321 35037 32355 35071
rect 33057 35037 33091 35071
rect 35541 35037 35575 35071
rect 35725 35037 35759 35071
rect 38025 35037 38059 35071
rect 38761 35037 38795 35071
rect 39865 35037 39899 35071
rect 40049 35037 40083 35071
rect 40693 35037 40727 35071
rect 41337 35037 41371 35071
rect 41981 35037 42015 35071
rect 15945 34969 15979 35003
rect 19533 34969 19567 35003
rect 19625 34969 19659 35003
rect 22100 34969 22134 35003
rect 25789 34969 25823 35003
rect 26893 34969 26927 35003
rect 26985 34969 27019 35003
rect 29828 34969 29862 35003
rect 37758 34969 37792 35003
rect 38485 34969 38519 35003
rect 25513 34901 25547 34935
rect 27261 34901 27295 34935
rect 31861 34901 31895 34935
rect 32229 34901 32263 34935
rect 35633 34901 35667 34935
rect 36645 34901 36679 34935
rect 41429 34901 41463 34935
rect 16957 34697 16991 34731
rect 22201 34697 22235 34731
rect 30297 34697 30331 34731
rect 30849 34697 30883 34731
rect 31217 34697 31251 34731
rect 33149 34697 33183 34731
rect 37933 34697 37967 34731
rect 39129 34697 39163 34731
rect 19438 34629 19472 34663
rect 32505 34629 32539 34663
rect 33301 34629 33335 34663
rect 33517 34629 33551 34663
rect 35072 34629 35106 34663
rect 37565 34629 37599 34663
rect 37770 34629 37804 34663
rect 38485 34629 38519 34663
rect 40233 34629 40267 34663
rect 41889 34629 41923 34663
rect 14473 34561 14507 34595
rect 14841 34561 14875 34595
rect 15485 34561 15519 34595
rect 15577 34561 15611 34595
rect 16681 34561 16715 34595
rect 18153 34561 18187 34595
rect 18245 34561 18279 34595
rect 18429 34561 18463 34595
rect 19080 34561 19114 34595
rect 19193 34561 19227 34595
rect 19349 34561 19383 34595
rect 19557 34561 19591 34595
rect 20913 34561 20947 34595
rect 22385 34561 22419 34595
rect 22569 34561 22603 34595
rect 22661 34561 22695 34595
rect 23673 34561 23707 34595
rect 25329 34561 25363 34595
rect 25513 34561 25547 34595
rect 25605 34561 25639 34595
rect 25697 34561 25731 34595
rect 27169 34561 27203 34595
rect 29929 34561 29963 34595
rect 30389 34561 30423 34595
rect 31033 34561 31067 34595
rect 31309 34561 31343 34595
rect 32137 34561 32171 34595
rect 34161 34561 34195 34595
rect 38945 34561 38979 34595
rect 14565 34493 14599 34527
rect 15301 34493 15335 34527
rect 16957 34493 16991 34527
rect 18337 34493 18371 34527
rect 22293 34493 22327 34527
rect 23581 34493 23615 34527
rect 25973 34493 26007 34527
rect 34805 34493 34839 34527
rect 38761 34493 38795 34527
rect 40049 34493 40083 34527
rect 15393 34425 15427 34459
rect 16773 34425 16807 34459
rect 17969 34425 18003 34459
rect 19717 34425 19751 34459
rect 24041 34425 24075 34459
rect 32689 34425 32723 34459
rect 14381 34357 14415 34391
rect 14749 34357 14783 34391
rect 21097 34357 21131 34391
rect 27077 34357 27111 34391
rect 30113 34357 30147 34391
rect 32505 34357 32539 34391
rect 33333 34357 33367 34391
rect 33977 34357 34011 34391
rect 36185 34357 36219 34391
rect 37749 34357 37783 34391
rect 38669 34357 38703 34391
rect 18521 34153 18555 34187
rect 20177 34153 20211 34187
rect 27169 34153 27203 34187
rect 29837 34153 29871 34187
rect 30205 34153 30239 34187
rect 31953 34153 31987 34187
rect 35265 34153 35299 34187
rect 35909 34153 35943 34187
rect 36921 34153 36955 34187
rect 37565 34153 37599 34187
rect 38301 34153 38335 34187
rect 15485 34085 15519 34119
rect 16957 34085 16991 34119
rect 18613 34085 18647 34119
rect 20729 34085 20763 34119
rect 27353 34085 27387 34119
rect 38853 34085 38887 34119
rect 16497 34017 16531 34051
rect 30297 34017 30331 34051
rect 35173 34017 35207 34051
rect 36277 34017 36311 34051
rect 37105 34017 37139 34051
rect 39865 34017 39899 34051
rect 14105 33949 14139 33983
rect 14372 33949 14406 33983
rect 16589 33949 16623 33983
rect 18153 33949 18187 33983
rect 18337 33949 18371 33983
rect 18429 33949 18463 33983
rect 18705 33949 18739 33983
rect 20085 33949 20119 33983
rect 21842 33949 21876 33983
rect 22109 33949 22143 33983
rect 26341 33949 26375 33983
rect 26525 33949 26559 33983
rect 27813 33949 27847 33983
rect 30021 33949 30055 33983
rect 33333 33949 33367 33983
rect 35357 33949 35391 33983
rect 35449 33949 35483 33983
rect 36093 33949 36127 33983
rect 36829 33949 36863 33983
rect 37565 33949 37599 33983
rect 37749 33949 37783 33983
rect 38669 33949 38703 33983
rect 40132 33949 40166 33983
rect 41705 33949 41739 33983
rect 26985 33881 27019 33915
rect 33088 33881 33122 33915
rect 37105 33881 37139 33915
rect 38577 33881 38611 33915
rect 26525 33813 26559 33847
rect 27185 33813 27219 33847
rect 27997 33813 28031 33847
rect 38485 33813 38519 33847
rect 41245 33813 41279 33847
rect 41797 33813 41831 33847
rect 16773 33609 16807 33643
rect 21833 33609 21867 33643
rect 27537 33609 27571 33643
rect 18981 33541 19015 33575
rect 19191 33541 19225 33575
rect 19901 33541 19935 33575
rect 21005 33541 21039 33575
rect 21985 33541 22019 33575
rect 22201 33541 22235 33575
rect 28650 33541 28684 33575
rect 33241 33541 33275 33575
rect 39221 33541 39255 33575
rect 41705 33541 41739 33575
rect 16865 33473 16899 33507
rect 18889 33473 18923 33507
rect 19073 33473 19107 33507
rect 20729 33473 20763 33507
rect 20913 33473 20947 33507
rect 21097 33473 21131 33507
rect 23029 33473 23063 33507
rect 23857 33473 23891 33507
rect 24961 33473 24995 33507
rect 25145 33473 25179 33507
rect 25605 33473 25639 33507
rect 25789 33473 25823 33507
rect 26249 33473 26283 33507
rect 26433 33473 26467 33507
rect 28917 33473 28951 33507
rect 32321 33473 32355 33507
rect 32505 33473 32539 33507
rect 33057 33473 33091 33507
rect 38209 33473 38243 33507
rect 41889 33473 41923 33507
rect 19349 33405 19383 33439
rect 38393 33405 38427 33439
rect 41337 33405 41371 33439
rect 21281 33337 21315 33371
rect 32413 33337 32447 33371
rect 38853 33337 38887 33371
rect 18705 33269 18739 33303
rect 19993 33269 20027 33303
rect 22017 33269 22051 33303
rect 23121 33269 23155 33303
rect 23673 33269 23707 33303
rect 24777 33269 24811 33303
rect 25697 33269 25731 33303
rect 26249 33269 26283 33303
rect 38025 33269 38059 33303
rect 39221 33269 39255 33303
rect 39405 33269 39439 33303
rect 18613 33065 18647 33099
rect 21281 33065 21315 33099
rect 26801 33065 26835 33099
rect 30113 33065 30147 33099
rect 32321 33065 32355 33099
rect 33241 33065 33275 33099
rect 38577 33065 38611 33099
rect 19349 32997 19383 33031
rect 23857 32997 23891 33031
rect 30941 32997 30975 33031
rect 19809 32929 19843 32963
rect 27905 32929 27939 32963
rect 32229 32929 32263 32963
rect 34989 32929 35023 32963
rect 38117 32929 38151 32963
rect 15301 32861 15335 32895
rect 16681 32861 16715 32895
rect 16865 32861 16899 32895
rect 17049 32861 17083 32895
rect 17785 32861 17819 32895
rect 17877 32861 17911 32895
rect 18521 32861 18555 32895
rect 18705 32861 18739 32895
rect 20085 32861 20119 32895
rect 20545 32861 20579 32895
rect 20729 32861 20763 32895
rect 21373 32861 21407 32895
rect 22477 32861 22511 32895
rect 22744 32861 22778 32895
rect 24593 32861 24627 32895
rect 24777 32861 24811 32895
rect 24895 32861 24929 32895
rect 25053 32861 25087 32895
rect 25513 32861 25547 32895
rect 25789 32861 25823 32895
rect 26939 32861 26973 32895
rect 27077 32861 27111 32895
rect 27353 32861 27387 32895
rect 27813 32861 27847 32895
rect 29929 32861 29963 32895
rect 30757 32861 30791 32895
rect 31493 32861 31527 32895
rect 32137 32861 32171 32895
rect 32413 32861 32447 32895
rect 33057 32861 33091 32895
rect 33241 32861 33275 32895
rect 34713 32861 34747 32895
rect 34805 32861 34839 32895
rect 36829 32861 36863 32895
rect 38209 32861 38243 32895
rect 38577 32861 38611 32895
rect 40325 32861 40359 32895
rect 19349 32793 19383 32827
rect 20637 32793 20671 32827
rect 24685 32793 24719 32827
rect 27169 32793 27203 32827
rect 36553 32793 36587 32827
rect 36737 32793 36771 32827
rect 40509 32793 40543 32827
rect 42165 32793 42199 32827
rect 15117 32725 15151 32759
rect 18061 32725 18095 32759
rect 19901 32725 19935 32759
rect 24409 32725 24443 32759
rect 31585 32725 31619 32759
rect 32597 32725 32631 32759
rect 33425 32725 33459 32759
rect 34989 32725 35023 32759
rect 36651 32725 36685 32759
rect 38761 32725 38795 32759
rect 18613 32521 18647 32555
rect 19073 32521 19107 32555
rect 20361 32521 20395 32555
rect 23397 32521 23431 32555
rect 26249 32521 26283 32555
rect 27077 32521 27111 32555
rect 28917 32521 28951 32555
rect 35909 32521 35943 32555
rect 36461 32521 36495 32555
rect 38669 32521 38703 32555
rect 39497 32521 39531 32555
rect 21189 32453 21223 32487
rect 37534 32453 37568 32487
rect 14473 32385 14507 32419
rect 14740 32385 14774 32419
rect 17500 32385 17534 32419
rect 19257 32385 19291 32419
rect 19441 32385 19475 32419
rect 20177 32385 20211 32419
rect 20361 32385 20395 32419
rect 23213 32385 23247 32419
rect 23949 32385 23983 32419
rect 24225 32385 24259 32419
rect 24961 32385 24995 32419
rect 25329 32385 25363 32419
rect 25789 32385 25823 32419
rect 26065 32385 26099 32419
rect 27169 32385 27203 32419
rect 28641 32385 28675 32419
rect 28733 32385 28767 32419
rect 29377 32385 29411 32419
rect 29644 32385 29678 32419
rect 31493 32385 31527 32419
rect 32689 32385 32723 32419
rect 34152 32385 34186 32419
rect 35725 32385 35759 32419
rect 36001 32385 36035 32419
rect 36737 32385 36771 32419
rect 37289 32385 37323 32419
rect 39129 32385 39163 32419
rect 39957 32385 39991 32419
rect 40224 32385 40258 32419
rect 17233 32317 17267 32351
rect 23029 32317 23063 32351
rect 25973 32317 26007 32351
rect 31217 32317 31251 32351
rect 32505 32317 32539 32351
rect 33885 32317 33919 32351
rect 36461 32317 36495 32351
rect 39221 32317 39255 32351
rect 21005 32249 21039 32283
rect 31309 32249 31343 32283
rect 31401 32249 31435 32283
rect 35725 32249 35759 32283
rect 15853 32181 15887 32215
rect 25329 32181 25363 32215
rect 25789 32181 25823 32215
rect 30757 32181 30791 32215
rect 35265 32181 35299 32215
rect 36645 32181 36679 32215
rect 39221 32181 39255 32215
rect 41337 32181 41371 32215
rect 17233 31977 17267 32011
rect 18245 31977 18279 32011
rect 24961 31977 24995 32011
rect 27169 31977 27203 32011
rect 15485 31909 15519 31943
rect 32321 31909 32355 31943
rect 14105 31841 14139 31875
rect 15945 31841 15979 31875
rect 20361 31841 20395 31875
rect 20453 31841 20487 31875
rect 26709 31841 26743 31875
rect 28549 31841 28583 31875
rect 30021 31841 30055 31875
rect 31861 31841 31895 31875
rect 33609 31841 33643 31875
rect 34713 31841 34747 31875
rect 34989 31841 35023 31875
rect 38393 31841 38427 31875
rect 38669 31841 38703 31875
rect 41337 31841 41371 31875
rect 16221 31773 16255 31807
rect 17417 31773 17451 31807
rect 17785 31773 17819 31807
rect 18429 31773 18463 31807
rect 20545 31773 20579 31807
rect 20637 31773 20671 31807
rect 22661 31773 22695 31807
rect 24869 31773 24903 31807
rect 26065 31773 26099 31807
rect 26228 31773 26262 31807
rect 26344 31773 26378 31807
rect 26453 31773 26487 31807
rect 28282 31773 28316 31807
rect 30205 31773 30239 31807
rect 30941 31773 30975 31807
rect 31125 31773 31159 31807
rect 31677 31773 31711 31807
rect 32873 31773 32907 31807
rect 33333 31773 33367 31807
rect 37013 31773 37047 31807
rect 37289 31773 37323 31807
rect 42165 31773 42199 31807
rect 14372 31705 14406 31739
rect 17509 31705 17543 31739
rect 17601 31705 17635 31739
rect 22394 31705 22428 31739
rect 32689 31705 32723 31739
rect 41981 31705 42015 31739
rect 20821 31637 20855 31671
rect 21281 31637 21315 31671
rect 30757 31637 30791 31671
rect 32505 31637 32539 31671
rect 32597 31637 32631 31671
rect 14289 31433 14323 31467
rect 15945 31433 15979 31467
rect 21281 31433 21315 31467
rect 26157 31433 26191 31467
rect 26985 31433 27019 31467
rect 29837 31433 29871 31467
rect 32337 31433 32371 31467
rect 34069 31433 34103 31467
rect 35633 31433 35667 31467
rect 38301 31433 38335 31467
rect 38485 31433 38519 31467
rect 39129 31433 39163 31467
rect 39497 31433 39531 31467
rect 40233 31433 40267 31467
rect 41521 31433 41555 31467
rect 15577 31365 15611 31399
rect 21925 31365 21959 31399
rect 24317 31365 24351 31399
rect 28457 31365 28491 31399
rect 32137 31365 32171 31399
rect 33425 31365 33459 31399
rect 33609 31365 33643 31399
rect 35541 31365 35575 31399
rect 35817 31365 35851 31399
rect 38209 31365 38243 31399
rect 14565 31297 14599 31331
rect 14657 31297 14691 31331
rect 14749 31297 14783 31331
rect 14933 31297 14967 31331
rect 15761 31297 15795 31331
rect 16681 31297 16715 31331
rect 16957 31297 16991 31331
rect 20637 31297 20671 31331
rect 20821 31297 20855 31331
rect 20913 31297 20947 31331
rect 21005 31297 21039 31331
rect 22017 31297 22051 31331
rect 23397 31297 23431 31331
rect 23581 31297 23615 31331
rect 24501 31297 24535 31331
rect 25973 31297 26007 31331
rect 26249 31297 26283 31331
rect 27261 31297 27295 31331
rect 27445 31297 27479 31331
rect 28641 31297 28675 31331
rect 29745 31297 29779 31331
rect 29929 31297 29963 31331
rect 30573 31297 30607 31331
rect 30757 31297 30791 31331
rect 31401 31297 31435 31331
rect 31493 31297 31527 31331
rect 34253 31297 34287 31331
rect 34621 31297 34655 31331
rect 34713 31297 34747 31331
rect 35449 31297 35483 31331
rect 37933 31297 37967 31331
rect 38117 31297 38151 31331
rect 39313 31297 39347 31331
rect 39589 31297 39623 31331
rect 40049 31297 40083 31331
rect 40785 31297 40819 31331
rect 41429 31297 41463 31331
rect 27169 31229 27203 31263
rect 27353 31229 27387 31263
rect 31217 31229 31251 31263
rect 31309 31161 31343 31195
rect 32505 31161 32539 31195
rect 35265 31161 35299 31195
rect 23489 31093 23523 31127
rect 25789 31093 25823 31127
rect 30757 31093 30791 31127
rect 32321 31093 32355 31127
rect 34345 31093 34379 31127
rect 15025 30889 15059 30923
rect 17601 30889 17635 30923
rect 21373 30889 21407 30923
rect 22569 30889 22603 30923
rect 25789 30889 25823 30923
rect 32137 30889 32171 30923
rect 32781 30889 32815 30923
rect 34897 30889 34931 30923
rect 35081 30889 35115 30923
rect 35633 30889 35667 30923
rect 38577 30889 38611 30923
rect 38761 30889 38795 30923
rect 41521 30889 41555 30923
rect 28825 30821 28859 30855
rect 20453 30753 20487 30787
rect 23305 30753 23339 30787
rect 27169 30753 27203 30787
rect 32597 30753 32631 30787
rect 35817 30753 35851 30787
rect 14289 30685 14323 30719
rect 14381 30685 14415 30719
rect 14933 30685 14967 30719
rect 15117 30685 15151 30719
rect 15761 30685 15795 30719
rect 15853 30685 15887 30719
rect 16503 30685 16537 30719
rect 16681 30685 16715 30719
rect 16773 30685 16807 30719
rect 16865 30685 16899 30719
rect 17601 30685 17635 30719
rect 17785 30685 17819 30719
rect 20637 30685 20671 30719
rect 20913 30685 20947 30719
rect 21557 30685 21591 30719
rect 21833 30685 21867 30719
rect 23213 30685 23247 30719
rect 23397 30685 23431 30719
rect 24685 30685 24719 30719
rect 24777 30685 24811 30719
rect 24874 30685 24908 30719
rect 25053 30685 25087 30719
rect 27813 30685 27847 30719
rect 30757 30685 30791 30719
rect 31013 30685 31047 30719
rect 32873 30685 32907 30719
rect 35541 30685 35575 30719
rect 36277 30685 36311 30719
rect 36461 30685 36495 30719
rect 37473 30685 37507 30719
rect 37565 30685 37599 30719
rect 37749 30685 37783 30719
rect 41429 30685 41463 30719
rect 16037 30617 16071 30651
rect 22661 30617 22695 30651
rect 26924 30617 26958 30651
rect 28641 30617 28675 30651
rect 34713 30617 34747 30651
rect 35817 30617 35851 30651
rect 38393 30617 38427 30651
rect 14105 30549 14139 30583
rect 17141 30549 17175 30583
rect 20821 30549 20855 30583
rect 21741 30549 21775 30583
rect 24409 30549 24443 30583
rect 27629 30549 27663 30583
rect 32597 30549 32631 30583
rect 34913 30549 34947 30583
rect 36369 30549 36403 30583
rect 37933 30549 37967 30583
rect 38593 30549 38627 30583
rect 13185 30345 13219 30379
rect 15117 30345 15151 30379
rect 16681 30345 16715 30379
rect 20755 30345 20789 30379
rect 23305 30345 23339 30379
rect 25513 30345 25547 30379
rect 25881 30345 25915 30379
rect 27997 30345 28031 30379
rect 35357 30345 35391 30379
rect 20545 30277 20579 30311
rect 24418 30277 24452 30311
rect 28702 30277 28736 30311
rect 33425 30277 33459 30311
rect 33793 30277 33827 30311
rect 34437 30277 34471 30311
rect 13093 30209 13127 30243
rect 13369 30209 13403 30243
rect 14013 30209 14047 30243
rect 14197 30209 14231 30243
rect 14289 30209 14323 30243
rect 14381 30209 14415 30243
rect 14565 30209 14599 30243
rect 15209 30209 15243 30243
rect 16957 30209 16991 30243
rect 17325 30209 17359 30243
rect 17877 30209 17911 30243
rect 18061 30209 18095 30243
rect 19645 30209 19679 30243
rect 22293 30209 22327 30243
rect 24685 30209 24719 30243
rect 25697 30209 25731 30243
rect 25973 30209 26007 30243
rect 26985 30209 27019 30243
rect 27169 30209 27203 30243
rect 27813 30209 27847 30243
rect 28457 30209 28491 30243
rect 32689 30209 32723 30243
rect 32873 30209 32907 30243
rect 33333 30209 33367 30243
rect 33609 30209 33643 30243
rect 34805 30209 34839 30243
rect 36470 30209 36504 30243
rect 36737 30209 36771 30243
rect 37565 30209 37599 30243
rect 37832 30209 37866 30243
rect 39405 30209 39439 30243
rect 39672 30209 39706 30243
rect 41797 30209 41831 30243
rect 16865 30141 16899 30175
rect 17233 30141 17267 30175
rect 19901 30141 19935 30175
rect 27077 30141 27111 30175
rect 13829 30073 13863 30107
rect 17969 30073 18003 30107
rect 38945 30073 38979 30107
rect 13369 30005 13403 30039
rect 18521 30005 18555 30039
rect 20729 30005 20763 30039
rect 20913 30005 20947 30039
rect 22385 30005 22419 30039
rect 29837 30005 29871 30039
rect 32689 30005 32723 30039
rect 34253 30005 34287 30039
rect 34437 30005 34471 30039
rect 40785 30005 40819 30039
rect 22845 29801 22879 29835
rect 25881 29801 25915 29835
rect 26065 29801 26099 29835
rect 29561 29801 29595 29835
rect 29745 29801 29779 29835
rect 33977 29801 34011 29835
rect 36093 29801 36127 29835
rect 37749 29801 37783 29835
rect 39865 29801 39899 29835
rect 14381 29733 14415 29767
rect 17141 29733 17175 29767
rect 19901 29733 19935 29767
rect 23489 29733 23523 29767
rect 38117 29733 38151 29767
rect 40233 29733 40267 29767
rect 14473 29665 14507 29699
rect 29009 29665 29043 29699
rect 38669 29665 38703 29699
rect 38853 29665 38887 29699
rect 11713 29597 11747 29631
rect 14289 29597 14323 29631
rect 14565 29597 14599 29631
rect 14749 29597 14783 29631
rect 15209 29597 15243 29631
rect 15485 29597 15519 29631
rect 15761 29597 15795 29631
rect 15945 29597 15979 29631
rect 16497 29597 16531 29631
rect 18521 29597 18555 29631
rect 19257 29597 19291 29631
rect 19441 29597 19475 29631
rect 19533 29597 19567 29631
rect 19625 29597 19659 29631
rect 20453 29597 20487 29631
rect 22937 29597 22971 29631
rect 28733 29597 28767 29631
rect 30389 29597 30423 29631
rect 32597 29597 32631 29631
rect 32853 29597 32887 29631
rect 34713 29597 34747 29631
rect 39129 29597 39163 29631
rect 40049 29597 40083 29631
rect 40325 29597 40359 29631
rect 11980 29529 12014 29563
rect 18254 29529 18288 29563
rect 20720 29529 20754 29563
rect 23673 29529 23707 29563
rect 25145 29529 25179 29563
rect 25697 29529 25731 29563
rect 29929 29529 29963 29563
rect 30634 29529 30668 29563
rect 34958 29529 34992 29563
rect 37749 29529 37783 29563
rect 39037 29529 39071 29563
rect 42073 29529 42107 29563
rect 13093 29461 13127 29495
rect 14105 29461 14139 29495
rect 15301 29461 15335 29495
rect 16589 29461 16623 29495
rect 21833 29461 21867 29495
rect 24869 29461 24903 29495
rect 25897 29461 25931 29495
rect 29719 29461 29753 29495
rect 31769 29461 31803 29495
rect 37565 29461 37599 29495
rect 41981 29461 42015 29495
rect 15761 29257 15795 29291
rect 15929 29257 15963 29291
rect 20821 29257 20855 29291
rect 23581 29257 23615 29291
rect 28733 29257 28767 29291
rect 29837 29257 29871 29291
rect 34713 29257 34747 29291
rect 37841 29257 37875 29291
rect 12348 29189 12382 29223
rect 16129 29189 16163 29223
rect 19441 29189 19475 29223
rect 24133 29189 24167 29223
rect 24349 29189 24383 29223
rect 25881 29189 25915 29223
rect 26081 29189 26115 29223
rect 12081 29121 12115 29155
rect 14841 29121 14875 29155
rect 16773 29121 16807 29155
rect 17049 29121 17083 29155
rect 19625 29121 19659 29155
rect 21005 29121 21039 29155
rect 22569 29121 22603 29155
rect 22752 29121 22786 29155
rect 23673 29121 23707 29155
rect 26985 29121 27019 29155
rect 28273 29121 28307 29155
rect 28365 29121 28399 29155
rect 28549 29121 28583 29155
rect 29193 29121 29227 29155
rect 29377 29121 29411 29155
rect 29469 29121 29503 29155
rect 29561 29121 29595 29155
rect 30757 29121 30791 29155
rect 34529 29121 34563 29155
rect 38025 29121 38059 29155
rect 14565 29053 14599 29087
rect 22661 29053 22695 29087
rect 22845 29053 22879 29087
rect 31033 29053 31067 29087
rect 23029 28985 23063 29019
rect 24501 28985 24535 29019
rect 26249 28985 26283 29019
rect 1685 28917 1719 28951
rect 13461 28917 13495 28951
rect 15945 28917 15979 28951
rect 24317 28917 24351 28951
rect 26065 28917 26099 28951
rect 27169 28917 27203 28951
rect 41797 28917 41831 28951
rect 14657 28713 14691 28747
rect 21741 28713 21775 28747
rect 23489 28645 23523 28679
rect 24869 28645 24903 28679
rect 28825 28645 28859 28679
rect 28917 28645 28951 28679
rect 1409 28577 1443 28611
rect 2789 28577 2823 28611
rect 14197 28577 14231 28611
rect 14381 28577 14415 28611
rect 14473 28577 14507 28611
rect 19625 28577 19659 28611
rect 22477 28577 22511 28611
rect 22661 28577 22695 28611
rect 25329 28577 25363 28611
rect 28089 28577 28123 28611
rect 41337 28577 41371 28611
rect 42165 28577 42199 28611
rect 13553 28509 13587 28543
rect 14289 28509 14323 28543
rect 16221 28509 16255 28543
rect 16589 28509 16623 28543
rect 17233 28509 17267 28543
rect 17417 28509 17451 28543
rect 21649 28509 21683 28543
rect 22385 28509 22419 28543
rect 22569 28509 22603 28543
rect 23305 28509 23339 28543
rect 25237 28509 25271 28543
rect 27005 28509 27039 28543
rect 27261 28509 27295 28543
rect 27813 28509 27847 28543
rect 27905 28509 27939 28543
rect 28549 28509 28583 28543
rect 28687 28509 28721 28543
rect 29009 28509 29043 28543
rect 29561 28509 29595 28543
rect 29745 28509 29779 28543
rect 30573 28509 30607 28543
rect 1593 28441 1627 28475
rect 16405 28441 16439 28475
rect 16497 28441 16531 28475
rect 19892 28441 19926 28475
rect 30818 28441 30852 28475
rect 41981 28441 42015 28475
rect 13461 28373 13495 28407
rect 16773 28373 16807 28407
rect 17417 28373 17451 28407
rect 21005 28373 21039 28407
rect 22845 28373 22879 28407
rect 25881 28373 25915 28407
rect 28089 28373 28123 28407
rect 29561 28373 29595 28407
rect 31953 28373 31987 28407
rect 2145 28169 2179 28203
rect 17785 28169 17819 28203
rect 20269 28169 20303 28203
rect 26341 28169 26375 28203
rect 28641 28169 28675 28203
rect 29745 28169 29779 28203
rect 41429 28169 41463 28203
rect 14657 28101 14691 28135
rect 16129 28101 16163 28135
rect 17049 28101 17083 28135
rect 19809 28101 19843 28135
rect 22845 28101 22879 28135
rect 26157 28101 26191 28135
rect 30389 28101 30423 28135
rect 31585 28101 31619 28135
rect 32781 28101 32815 28135
rect 33577 28101 33611 28135
rect 33793 28101 33827 28135
rect 2237 28033 2271 28067
rect 12725 28033 12759 28067
rect 14473 28033 14507 28067
rect 15577 28033 15611 28067
rect 15853 28033 15887 28067
rect 15945 28033 15979 28067
rect 16819 28033 16853 28067
rect 16957 28033 16991 28067
rect 17232 28033 17266 28067
rect 17325 28033 17359 28067
rect 18153 28033 18187 28067
rect 18245 28033 18279 28067
rect 18797 28033 18831 28067
rect 19625 28033 19659 28067
rect 20453 28033 20487 28067
rect 24124 28033 24158 28067
rect 25973 28033 26007 28067
rect 28273 28033 28307 28067
rect 28457 28033 28491 28067
rect 29101 28033 29135 28067
rect 29264 28033 29298 28067
rect 29364 28033 29398 28067
rect 29489 28033 29523 28067
rect 31401 28033 31435 28067
rect 32597 28033 32631 28067
rect 34897 28033 34931 28067
rect 41337 28033 41371 28067
rect 15669 27965 15703 27999
rect 17969 27965 18003 27999
rect 18061 27965 18095 27999
rect 23029 27965 23063 27999
rect 23857 27965 23891 27999
rect 28181 27965 28215 27999
rect 28365 27965 28399 27999
rect 32965 27897 32999 27931
rect 12541 27829 12575 27863
rect 14841 27829 14875 27863
rect 16681 27829 16715 27863
rect 18981 27829 19015 27863
rect 25237 27829 25271 27863
rect 30297 27829 30331 27863
rect 33425 27829 33459 27863
rect 33609 27829 33643 27863
rect 34897 27829 34931 27863
rect 20361 27625 20395 27659
rect 20545 27625 20579 27659
rect 22569 27625 22603 27659
rect 24409 27625 24443 27659
rect 25973 27625 26007 27659
rect 28181 27625 28215 27659
rect 28825 27625 28859 27659
rect 29561 27625 29595 27659
rect 31585 27625 31619 27659
rect 15393 27557 15427 27591
rect 16865 27557 16899 27591
rect 18613 27557 18647 27591
rect 21005 27557 21039 27591
rect 22385 27557 22419 27591
rect 23765 27557 23799 27591
rect 29745 27557 29779 27591
rect 30849 27557 30883 27591
rect 11897 27489 11931 27523
rect 16405 27489 16439 27523
rect 23397 27489 23431 27523
rect 32781 27489 32815 27523
rect 12164 27421 12198 27455
rect 14473 27421 14507 27455
rect 14657 27421 14691 27455
rect 15117 27421 15151 27455
rect 16313 27421 16347 27455
rect 16589 27421 16623 27455
rect 16681 27421 16715 27455
rect 19993 27421 20027 27455
rect 21189 27421 21223 27455
rect 21465 27421 21499 27455
rect 22937 27421 22971 27455
rect 24593 27421 24627 27455
rect 25881 27421 25915 27455
rect 26065 27421 26099 27455
rect 26617 27421 26651 27455
rect 27997 27421 28031 27455
rect 28181 27421 28215 27455
rect 32137 27421 32171 27455
rect 41429 27421 41463 27455
rect 15393 27353 15427 27387
rect 18337 27353 18371 27387
rect 20361 27353 20395 27387
rect 28793 27353 28827 27387
rect 29009 27353 29043 27387
rect 30021 27353 30055 27387
rect 30849 27353 30883 27387
rect 33026 27353 33060 27387
rect 13277 27285 13311 27319
rect 14657 27285 14691 27319
rect 15209 27285 15243 27319
rect 21373 27285 21407 27319
rect 22569 27285 22603 27319
rect 23857 27285 23891 27319
rect 26709 27285 26743 27319
rect 28641 27285 28675 27319
rect 31309 27285 31343 27319
rect 31401 27285 31435 27319
rect 32321 27285 32355 27319
rect 34161 27285 34195 27319
rect 41521 27285 41555 27319
rect 13001 27081 13035 27115
rect 20637 27081 20671 27115
rect 23213 27081 23247 27115
rect 24041 27081 24075 27115
rect 28089 27081 28123 27115
rect 23673 27013 23707 27047
rect 23873 27013 23907 27047
rect 41705 27013 41739 27047
rect 13185 26945 13219 26979
rect 15301 26945 15335 26979
rect 15577 26945 15611 26979
rect 16681 26945 16715 26979
rect 19818 26945 19852 26979
rect 20085 26945 20119 26979
rect 20545 26945 20579 26979
rect 21833 26945 21867 26979
rect 22089 26945 22123 26979
rect 26065 26945 26099 26979
rect 28273 26945 28307 26979
rect 28917 26945 28951 26979
rect 29193 26945 29227 26979
rect 30941 26945 30975 26979
rect 31401 26945 31435 26979
rect 32781 26945 32815 26979
rect 32965 26945 32999 26979
rect 33057 26945 33091 26979
rect 33149 26945 33183 26979
rect 33885 26945 33919 26979
rect 34141 26945 34175 26979
rect 13369 26877 13403 26911
rect 15485 26877 15519 26911
rect 16957 26877 16991 26911
rect 21005 26877 21039 26911
rect 28457 26877 28491 26911
rect 31217 26877 31251 26911
rect 33425 26877 33459 26911
rect 41337 26877 41371 26911
rect 41889 26877 41923 26911
rect 15393 26809 15427 26843
rect 15761 26741 15795 26775
rect 16773 26741 16807 26775
rect 16865 26741 16899 26775
rect 18705 26741 18739 26775
rect 20821 26741 20855 26775
rect 23857 26741 23891 26775
rect 26249 26741 26283 26775
rect 31033 26741 31067 26775
rect 31585 26741 31619 26775
rect 35265 26741 35299 26775
rect 16405 26537 16439 26571
rect 19533 26537 19567 26571
rect 19901 26537 19935 26571
rect 21833 26537 21867 26571
rect 25421 26537 25455 26571
rect 25605 26537 25639 26571
rect 29561 26537 29595 26571
rect 30021 26537 30055 26571
rect 32045 26537 32079 26571
rect 34069 26537 34103 26571
rect 41797 26537 41831 26571
rect 13553 26469 13587 26503
rect 15577 26469 15611 26503
rect 29009 26469 29043 26503
rect 32413 26469 32447 26503
rect 33517 26469 33551 26503
rect 12173 26401 12207 26435
rect 14381 26401 14415 26435
rect 14749 26401 14783 26435
rect 15669 26401 15703 26435
rect 16313 26401 16347 26435
rect 19993 26401 20027 26435
rect 20637 26401 20671 26435
rect 23397 26401 23431 26435
rect 26065 26401 26099 26435
rect 28365 26401 28399 26435
rect 29837 26401 29871 26435
rect 31033 26401 31067 26435
rect 14289 26333 14323 26367
rect 15393 26333 15427 26367
rect 16497 26333 16531 26367
rect 16589 26333 16623 26367
rect 17233 26333 17267 26367
rect 19717 26333 19751 26367
rect 20545 26333 20579 26367
rect 20729 26333 20763 26367
rect 21189 26333 21223 26367
rect 21373 26333 21407 26367
rect 21468 26333 21502 26367
rect 21603 26333 21637 26367
rect 23121 26333 23155 26367
rect 24593 26333 24627 26367
rect 25053 26333 25087 26367
rect 26332 26333 26366 26367
rect 28641 26333 28675 26367
rect 28850 26333 28884 26367
rect 30113 26333 30147 26367
rect 30757 26333 30791 26367
rect 32045 26333 32079 26367
rect 32229 26333 32263 26367
rect 33316 26333 33350 26367
rect 33977 26333 34011 26367
rect 34161 26333 34195 26367
rect 34897 26333 34931 26367
rect 12440 26265 12474 26299
rect 14105 26265 14139 26299
rect 17141 26265 17175 26299
rect 34805 26265 34839 26299
rect 15209 26197 15243 26231
rect 24409 26197 24443 26231
rect 25421 26197 25455 26231
rect 27445 26197 27479 26231
rect 28733 26197 28767 26231
rect 14381 25993 14415 26027
rect 15485 25993 15519 26027
rect 20821 25993 20855 26027
rect 20984 25993 21018 26027
rect 25513 25993 25547 26027
rect 28641 25993 28675 26027
rect 29009 25993 29043 26027
rect 31033 25993 31067 26027
rect 32505 25993 32539 26027
rect 33885 25993 33919 26027
rect 21189 25925 21223 25959
rect 23940 25925 23974 25959
rect 25881 25925 25915 25959
rect 14565 25857 14599 25891
rect 14749 25857 14783 25891
rect 15393 25857 15427 25891
rect 15669 25857 15703 25891
rect 18438 25857 18472 25891
rect 18705 25857 18739 25891
rect 23029 25857 23063 25891
rect 23673 25857 23707 25891
rect 25697 25857 25731 25891
rect 25973 25857 26007 25891
rect 27353 25857 27387 25891
rect 28549 25857 28583 25891
rect 28825 25857 28859 25891
rect 29909 25857 29943 25891
rect 32321 25857 32355 25891
rect 33885 25857 33919 25891
rect 34069 25857 34103 25891
rect 14841 25789 14875 25823
rect 27261 25789 27295 25823
rect 29653 25789 29687 25823
rect 32137 25789 32171 25823
rect 15853 25721 15887 25755
rect 25053 25721 25087 25755
rect 17325 25653 17359 25687
rect 21005 25653 21039 25687
rect 23121 25653 23155 25687
rect 26985 25653 27019 25687
rect 27169 25653 27203 25687
rect 41797 25653 41831 25687
rect 15209 25449 15243 25483
rect 15393 25449 15427 25483
rect 24409 25449 24443 25483
rect 25513 25449 25547 25483
rect 28917 25449 28951 25483
rect 30113 25449 30147 25483
rect 16221 25313 16255 25347
rect 17601 25313 17635 25347
rect 24568 25313 24602 25347
rect 24685 25313 24719 25347
rect 25053 25313 25087 25347
rect 25881 25313 25915 25347
rect 26617 25313 26651 25347
rect 26893 25313 26927 25347
rect 31401 25313 31435 25347
rect 14565 25245 14599 25279
rect 15393 25245 15427 25279
rect 15577 25245 15611 25279
rect 16497 25245 16531 25279
rect 17877 25245 17911 25279
rect 20177 25245 20211 25279
rect 20361 25245 20395 25279
rect 25697 25245 25731 25279
rect 28549 25245 28583 25279
rect 30389 25245 30423 25279
rect 30573 25245 30607 25279
rect 31309 25245 31343 25279
rect 31585 25245 31619 25279
rect 32413 25245 32447 25279
rect 32689 25245 32723 25279
rect 33333 25245 33367 25279
rect 33517 25245 33551 25279
rect 40509 25245 40543 25279
rect 41337 25245 41371 25279
rect 41797 25245 41831 25279
rect 14657 25177 14691 25211
rect 28733 25177 28767 25211
rect 32505 25177 32539 25211
rect 41889 25177 41923 25211
rect 20269 25109 20303 25143
rect 24777 25109 24811 25143
rect 30297 25109 30331 25143
rect 31769 25109 31803 25143
rect 32873 25109 32907 25143
rect 33333 25109 33367 25143
rect 41245 25109 41279 25143
rect 14289 24905 14323 24939
rect 25681 24905 25715 24939
rect 27353 24905 27387 24939
rect 28641 24905 28675 24939
rect 29561 24905 29595 24939
rect 31417 24905 31451 24939
rect 15669 24837 15703 24871
rect 15879 24837 15913 24871
rect 25881 24837 25915 24871
rect 27261 24837 27295 24871
rect 31217 24837 31251 24871
rect 40233 24837 40267 24871
rect 12909 24769 12943 24803
rect 13176 24769 13210 24803
rect 14933 24769 14967 24803
rect 15577 24769 15611 24803
rect 15761 24769 15795 24803
rect 16037 24769 16071 24803
rect 17049 24769 17083 24803
rect 17417 24769 17451 24803
rect 19533 24769 19567 24803
rect 19789 24769 19823 24803
rect 22201 24769 22235 24803
rect 23029 24769 23063 24803
rect 27169 24769 27203 24803
rect 28825 24769 28859 24803
rect 29377 24769 29411 24803
rect 32321 24769 32355 24803
rect 32505 24772 32539 24806
rect 32600 24769 32634 24803
rect 32689 24769 32723 24803
rect 34538 24769 34572 24803
rect 34805 24769 34839 24803
rect 36378 24769 36412 24803
rect 36645 24769 36679 24803
rect 39313 24769 39347 24803
rect 40049 24769 40083 24803
rect 14841 24701 14875 24735
rect 17325 24701 17359 24735
rect 22293 24701 22327 24735
rect 26985 24701 27019 24735
rect 32965 24701 32999 24735
rect 41245 24701 41279 24735
rect 15393 24633 15427 24667
rect 17509 24633 17543 24667
rect 25513 24633 25547 24667
rect 27537 24633 27571 24667
rect 17141 24565 17175 24599
rect 20913 24565 20947 24599
rect 22569 24565 22603 24599
rect 23213 24565 23247 24599
rect 25697 24565 25731 24599
rect 31401 24565 31435 24599
rect 31585 24565 31619 24599
rect 33425 24565 33459 24599
rect 35265 24565 35299 24599
rect 39497 24565 39531 24599
rect 13461 24361 13495 24395
rect 15025 24361 15059 24395
rect 15577 24361 15611 24395
rect 17141 24361 17175 24395
rect 19625 24361 19659 24395
rect 20821 24361 20855 24395
rect 23397 24361 23431 24395
rect 29745 24361 29779 24395
rect 30573 24361 30607 24395
rect 31493 24361 31527 24395
rect 32689 24361 32723 24395
rect 33333 24361 33367 24395
rect 34161 24361 34195 24395
rect 21557 24293 21591 24327
rect 26249 24293 26283 24327
rect 29009 24293 29043 24327
rect 32321 24293 32355 24327
rect 32873 24293 32907 24327
rect 37565 24293 37599 24327
rect 3801 24225 3835 24259
rect 5641 24225 5675 24259
rect 14841 24225 14875 24259
rect 17233 24225 17267 24259
rect 18429 24225 18463 24259
rect 21005 24225 21039 24259
rect 23765 24225 23799 24259
rect 24685 24225 24719 24259
rect 26801 24225 26835 24259
rect 31585 24225 31619 24259
rect 40049 24225 40083 24259
rect 40509 24225 40543 24259
rect 13369 24157 13403 24191
rect 13553 24157 13587 24191
rect 14105 24157 14139 24191
rect 14197 24157 14231 24191
rect 15117 24157 15151 24191
rect 15945 24157 15979 24191
rect 16957 24157 16991 24191
rect 17049 24157 17083 24191
rect 18245 24157 18279 24191
rect 19901 24157 19935 24191
rect 19993 24157 20027 24191
rect 20085 24157 20119 24191
rect 20269 24157 20303 24191
rect 22109 24157 22143 24191
rect 22385 24157 22419 24191
rect 23581 24157 23615 24191
rect 24409 24157 24443 24191
rect 24501 24157 24535 24191
rect 26065 24157 26099 24191
rect 26709 24157 26743 24191
rect 28733 24157 28767 24191
rect 28825 24157 28859 24191
rect 30481 24157 30515 24191
rect 30665 24157 30699 24191
rect 31309 24157 31343 24191
rect 33517 24157 33551 24191
rect 33977 24157 34011 24191
rect 37749 24157 37783 24191
rect 39129 24157 39163 24191
rect 5457 24089 5491 24123
rect 14381 24089 14415 24123
rect 14841 24089 14875 24123
rect 15761 24089 15795 24123
rect 21557 24089 21591 24123
rect 29009 24089 29043 24123
rect 29561 24089 29595 24123
rect 32689 24089 32723 24123
rect 39221 24089 39255 24123
rect 40233 24089 40267 24123
rect 14289 24021 14323 24055
rect 18061 24021 18095 24055
rect 21097 24021 21131 24055
rect 24685 24021 24719 24055
rect 29761 24021 29795 24055
rect 29929 24021 29963 24055
rect 31125 24021 31159 24055
rect 3433 23817 3467 23851
rect 16773 23817 16807 23851
rect 20729 23817 20763 23851
rect 22201 23817 22235 23851
rect 24501 23817 24535 23851
rect 25605 23817 25639 23851
rect 29745 23817 29779 23851
rect 32321 23817 32355 23851
rect 23366 23749 23400 23783
rect 3341 23681 3375 23715
rect 14637 23681 14671 23715
rect 16865 23681 16899 23715
rect 17684 23681 17718 23715
rect 19441 23681 19475 23715
rect 20913 23681 20947 23715
rect 21005 23681 21039 23715
rect 24961 23681 24995 23715
rect 25145 23681 25179 23715
rect 25421 23681 25455 23715
rect 26065 23681 26099 23715
rect 26433 23681 26467 23715
rect 26985 23681 27019 23715
rect 27169 23681 27203 23715
rect 27537 23681 27571 23715
rect 28181 23681 28215 23715
rect 28344 23687 28378 23721
rect 28444 23681 28478 23715
rect 28549 23681 28583 23715
rect 29285 23681 29319 23715
rect 29748 23681 29782 23715
rect 30665 23681 30699 23715
rect 30757 23681 30791 23715
rect 32137 23681 32171 23715
rect 32229 23681 32263 23715
rect 35265 23681 35299 23715
rect 35521 23681 35555 23715
rect 37749 23681 37783 23715
rect 38016 23681 38050 23715
rect 41889 23681 41923 23715
rect 14381 23613 14415 23647
rect 17417 23613 17451 23647
rect 19533 23613 19567 23647
rect 21097 23613 21131 23647
rect 21189 23613 21223 23647
rect 22293 23613 22327 23647
rect 22477 23613 22511 23647
rect 23121 23613 23155 23647
rect 26249 23613 26283 23647
rect 27261 23613 27295 23647
rect 27353 23613 27387 23647
rect 27721 23613 27755 23647
rect 30573 23613 30607 23647
rect 30849 23613 30883 23647
rect 32597 23613 32631 23647
rect 41337 23613 41371 23647
rect 41705 23613 41739 23647
rect 15761 23545 15795 23579
rect 18797 23545 18831 23579
rect 19809 23545 19843 23579
rect 21833 23477 21867 23511
rect 26249 23477 26283 23511
rect 26341 23477 26375 23511
rect 28825 23477 28859 23511
rect 29377 23477 29411 23511
rect 29929 23477 29963 23511
rect 30389 23477 30423 23511
rect 39129 23477 39163 23511
rect 19441 23273 19475 23307
rect 20821 23273 20855 23307
rect 23857 23273 23891 23307
rect 26893 23273 26927 23307
rect 32229 23273 32263 23307
rect 38669 23273 38703 23307
rect 38209 23205 38243 23239
rect 17877 23137 17911 23171
rect 23397 23137 23431 23171
rect 24409 23137 24443 23171
rect 24685 23137 24719 23171
rect 29561 23137 29595 23171
rect 30113 23137 30147 23171
rect 30849 23137 30883 23171
rect 34897 23137 34931 23171
rect 39037 23137 39071 23171
rect 40509 23137 40543 23171
rect 40785 23137 40819 23171
rect 1685 23069 1719 23103
rect 18153 23069 18187 23103
rect 19625 23069 19659 23103
rect 19809 23069 19843 23103
rect 19993 23069 20027 23103
rect 20821 23069 20855 23103
rect 21097 23069 21131 23103
rect 22477 23069 22511 23103
rect 23305 23069 23339 23103
rect 23581 23069 23615 23103
rect 23673 23069 23707 23103
rect 28181 23069 28215 23103
rect 29745 23069 29779 23103
rect 31116 23069 31150 23103
rect 36829 23069 36863 23103
rect 38853 23069 38887 23103
rect 40325 23069 40359 23103
rect 19717 23001 19751 23035
rect 20913 23001 20947 23035
rect 22569 23001 22603 23035
rect 28733 23001 28767 23035
rect 30021 23001 30055 23035
rect 35142 23001 35176 23035
rect 37096 23001 37130 23035
rect 28825 22933 28859 22967
rect 17877 22729 17911 22763
rect 25973 22729 26007 22763
rect 38301 22729 38335 22763
rect 28181 22661 28215 22695
rect 2145 22593 2179 22627
rect 18061 22593 18095 22627
rect 18613 22593 18647 22627
rect 22661 22593 22695 22627
rect 23489 22593 23523 22627
rect 23765 22593 23799 22627
rect 23857 22593 23891 22627
rect 25513 22593 25547 22627
rect 25605 22593 25639 22627
rect 25789 22593 25823 22627
rect 26985 22593 27019 22627
rect 27169 22593 27203 22627
rect 27537 22593 27571 22627
rect 28365 22593 28399 22627
rect 28457 22593 28491 22627
rect 29101 22593 29135 22627
rect 29193 22593 29227 22627
rect 29469 22593 29503 22627
rect 30113 22593 30147 22627
rect 30297 22593 30331 22627
rect 32137 22593 32171 22627
rect 32321 22593 32355 22627
rect 32413 22593 32447 22627
rect 34906 22593 34940 22627
rect 35173 22593 35207 22627
rect 38117 22593 38151 22627
rect 38761 22593 38795 22627
rect 39017 22593 39051 22627
rect 40785 22593 40819 22627
rect 41429 22593 41463 22627
rect 22937 22525 22971 22559
rect 27261 22525 27295 22559
rect 27353 22525 27387 22559
rect 40969 22525 41003 22559
rect 23581 22457 23615 22491
rect 24041 22457 24075 22491
rect 27721 22457 27755 22491
rect 40141 22457 40175 22491
rect 2053 22389 2087 22423
rect 18797 22389 18831 22423
rect 28181 22389 28215 22423
rect 28917 22389 28951 22423
rect 29377 22389 29411 22423
rect 29929 22389 29963 22423
rect 32137 22389 32171 22423
rect 40601 22389 40635 22423
rect 41521 22389 41555 22423
rect 18245 22185 18279 22219
rect 20821 22185 20855 22219
rect 22753 22185 22787 22219
rect 24501 22185 24535 22219
rect 26709 22185 26743 22219
rect 29745 22185 29779 22219
rect 29837 22185 29871 22219
rect 31953 22185 31987 22219
rect 20729 22117 20763 22151
rect 25605 22117 25639 22151
rect 28733 22117 28767 22151
rect 32045 22117 32079 22151
rect 1409 22049 1443 22083
rect 1593 22049 1627 22083
rect 1869 22049 1903 22083
rect 15945 22049 15979 22083
rect 16221 22049 16255 22083
rect 20637 22049 20671 22083
rect 27813 22049 27847 22083
rect 29745 22049 29779 22083
rect 30481 22049 30515 22083
rect 31861 22049 31895 22083
rect 34713 22049 34747 22083
rect 39313 22049 39347 22083
rect 40509 22049 40543 22083
rect 42165 22049 42199 22083
rect 15485 21981 15519 22015
rect 16313 21981 16347 22015
rect 17969 21981 18003 22015
rect 18061 21981 18095 22015
rect 19809 21981 19843 22015
rect 20913 21981 20947 22015
rect 21373 21981 21407 22015
rect 24409 21981 24443 22015
rect 24593 21981 24627 22015
rect 25789 21981 25823 22015
rect 27077 21981 27111 22015
rect 28630 21981 28664 22015
rect 28917 21981 28951 22015
rect 29929 21981 29963 22015
rect 30389 21981 30423 22015
rect 32137 21981 32171 22015
rect 32781 21981 32815 22015
rect 33037 21981 33071 22015
rect 34989 21981 35023 22015
rect 36001 21981 36035 22015
rect 36185 21981 36219 22015
rect 39037 21981 39071 22015
rect 39129 21981 39163 22015
rect 40325 21981 40359 22015
rect 15240 21913 15274 21947
rect 21640 21913 21674 21947
rect 25973 21913 26007 21947
rect 26893 21913 26927 21947
rect 27629 21913 27663 21947
rect 29561 21913 29595 21947
rect 14105 21845 14139 21879
rect 19717 21845 19751 21879
rect 28641 21845 28675 21879
rect 34161 21845 34195 21879
rect 36369 21845 36403 21879
rect 14657 21641 14691 21675
rect 22017 21641 22051 21675
rect 22937 21641 22971 21675
rect 24041 21641 24075 21675
rect 25421 21641 25455 21675
rect 26065 21641 26099 21675
rect 29745 21641 29779 21675
rect 32305 21641 32339 21675
rect 38669 21641 38703 21675
rect 19226 21573 19260 21607
rect 21833 21573 21867 21607
rect 32505 21573 32539 21607
rect 35633 21573 35667 21607
rect 41889 21573 41923 21607
rect 6377 21505 6411 21539
rect 14749 21505 14783 21539
rect 15301 21505 15335 21539
rect 16681 21505 16715 21539
rect 16948 21505 16982 21539
rect 18981 21505 19015 21539
rect 22109 21505 22143 21539
rect 22753 21505 22787 21539
rect 24317 21505 24351 21539
rect 24593 21505 24627 21539
rect 25053 21505 25087 21539
rect 25973 21505 26007 21539
rect 27353 21505 27387 21539
rect 27537 21505 27571 21539
rect 28549 21505 28583 21539
rect 28733 21505 28767 21539
rect 29285 21505 29319 21539
rect 29561 21505 29595 21539
rect 35541 21505 35575 21539
rect 35725 21505 35759 21539
rect 36185 21505 36219 21539
rect 36369 21505 36403 21539
rect 38485 21505 38519 21539
rect 39589 21505 39623 21539
rect 1869 21437 1903 21471
rect 2053 21437 2087 21471
rect 2789 21437 2823 21471
rect 7113 21437 7147 21471
rect 15577 21437 15611 21471
rect 24133 21437 24167 21471
rect 25145 21437 25179 21471
rect 27721 21437 27755 21471
rect 37565 21437 37599 21471
rect 38025 21437 38059 21471
rect 40049 21437 40083 21471
rect 40233 21437 40267 21471
rect 21833 21369 21867 21403
rect 29377 21369 29411 21403
rect 29469 21369 29503 21403
rect 32137 21369 32171 21403
rect 37933 21369 37967 21403
rect 18061 21301 18095 21335
rect 20361 21301 20395 21335
rect 25145 21301 25179 21335
rect 28733 21301 28767 21335
rect 32321 21301 32355 21335
rect 36185 21301 36219 21335
rect 1961 21097 1995 21131
rect 2697 21097 2731 21131
rect 7481 21097 7515 21131
rect 15485 21097 15519 21131
rect 17233 21097 17267 21131
rect 20821 21097 20855 21131
rect 28917 21097 28951 21131
rect 31033 21097 31067 21131
rect 37197 21097 37231 21131
rect 38117 21097 38151 21131
rect 39313 21097 39347 21131
rect 40969 21097 41003 21131
rect 41613 21097 41647 21131
rect 17693 21029 17727 21063
rect 27077 21029 27111 21063
rect 30665 21029 30699 21063
rect 33057 21029 33091 21063
rect 36277 21029 36311 21063
rect 13461 20961 13495 20995
rect 16129 20961 16163 20995
rect 20913 20961 20947 20995
rect 25513 20961 25547 20995
rect 33701 20961 33735 20995
rect 36001 20961 36035 20995
rect 36829 20961 36863 20995
rect 37013 20961 37047 20995
rect 2789 20893 2823 20927
rect 5733 20893 5767 20927
rect 6193 20893 6227 20927
rect 13369 20893 13403 20927
rect 13553 20893 13587 20927
rect 14381 20893 14415 20927
rect 14473 20893 14507 20927
rect 14565 20893 14599 20927
rect 14749 20893 14783 20927
rect 15669 20893 15703 20927
rect 16589 20893 16623 20927
rect 16864 20893 16898 20927
rect 17049 20893 17083 20927
rect 17969 20893 18003 20927
rect 19257 20893 19291 20927
rect 19441 20893 19475 20927
rect 19625 20893 19659 20927
rect 20269 20893 20303 20927
rect 21097 20893 21131 20927
rect 21925 20893 21959 20927
rect 24593 20893 24627 20927
rect 25237 20893 25271 20927
rect 27077 20893 27111 20927
rect 27261 20893 27295 20927
rect 27905 20893 27939 20927
rect 28733 20893 28767 20927
rect 28917 20893 28951 20927
rect 31677 20893 31711 20927
rect 33793 20893 33827 20927
rect 34713 20893 34747 20927
rect 34989 20893 35023 20927
rect 35081 20893 35115 20927
rect 35909 20893 35943 20927
rect 36921 20893 36955 20927
rect 37657 20893 37691 20927
rect 37749 20893 37783 20927
rect 37933 20893 37967 20927
rect 39129 20893 39163 20927
rect 40049 20893 40083 20927
rect 40233 20893 40267 20927
rect 40325 20893 40359 20927
rect 40877 20893 40911 20927
rect 41521 20893 41555 20927
rect 5457 20825 5491 20859
rect 15761 20825 15795 20859
rect 15853 20825 15887 20859
rect 15991 20825 16025 20859
rect 16727 20825 16761 20859
rect 16957 20825 16991 20859
rect 17693 20825 17727 20859
rect 17877 20825 17911 20859
rect 20821 20825 20855 20859
rect 24777 20825 24811 20859
rect 26709 20825 26743 20859
rect 27721 20825 27755 20859
rect 28089 20825 28123 20859
rect 31033 20825 31067 20859
rect 31922 20825 31956 20859
rect 34897 20825 34931 20859
rect 14105 20757 14139 20791
rect 20085 20757 20119 20791
rect 21281 20757 21315 20791
rect 21833 20757 21867 20791
rect 31217 20757 31251 20791
rect 34161 20757 34195 20791
rect 35265 20757 35299 20791
rect 5733 20553 5767 20587
rect 16957 20553 16991 20587
rect 21005 20553 21039 20587
rect 24225 20553 24259 20587
rect 24777 20553 24811 20587
rect 27537 20553 27571 20587
rect 28733 20553 28767 20587
rect 30021 20553 30055 20587
rect 31585 20553 31619 20587
rect 32137 20553 32171 20587
rect 32505 20553 32539 20587
rect 33977 20553 34011 20587
rect 40233 20553 40267 20587
rect 13176 20485 13210 20519
rect 14841 20485 14875 20519
rect 19892 20485 19926 20519
rect 25237 20485 25271 20519
rect 27077 20485 27111 20519
rect 36277 20485 36311 20519
rect 38393 20485 38427 20519
rect 39098 20485 39132 20519
rect 15071 20451 15105 20485
rect 5549 20417 5583 20451
rect 6377 20417 6411 20451
rect 15669 20417 15703 20451
rect 16865 20417 16899 20451
rect 17049 20417 17083 20451
rect 18705 20417 18739 20451
rect 24133 20417 24167 20451
rect 24317 20417 24351 20451
rect 24961 20417 24995 20451
rect 26249 20417 26283 20451
rect 28181 20417 28215 20451
rect 28549 20417 28583 20451
rect 29929 20417 29963 20451
rect 30757 20417 30791 20451
rect 30941 20417 30975 20451
rect 31401 20417 31435 20451
rect 32321 20417 32355 20451
rect 32597 20417 32631 20451
rect 33885 20417 33919 20451
rect 34069 20417 34103 20451
rect 37749 20417 37783 20451
rect 37933 20417 37967 20451
rect 38209 20417 38243 20451
rect 40969 20417 41003 20451
rect 41613 20417 41647 20451
rect 7205 20349 7239 20383
rect 12909 20349 12943 20383
rect 15761 20349 15795 20383
rect 18521 20349 18555 20383
rect 19625 20349 19659 20383
rect 25145 20349 25179 20383
rect 30113 20349 30147 20383
rect 38853 20349 38887 20383
rect 14289 20281 14323 20315
rect 15209 20281 15243 20315
rect 27445 20281 27479 20315
rect 36645 20281 36679 20315
rect 1685 20213 1719 20247
rect 15025 20213 15059 20247
rect 15853 20213 15887 20247
rect 16037 20213 16071 20247
rect 18889 20213 18923 20247
rect 25237 20213 25271 20247
rect 26433 20213 26467 20247
rect 28549 20213 28583 20247
rect 29561 20213 29595 20247
rect 30757 20213 30791 20247
rect 36737 20213 36771 20247
rect 41061 20213 41095 20247
rect 41705 20213 41739 20247
rect 18429 19941 18463 19975
rect 20729 19941 20763 19975
rect 24501 19941 24535 19975
rect 30389 19941 30423 19975
rect 32505 19941 32539 19975
rect 1409 19873 1443 19907
rect 1869 19873 1903 19907
rect 6745 19873 6779 19907
rect 11621 19873 11655 19907
rect 15761 19873 15795 19907
rect 24869 19873 24903 19907
rect 25513 19873 25547 19907
rect 25789 19873 25823 19907
rect 27077 19873 27111 19907
rect 27353 19873 27387 19907
rect 28089 19873 28123 19907
rect 34805 19873 34839 19907
rect 36911 19873 36945 19907
rect 38577 19873 38611 19907
rect 40509 19873 40543 19907
rect 6193 19805 6227 19839
rect 10333 19805 10367 19839
rect 10517 19805 10551 19839
rect 11069 19805 11103 19839
rect 16037 19805 16071 19839
rect 19349 19805 19383 19839
rect 21741 19805 21775 19839
rect 22385 19805 22419 19839
rect 24685 19805 24719 19839
rect 24777 19805 24811 19839
rect 24961 19805 24995 19839
rect 26985 19805 27019 19839
rect 27905 19805 27939 19839
rect 30113 19805 30147 19839
rect 30205 19805 30239 19839
rect 30389 19805 30423 19839
rect 32321 19805 32355 19839
rect 32597 19805 32631 19839
rect 34897 19805 34931 19839
rect 36829 19805 36863 19839
rect 37013 19805 37047 19839
rect 37565 19805 37599 19839
rect 37841 19805 37875 19839
rect 38485 19805 38519 19839
rect 38669 19805 38703 19839
rect 39129 19805 39163 19839
rect 40325 19805 40359 19839
rect 1593 19737 1627 19771
rect 18613 19737 18647 19771
rect 19616 19737 19650 19771
rect 21925 19737 21959 19771
rect 22652 19737 22686 19771
rect 37657 19737 37691 19771
rect 42165 19737 42199 19771
rect 23765 19669 23799 19703
rect 32137 19669 32171 19703
rect 35265 19669 35299 19703
rect 36645 19669 36679 19703
rect 38025 19669 38059 19703
rect 39221 19669 39255 19703
rect 2053 19465 2087 19499
rect 19625 19465 19659 19499
rect 23765 19465 23799 19499
rect 24317 19465 24351 19499
rect 25237 19465 25271 19499
rect 27077 19465 27111 19499
rect 32413 19465 32447 19499
rect 37657 19465 37691 19499
rect 11989 19397 12023 19431
rect 15761 19397 15795 19431
rect 15853 19397 15887 19431
rect 15991 19397 16025 19431
rect 32505 19397 32539 19431
rect 40233 19397 40267 19431
rect 2145 19329 2179 19363
rect 10517 19329 10551 19363
rect 10793 19329 10827 19363
rect 11621 19329 11655 19363
rect 12909 19329 12943 19363
rect 13176 19329 13210 19363
rect 15485 19329 15519 19363
rect 15669 19329 15703 19363
rect 16129 19329 16163 19363
rect 16865 19329 16899 19363
rect 17792 19329 17826 19363
rect 18052 19329 18086 19363
rect 19809 19329 19843 19363
rect 22385 19329 22419 19363
rect 22641 19329 22675 19363
rect 24225 19329 24259 19363
rect 24501 19329 24535 19363
rect 25145 19329 25179 19363
rect 25789 19329 25823 19363
rect 25973 19329 26007 19363
rect 27169 19329 27203 19363
rect 28733 19329 28767 19363
rect 29193 19329 29227 19363
rect 29837 19329 29871 19363
rect 30021 19329 30055 19363
rect 32597 19329 32631 19363
rect 34897 19329 34931 19363
rect 37473 19329 37507 19363
rect 40049 19329 40083 19363
rect 16681 19261 16715 19295
rect 24593 19261 24627 19295
rect 28917 19261 28951 19295
rect 30113 19261 30147 19295
rect 32137 19261 32171 19295
rect 34989 19261 35023 19295
rect 41245 19261 41279 19295
rect 25789 19193 25823 19227
rect 29055 19193 29089 19227
rect 35265 19193 35299 19227
rect 39589 19193 39623 19227
rect 14289 19125 14323 19159
rect 17049 19125 17083 19159
rect 19165 19125 19199 19159
rect 24409 19125 24443 19159
rect 28825 19125 28859 19159
rect 29653 19125 29687 19159
rect 17969 18921 18003 18955
rect 20269 18921 20303 18955
rect 33609 18921 33643 18955
rect 13553 18853 13587 18887
rect 19625 18853 19659 18887
rect 22753 18853 22787 18887
rect 25789 18853 25823 18887
rect 14565 18785 14599 18819
rect 15393 18785 15427 18819
rect 15669 18785 15703 18819
rect 24409 18785 24443 18819
rect 29745 18785 29779 18819
rect 30205 18785 30239 18819
rect 40417 18785 40451 18819
rect 11069 18717 11103 18751
rect 14749 18717 14783 18751
rect 16957 18717 16991 18751
rect 17417 18717 17451 18751
rect 17785 18717 17819 18751
rect 20913 18717 20947 18751
rect 22937 18717 22971 18751
rect 28641 18717 28675 18751
rect 29837 18717 29871 18751
rect 30665 18717 30699 18751
rect 30849 18717 30883 18751
rect 32229 18717 32263 18751
rect 32496 18717 32530 18751
rect 38945 18717 38979 18751
rect 39037 18717 39071 18751
rect 40233 18717 40267 18751
rect 11621 18649 11655 18683
rect 13369 18649 13403 18683
rect 16681 18649 16715 18683
rect 17601 18649 17635 18683
rect 17693 18649 17727 18683
rect 19257 18649 19291 18683
rect 20361 18649 20395 18683
rect 21158 18649 21192 18683
rect 24654 18649 24688 18683
rect 28825 18649 28859 18683
rect 30113 18649 30147 18683
rect 42073 18649 42107 18683
rect 14933 18581 14967 18615
rect 19717 18581 19751 18615
rect 22293 18581 22327 18615
rect 29009 18581 29043 18615
rect 29561 18581 29595 18615
rect 30757 18581 30791 18615
rect 39221 18581 39255 18615
rect 22293 18377 22327 18411
rect 28641 18377 28675 18411
rect 38945 18377 38979 18411
rect 39589 18377 39623 18411
rect 16129 18309 16163 18343
rect 17601 18309 17635 18343
rect 29461 18309 29495 18343
rect 32229 18309 32263 18343
rect 32413 18309 32447 18343
rect 37832 18309 37866 18343
rect 11796 18241 11830 18275
rect 15209 18241 15243 18275
rect 15856 18241 15890 18275
rect 15945 18241 15979 18275
rect 16681 18241 16715 18275
rect 16865 18241 16899 18275
rect 17509 18241 17543 18275
rect 17693 18241 17727 18275
rect 18613 18241 18647 18275
rect 18889 18241 18923 18275
rect 19993 18241 20027 18275
rect 28733 18241 28767 18275
rect 29193 18241 29227 18275
rect 29377 18241 29411 18275
rect 29607 18241 29641 18275
rect 30665 18241 30699 18275
rect 33425 18241 33459 18275
rect 33681 18241 33715 18275
rect 37565 18241 37599 18275
rect 39405 18241 39439 18275
rect 11529 18173 11563 18207
rect 14473 18173 14507 18207
rect 14933 18173 14967 18207
rect 15025 18173 15059 18207
rect 21833 18173 21867 18207
rect 30573 18173 30607 18207
rect 41337 18173 41371 18207
rect 41705 18173 41739 18207
rect 41889 18173 41923 18207
rect 12909 18105 12943 18139
rect 16129 18105 16163 18139
rect 22201 18105 22235 18139
rect 14243 18037 14277 18071
rect 15393 18037 15427 18071
rect 17049 18037 17083 18071
rect 20177 18037 20211 18071
rect 29745 18037 29779 18071
rect 31033 18037 31067 18071
rect 34805 18037 34839 18071
rect 14105 17833 14139 17867
rect 15209 17833 15243 17867
rect 15393 17833 15427 17867
rect 16681 17833 16715 17867
rect 16865 17833 16899 17867
rect 40693 17833 40727 17867
rect 41429 17833 41463 17867
rect 41981 17833 42015 17867
rect 13553 17765 13587 17799
rect 19349 17765 19383 17799
rect 30757 17765 30791 17799
rect 19257 17697 19291 17731
rect 29009 17697 29043 17731
rect 31309 17697 31343 17731
rect 36369 17697 36403 17731
rect 2053 17629 2087 17663
rect 2973 17629 3007 17663
rect 11069 17629 11103 17663
rect 11529 17629 11563 17663
rect 13277 17629 13311 17663
rect 14289 17629 14323 17663
rect 14381 17629 14415 17663
rect 14749 17629 14783 17663
rect 17785 17629 17819 17663
rect 17877 17629 17911 17663
rect 18061 17629 18095 17663
rect 18153 17629 18187 17663
rect 19533 17629 19567 17663
rect 20269 17629 20303 17663
rect 22477 17629 22511 17663
rect 27169 17629 27203 17663
rect 28742 17629 28776 17663
rect 30665 17629 30699 17663
rect 31565 17629 31599 17663
rect 34805 17629 34839 17663
rect 34989 17629 35023 17663
rect 36636 17629 36670 17663
rect 38485 17629 38519 17663
rect 38761 17629 38795 17663
rect 41337 17629 41371 17663
rect 15347 17595 15381 17629
rect 13553 17561 13587 17595
rect 14473 17561 14507 17595
rect 14591 17561 14625 17595
rect 15577 17561 15611 17595
rect 16497 17561 16531 17595
rect 16697 17561 16731 17595
rect 20514 17561 20548 17595
rect 22722 17561 22756 17595
rect 26902 17561 26936 17595
rect 30021 17561 30055 17595
rect 2881 17493 2915 17527
rect 13369 17493 13403 17527
rect 17601 17493 17635 17527
rect 19717 17493 19751 17527
rect 21649 17493 21683 17527
rect 23857 17493 23891 17527
rect 25789 17493 25823 17527
rect 27629 17493 27663 17527
rect 30113 17493 30147 17527
rect 32689 17493 32723 17527
rect 34897 17493 34931 17527
rect 37749 17493 37783 17527
rect 14565 17289 14599 17323
rect 18981 17289 19015 17323
rect 2145 17221 2179 17255
rect 13737 17221 13771 17255
rect 15209 17221 15243 17255
rect 29644 17221 29678 17255
rect 1961 17153 1995 17187
rect 11529 17153 11563 17187
rect 11796 17153 11830 17187
rect 13369 17153 13403 17187
rect 13553 17153 13587 17187
rect 13645 17153 13679 17187
rect 13855 17153 13889 17187
rect 14013 17153 14047 17187
rect 14473 17153 14507 17187
rect 14657 17153 14691 17187
rect 15485 17153 15519 17187
rect 17233 17153 17267 17187
rect 18061 17153 18095 17187
rect 18889 17153 18923 17187
rect 19073 17153 19107 17187
rect 20361 17153 20395 17187
rect 21833 17153 21867 17187
rect 22733 17153 22767 17187
rect 25421 17153 25455 17187
rect 25605 17153 25639 17187
rect 29377 17153 29411 17187
rect 34805 17153 34839 17187
rect 34897 17153 34931 17187
rect 37841 17153 37875 17187
rect 37933 17153 37967 17187
rect 2789 17085 2823 17119
rect 15393 17085 15427 17119
rect 16957 17085 16991 17119
rect 18153 17085 18187 17119
rect 20637 17085 20671 17119
rect 22477 17085 22511 17119
rect 26433 17085 26467 17119
rect 22017 17017 22051 17051
rect 12909 16949 12943 16983
rect 15209 16949 15243 16983
rect 15669 16949 15703 16983
rect 16681 16949 16715 16983
rect 17141 16949 17175 16983
rect 18061 16949 18095 16983
rect 18429 16949 18463 16983
rect 23857 16949 23891 16983
rect 30757 16949 30791 16983
rect 34621 16949 34655 16983
rect 37657 16949 37691 16983
rect 41797 16949 41831 16983
rect 15117 16745 15151 16779
rect 16313 16745 16347 16779
rect 17877 16745 17911 16779
rect 21189 16745 21223 16779
rect 21373 16745 21407 16779
rect 24409 16745 24443 16779
rect 27445 16745 27479 16779
rect 28089 16745 28123 16779
rect 17785 16677 17819 16711
rect 20821 16677 20855 16711
rect 25789 16677 25823 16711
rect 31217 16677 31251 16711
rect 33885 16677 33919 16711
rect 1869 16609 1903 16643
rect 13553 16609 13587 16643
rect 14473 16609 14507 16643
rect 15209 16609 15243 16643
rect 16405 16609 16439 16643
rect 17233 16609 17267 16643
rect 17693 16609 17727 16643
rect 19901 16609 19935 16643
rect 20361 16609 20395 16643
rect 22201 16609 22235 16643
rect 24501 16609 24535 16643
rect 26433 16609 26467 16643
rect 41705 16609 41739 16643
rect 42165 16609 42199 16643
rect 1409 16541 1443 16575
rect 13277 16541 13311 16575
rect 14289 16541 14323 16575
rect 15117 16541 15151 16575
rect 16129 16541 16163 16575
rect 16865 16541 16899 16575
rect 17969 16541 18003 16575
rect 19257 16541 19291 16575
rect 19441 16541 19475 16575
rect 19993 16541 20027 16575
rect 20177 16541 20211 16575
rect 22017 16541 22051 16575
rect 24685 16541 24719 16575
rect 25421 16541 25455 16575
rect 25605 16541 25639 16575
rect 25789 16541 25823 16575
rect 26617 16541 26651 16575
rect 28181 16541 28215 16575
rect 30849 16541 30883 16575
rect 30941 16541 30975 16575
rect 31033 16541 31067 16575
rect 32500 16541 32534 16575
rect 32597 16541 32631 16575
rect 32872 16541 32906 16575
rect 32965 16541 32999 16575
rect 33609 16541 33643 16575
rect 34989 16541 35023 16575
rect 35173 16541 35207 16575
rect 37657 16541 37691 16575
rect 1593 16473 1627 16507
rect 17049 16473 17083 16507
rect 19349 16473 19383 16507
rect 21833 16473 21867 16507
rect 24409 16473 24443 16507
rect 26801 16473 26835 16507
rect 27353 16473 27387 16507
rect 32689 16473 32723 16507
rect 41981 16473 42015 16507
rect 14105 16405 14139 16439
rect 15485 16405 15519 16439
rect 15945 16405 15979 16439
rect 21189 16405 21223 16439
rect 24869 16405 24903 16439
rect 32321 16405 32355 16439
rect 34069 16405 34103 16439
rect 35081 16405 35115 16439
rect 37473 16405 37507 16439
rect 2145 16201 2179 16235
rect 18061 16201 18095 16235
rect 20729 16201 20763 16235
rect 41429 16201 41463 16235
rect 14749 16133 14783 16167
rect 22262 16133 22296 16167
rect 31033 16133 31067 16167
rect 32229 16133 32263 16167
rect 14979 16099 15013 16133
rect 1409 16065 1443 16099
rect 2237 16065 2271 16099
rect 12817 16065 12851 16099
rect 13001 16065 13035 16099
rect 15761 16065 15795 16099
rect 17969 16065 18003 16099
rect 18245 16065 18279 16099
rect 19605 16065 19639 16099
rect 22017 16065 22051 16099
rect 24317 16065 24351 16099
rect 24593 16065 24627 16099
rect 24777 16065 24811 16099
rect 25237 16065 25271 16099
rect 26249 16065 26283 16099
rect 26433 16065 26467 16099
rect 26985 16065 27019 16099
rect 27241 16065 27275 16099
rect 29101 16065 29135 16099
rect 30665 16065 30699 16099
rect 31125 16065 31159 16099
rect 32597 16065 32631 16099
rect 33425 16065 33459 16099
rect 34437 16065 34471 16099
rect 35449 16065 35483 16099
rect 37289 16065 37323 16099
rect 40877 16065 40911 16099
rect 41337 16065 41371 16099
rect 13461 15997 13495 16031
rect 13737 15997 13771 16031
rect 18429 15997 18463 16031
rect 19349 15997 19383 16031
rect 25329 15997 25363 16031
rect 26341 15997 26375 16031
rect 28825 15997 28859 16031
rect 29009 15997 29043 16031
rect 30849 15997 30883 16031
rect 32689 15997 32723 16031
rect 33333 15997 33367 16031
rect 33793 15997 33827 16031
rect 34345 15997 34379 16031
rect 35357 15997 35391 16031
rect 37473 15997 37507 16031
rect 38945 15997 38979 16031
rect 23397 15929 23431 15963
rect 28365 15929 28399 15963
rect 13001 15861 13035 15895
rect 14933 15861 14967 15895
rect 15117 15861 15151 15895
rect 15669 15861 15703 15895
rect 24455 15861 24489 15895
rect 24685 15861 24719 15895
rect 25237 15861 25271 15895
rect 25605 15861 25639 15895
rect 28917 15861 28951 15895
rect 32321 15861 32355 15895
rect 34713 15861 34747 15895
rect 35817 15861 35851 15895
rect 40233 15861 40267 15895
rect 40785 15861 40819 15895
rect 11529 15657 11563 15691
rect 13553 15657 13587 15691
rect 18153 15657 18187 15691
rect 21649 15657 21683 15691
rect 28825 15657 28859 15691
rect 33701 15657 33735 15691
rect 37289 15657 37323 15691
rect 34989 15589 35023 15623
rect 12909 15521 12943 15555
rect 15392 15521 15426 15555
rect 15485 15521 15519 15555
rect 16129 15521 16163 15555
rect 24961 15521 24995 15555
rect 29561 15521 29595 15555
rect 34713 15521 34747 15555
rect 35633 15521 35667 15555
rect 40325 15521 40359 15555
rect 40509 15521 40543 15555
rect 42165 15521 42199 15555
rect 1777 15453 1811 15487
rect 13369 15453 13403 15487
rect 13553 15453 13587 15487
rect 14105 15453 14139 15487
rect 14381 15453 14415 15487
rect 14473 15453 14507 15487
rect 15209 15453 15243 15487
rect 15301 15453 15335 15487
rect 16221 15453 16255 15487
rect 16405 15453 16439 15487
rect 17417 15453 17451 15487
rect 17601 15453 17635 15487
rect 18061 15453 18095 15487
rect 18337 15453 18371 15487
rect 20821 15453 20855 15487
rect 21373 15453 21407 15487
rect 21833 15453 21867 15487
rect 25053 15453 25087 15487
rect 27445 15453 27479 15487
rect 27712 15453 27746 15487
rect 29817 15453 29851 15487
rect 33241 15453 33275 15487
rect 33333 15453 33367 15487
rect 33517 15453 33551 15487
rect 35909 15453 35943 15487
rect 37197 15453 37231 15487
rect 12664 15385 12698 15419
rect 14289 15385 14323 15419
rect 19625 15385 19659 15419
rect 19809 15385 19843 15419
rect 20637 15385 20671 15419
rect 21465 15385 21499 15419
rect 14657 15317 14691 15351
rect 15669 15317 15703 15351
rect 17509 15317 17543 15351
rect 18521 15317 18555 15351
rect 25421 15317 25455 15351
rect 30941 15317 30975 15351
rect 35173 15317 35207 15351
rect 13185 15113 13219 15147
rect 18061 15113 18095 15147
rect 24987 15113 25021 15147
rect 14749 15045 14783 15079
rect 15945 15045 15979 15079
rect 16926 15045 16960 15079
rect 22753 15045 22787 15079
rect 23673 15045 23707 15079
rect 24777 15045 24811 15079
rect 30941 15045 30975 15079
rect 1777 14977 1811 15011
rect 13461 14977 13495 15011
rect 13550 14983 13584 15017
rect 13645 14977 13679 15011
rect 13829 14977 13863 15011
rect 14381 14977 14415 15011
rect 14841 14977 14875 15011
rect 15301 14977 15335 15011
rect 15485 14977 15519 15011
rect 15577 14977 15611 15011
rect 15669 14977 15703 15011
rect 18797 14977 18831 15011
rect 19993 14977 20027 15011
rect 20729 14977 20763 15011
rect 20913 14977 20947 15011
rect 30113 14977 30147 15011
rect 30297 14977 30331 15011
rect 30757 14977 30791 15011
rect 35357 14977 35391 15011
rect 35541 14977 35575 15011
rect 1961 14909 1995 14943
rect 2789 14909 2823 14943
rect 14565 14909 14599 14943
rect 16681 14909 16715 14943
rect 19717 14909 19751 14943
rect 20637 14909 20671 14943
rect 22385 14909 22419 14943
rect 41337 14909 41371 14943
rect 41705 14909 41739 14943
rect 41889 14909 41923 14943
rect 19073 14841 19107 14875
rect 19257 14841 19291 14875
rect 20177 14841 20211 14875
rect 22937 14841 22971 14875
rect 19809 14773 19843 14807
rect 21097 14773 21131 14807
rect 22753 14773 22787 14807
rect 23581 14773 23615 14807
rect 24961 14773 24995 14807
rect 25145 14773 25179 14807
rect 30205 14773 30239 14807
rect 31125 14773 31159 14807
rect 35725 14773 35759 14807
rect 2237 14569 2271 14603
rect 13369 14569 13403 14603
rect 19625 14569 19659 14603
rect 20729 14569 20763 14603
rect 21741 14569 21775 14603
rect 24869 14569 24903 14603
rect 35541 14569 35575 14603
rect 35817 14569 35851 14603
rect 41429 14569 41463 14603
rect 41981 14569 42015 14603
rect 23581 14501 23615 14535
rect 15485 14433 15519 14467
rect 15761 14433 15795 14467
rect 15853 14433 15887 14467
rect 17601 14433 17635 14467
rect 17877 14433 17911 14467
rect 19257 14433 19291 14467
rect 20361 14433 20395 14467
rect 2329 14365 2363 14399
rect 12357 14365 12391 14399
rect 13277 14365 13311 14399
rect 13461 14365 13495 14399
rect 14657 14365 14691 14399
rect 14749 14365 14783 14399
rect 14841 14365 14875 14399
rect 15025 14365 15059 14399
rect 15669 14365 15703 14399
rect 15945 14365 15979 14399
rect 19441 14365 19475 14399
rect 20269 14365 20303 14399
rect 20545 14365 20579 14399
rect 21373 14365 21407 14399
rect 23397 14365 23431 14399
rect 26249 14365 26283 14399
rect 26709 14365 26743 14399
rect 26976 14365 27010 14399
rect 29561 14365 29595 14399
rect 29828 14365 29862 14399
rect 32045 14365 32079 14399
rect 33609 14365 33643 14399
rect 33793 14365 33827 14399
rect 34897 14365 34931 14399
rect 35725 14365 35759 14399
rect 36093 14365 36127 14399
rect 36553 14365 36587 14399
rect 36737 14365 36771 14399
rect 41337 14365 41371 14399
rect 21741 14297 21775 14331
rect 26004 14297 26038 14331
rect 33057 14297 33091 14331
rect 35081 14297 35115 14331
rect 12173 14229 12207 14263
rect 14381 14229 14415 14263
rect 21925 14229 21959 14263
rect 28089 14229 28123 14263
rect 30941 14229 30975 14263
rect 33701 14229 33735 14263
rect 34713 14229 34747 14263
rect 36645 14229 36679 14263
rect 15485 14025 15519 14059
rect 16681 14025 16715 14059
rect 19901 14025 19935 14059
rect 24593 14025 24627 14059
rect 26157 14025 26191 14059
rect 32229 14025 32263 14059
rect 33333 14025 33367 14059
rect 14372 13957 14406 13991
rect 16833 13957 16867 13991
rect 17049 13957 17083 13991
rect 21925 13957 21959 13991
rect 22109 13957 22143 13991
rect 22814 13957 22848 13991
rect 27721 13957 27755 13991
rect 31585 13957 31619 13991
rect 34713 13957 34747 13991
rect 11805 13889 11839 13923
rect 14105 13889 14139 13923
rect 18061 13889 18095 13923
rect 19809 13889 19843 13923
rect 19993 13889 20027 13923
rect 20453 13889 20487 13923
rect 22569 13889 22603 13923
rect 24777 13889 24811 13923
rect 25237 13889 25271 13923
rect 25421 13889 25455 13923
rect 26341 13889 26375 13923
rect 30113 13889 30147 13923
rect 30297 13889 30331 13923
rect 31125 13889 31159 13923
rect 32137 13889 32171 13923
rect 32321 13889 32355 13923
rect 33241 13889 33275 13923
rect 34529 13889 34563 13923
rect 34621 13889 34655 13923
rect 34831 13889 34865 13923
rect 35633 13889 35667 13923
rect 1961 13821 1995 13855
rect 2145 13821 2179 13855
rect 2881 13821 2915 13855
rect 11989 13821 12023 13855
rect 13645 13821 13679 13855
rect 18245 13821 18279 13855
rect 20729 13821 20763 13855
rect 31217 13821 31251 13855
rect 33425 13821 33459 13855
rect 34989 13821 35023 13855
rect 35909 13821 35943 13855
rect 20637 13753 20671 13787
rect 23949 13753 23983 13787
rect 27537 13753 27571 13787
rect 16865 13685 16899 13719
rect 17877 13685 17911 13719
rect 20545 13685 20579 13719
rect 25329 13685 25363 13719
rect 30113 13685 30147 13719
rect 30941 13685 30975 13719
rect 32873 13685 32907 13719
rect 34345 13685 34379 13719
rect 41797 13685 41831 13719
rect 2053 13481 2087 13515
rect 2789 13481 2823 13515
rect 12081 13481 12115 13515
rect 21557 13481 21591 13515
rect 21925 13481 21959 13515
rect 24869 13481 24903 13515
rect 25421 13481 25455 13515
rect 28181 13481 28215 13515
rect 28365 13481 28399 13515
rect 34713 13481 34747 13515
rect 36829 13481 36863 13515
rect 17693 13413 17727 13447
rect 17601 13345 17635 13379
rect 20269 13345 20303 13379
rect 22477 13345 22511 13379
rect 25789 13345 25823 13379
rect 29929 13345 29963 13379
rect 32045 13345 32079 13379
rect 33425 13345 33459 13379
rect 33517 13345 33551 13379
rect 35449 13345 35483 13379
rect 41337 13345 41371 13379
rect 42165 13345 42199 13379
rect 2881 13277 2915 13311
rect 12173 13277 12207 13311
rect 12817 13277 12851 13311
rect 16129 13277 16163 13311
rect 16405 13277 16439 13311
rect 16589 13277 16623 13311
rect 17877 13277 17911 13311
rect 20545 13277 20579 13311
rect 21557 13277 21591 13311
rect 21649 13277 21683 13311
rect 22733 13277 22767 13311
rect 24685 13277 24719 13311
rect 24869 13277 24903 13311
rect 25329 13277 25363 13311
rect 26341 13277 26375 13311
rect 28733 13277 28767 13311
rect 30113 13277 30147 13311
rect 31033 13277 31067 13311
rect 31401 13277 31435 13311
rect 33333 13277 33367 13311
rect 34713 13277 34747 13311
rect 34989 13277 35023 13311
rect 35725 13277 35759 13311
rect 36737 13277 36771 13311
rect 36921 13277 36955 13311
rect 37381 13277 37415 13311
rect 16221 13209 16255 13243
rect 30297 13209 30331 13243
rect 41981 13209 42015 13243
rect 12725 13141 12759 13175
rect 18061 13141 18095 13175
rect 23857 13141 23891 13175
rect 26525 13141 26559 13175
rect 28365 13141 28399 13175
rect 32965 13141 32999 13175
rect 34897 13141 34931 13175
rect 37473 13141 37507 13175
rect 19717 12937 19751 12971
rect 21189 12937 21223 12971
rect 29285 12937 29319 12971
rect 32229 12937 32263 12971
rect 33609 12937 33643 12971
rect 34069 12937 34103 12971
rect 34897 12937 34931 12971
rect 35541 12937 35575 12971
rect 36001 12937 36035 12971
rect 41521 12937 41555 12971
rect 12357 12869 12391 12903
rect 15025 12869 15059 12903
rect 18582 12869 18616 12903
rect 22017 12869 22051 12903
rect 26341 12869 26375 12903
rect 31309 12869 31343 12903
rect 15209 12801 15243 12835
rect 15853 12801 15887 12835
rect 16129 12801 16163 12835
rect 16681 12801 16715 12835
rect 18337 12801 18371 12835
rect 20913 12801 20947 12835
rect 21005 12801 21039 12835
rect 21833 12801 21867 12835
rect 23949 12801 23983 12835
rect 24225 12801 24259 12835
rect 25053 12801 25087 12835
rect 27252 12801 27286 12835
rect 28825 12801 28859 12835
rect 29101 12801 29135 12835
rect 30297 12801 30331 12835
rect 30573 12801 30607 12835
rect 30757 12801 30791 12835
rect 32137 12801 32171 12835
rect 32321 12801 32355 12835
rect 33977 12801 34011 12835
rect 35357 12801 35391 12835
rect 36139 12801 36173 12835
rect 36277 12801 36311 12835
rect 36369 12801 36403 12835
rect 36497 12801 36531 12835
rect 36645 12801 36679 12835
rect 37841 12801 37875 12835
rect 41429 12801 41463 12835
rect 12173 12733 12207 12767
rect 13737 12733 13771 12767
rect 15945 12733 15979 12767
rect 16957 12733 16991 12767
rect 24133 12733 24167 12767
rect 25145 12733 25179 12767
rect 26985 12733 27019 12767
rect 29009 12733 29043 12767
rect 34253 12733 34287 12767
rect 35265 12733 35299 12767
rect 15669 12665 15703 12699
rect 26157 12665 26191 12699
rect 31493 12665 31527 12699
rect 37657 12665 37691 12699
rect 1685 12597 1719 12631
rect 16129 12597 16163 12631
rect 22201 12597 22235 12631
rect 24225 12597 24259 12631
rect 24409 12597 24443 12631
rect 25421 12597 25455 12631
rect 28365 12597 28399 12631
rect 28825 12597 28859 12631
rect 30573 12597 30607 12631
rect 40785 12597 40819 12631
rect 12725 12393 12759 12427
rect 15669 12393 15703 12427
rect 16221 12393 16255 12427
rect 17233 12393 17267 12427
rect 20177 12393 20211 12427
rect 20361 12393 20395 12427
rect 24409 12393 24443 12427
rect 24777 12393 24811 12427
rect 27445 12393 27479 12427
rect 34897 12393 34931 12427
rect 17601 12325 17635 12359
rect 19349 12325 19383 12359
rect 1409 12257 1443 12291
rect 2789 12257 2823 12291
rect 14289 12257 14323 12291
rect 21005 12257 21039 12291
rect 28549 12257 28583 12291
rect 29009 12257 29043 12291
rect 30205 12257 30239 12291
rect 31125 12257 31159 12291
rect 32505 12257 32539 12291
rect 33885 12257 33919 12291
rect 34161 12257 34195 12291
rect 36921 12257 36955 12291
rect 40325 12257 40359 12291
rect 42165 12257 42199 12291
rect 12909 12189 12943 12223
rect 16405 12189 16439 12223
rect 18245 12189 18279 12223
rect 18521 12189 18555 12223
rect 19257 12189 19291 12223
rect 19441 12189 19475 12223
rect 21189 12189 21223 12223
rect 24409 12189 24443 12223
rect 24593 12189 24627 12223
rect 26065 12189 26099 12223
rect 26332 12189 26366 12223
rect 28641 12189 28675 12223
rect 30481 12189 30515 12223
rect 32321 12189 32355 12223
rect 32413 12189 32447 12223
rect 36001 12189 36035 12223
rect 36829 12189 36863 12223
rect 37013 12189 37047 12223
rect 1593 12121 1627 12155
rect 14556 12121 14590 12155
rect 16589 12121 16623 12155
rect 18429 12121 18463 12155
rect 20545 12121 20579 12155
rect 34881 12121 34915 12155
rect 35081 12121 35115 12155
rect 36185 12121 36219 12155
rect 40509 12121 40543 12155
rect 17049 12053 17083 12087
rect 17233 12053 17267 12087
rect 18061 12053 18095 12087
rect 20345 12053 20379 12087
rect 31953 12053 31987 12087
rect 34713 12053 34747 12087
rect 36369 12053 36403 12087
rect 2145 11849 2179 11883
rect 14749 11849 14783 11883
rect 16773 11849 16807 11883
rect 19901 11849 19935 11883
rect 23857 11849 23891 11883
rect 24317 11849 24351 11883
rect 28365 11849 28399 11883
rect 41521 11849 41555 11883
rect 19073 11781 19107 11815
rect 19289 11781 19323 11815
rect 27230 11781 27264 11815
rect 34437 11781 34471 11815
rect 2237 11713 2271 11747
rect 9413 11713 9447 11747
rect 14933 11713 14967 11747
rect 16957 11713 16991 11747
rect 17693 11713 17727 11747
rect 21025 11713 21059 11747
rect 21281 11713 21315 11747
rect 22477 11713 22511 11747
rect 22733 11713 22767 11747
rect 25430 11713 25464 11747
rect 26985 11713 27019 11747
rect 30665 11713 30699 11747
rect 33425 11713 33459 11747
rect 33701 11713 33735 11747
rect 33885 11713 33919 11747
rect 34345 11713 34379 11747
rect 34621 11713 34655 11747
rect 35082 11735 35116 11769
rect 35817 11713 35851 11747
rect 41613 11713 41647 11747
rect 17141 11645 17175 11679
rect 17969 11645 18003 11679
rect 25697 11645 25731 11679
rect 35357 11645 35391 11679
rect 36093 11645 36127 11679
rect 35173 11577 35207 11611
rect 9321 11509 9355 11543
rect 19257 11509 19291 11543
rect 19441 11509 19475 11543
rect 30481 11509 30515 11543
rect 33241 11509 33275 11543
rect 34345 11509 34379 11543
rect 35265 11509 35299 11543
rect 40785 11509 40819 11543
rect 19533 11305 19567 11339
rect 21005 11305 21039 11339
rect 21649 11305 21683 11339
rect 22845 11305 22879 11339
rect 36829 11305 36863 11339
rect 33885 11237 33919 11271
rect 33977 11169 34011 11203
rect 34713 11169 34747 11203
rect 36093 11169 36127 11203
rect 36185 11169 36219 11203
rect 40325 11169 40359 11203
rect 1685 11101 1719 11135
rect 17233 11101 17267 11135
rect 17785 11101 17819 11135
rect 18061 11101 18095 11135
rect 19717 11101 19751 11135
rect 19993 11101 20027 11135
rect 21097 11101 21131 11135
rect 21833 11101 21867 11135
rect 22661 11101 22695 11135
rect 26341 11101 26375 11135
rect 33514 11101 33548 11135
rect 34897 11101 34931 11135
rect 35081 11101 35115 11135
rect 36001 11101 36035 11135
rect 36829 11101 36863 11135
rect 37013 11101 37047 11135
rect 37473 11101 37507 11135
rect 37657 11101 37691 11135
rect 40509 11033 40543 11067
rect 42165 11033 42199 11067
rect 17141 10965 17175 10999
rect 19901 10965 19935 10999
rect 25697 10965 25731 10999
rect 33333 10965 33367 10999
rect 33517 10965 33551 10999
rect 35633 10965 35667 10999
rect 37565 10965 37599 10999
rect 21281 10761 21315 10795
rect 23857 10761 23891 10795
rect 25697 10761 25731 10795
rect 28365 10761 28399 10795
rect 32873 10761 32907 10795
rect 34989 10761 35023 10795
rect 41429 10761 41463 10795
rect 18153 10693 18187 10727
rect 24562 10693 24596 10727
rect 28825 10693 28859 10727
rect 30674 10693 30708 10727
rect 1685 10625 1719 10659
rect 14749 10625 14783 10659
rect 15005 10625 15039 10659
rect 18521 10625 18555 10659
rect 19349 10625 19383 10659
rect 19441 10625 19475 10659
rect 19901 10625 19935 10659
rect 20157 10625 20191 10659
rect 23029 10625 23063 10659
rect 23213 10625 23247 10659
rect 23673 10625 23707 10659
rect 28733 10625 28767 10659
rect 30941 10625 30975 10659
rect 31585 10625 31619 10659
rect 32965 10625 32999 10659
rect 34897 10625 34931 10659
rect 36001 10625 36035 10659
rect 36093 10625 36127 10659
rect 36185 10625 36219 10659
rect 36369 10625 36403 10659
rect 41521 10625 41555 10659
rect 1869 10557 1903 10591
rect 2789 10557 2823 10591
rect 16681 10557 16715 10591
rect 16957 10557 16991 10591
rect 19165 10557 19199 10591
rect 22845 10557 22879 10591
rect 24317 10557 24351 10591
rect 28917 10557 28951 10591
rect 33057 10557 33091 10591
rect 35081 10557 35115 10591
rect 16129 10489 16163 10523
rect 17969 10421 18003 10455
rect 18153 10421 18187 10455
rect 19257 10421 19291 10455
rect 29561 10421 29595 10455
rect 31401 10421 31435 10455
rect 32505 10421 32539 10455
rect 34529 10421 34563 10455
rect 35725 10421 35759 10455
rect 40693 10421 40727 10455
rect 2053 10217 2087 10251
rect 14841 10217 14875 10251
rect 15853 10217 15887 10251
rect 16497 10217 16531 10251
rect 16681 10217 16715 10251
rect 18705 10217 18739 10251
rect 19625 10217 19659 10251
rect 22569 10217 22603 10251
rect 23213 10217 23247 10251
rect 32597 10217 32631 10251
rect 35173 10217 35207 10251
rect 35725 10217 35759 10251
rect 17325 10081 17359 10115
rect 33057 10081 33091 10115
rect 33149 10081 33183 10115
rect 34989 10081 35023 10115
rect 40325 10081 40359 10115
rect 42165 10081 42199 10115
rect 2145 10013 2179 10047
rect 2789 10013 2823 10047
rect 15117 10013 15151 10047
rect 15577 10013 15611 10047
rect 15853 10013 15887 10047
rect 19625 10013 19659 10047
rect 19901 10013 19935 10047
rect 21925 10013 21959 10047
rect 22385 10013 22419 10047
rect 23029 10013 23063 10047
rect 25421 10013 25455 10047
rect 27353 10013 27387 10047
rect 31401 10013 31435 10047
rect 32965 10013 32999 10047
rect 35265 10013 35299 10047
rect 35725 10013 35759 10047
rect 35909 10013 35943 10047
rect 36001 10013 36035 10047
rect 14841 9945 14875 9979
rect 16313 9945 16347 9979
rect 17592 9945 17626 9979
rect 19809 9945 19843 9979
rect 25688 9945 25722 9979
rect 27620 9945 27654 9979
rect 31134 9945 31168 9979
rect 40509 9945 40543 9979
rect 15025 9877 15059 9911
rect 15669 9877 15703 9911
rect 16513 9877 16547 9911
rect 21741 9877 21775 9911
rect 28733 9877 28767 9911
rect 30021 9877 30055 9911
rect 34713 9877 34747 9911
rect 18613 9673 18647 9707
rect 27905 9673 27939 9707
rect 30021 9673 30055 9707
rect 30481 9673 30515 9707
rect 15577 9605 15611 9639
rect 26249 9605 26283 9639
rect 33333 9605 33367 9639
rect 33977 9605 34011 9639
rect 41429 9605 41463 9639
rect 2329 9537 2363 9571
rect 2973 9537 3007 9571
rect 15761 9537 15795 9571
rect 15853 9537 15887 9571
rect 18429 9537 18463 9571
rect 21833 9537 21867 9571
rect 22017 9537 22051 9571
rect 22661 9537 22695 9571
rect 23572 9537 23606 9571
rect 25329 9537 25363 9571
rect 25421 9537 25455 9571
rect 25605 9537 25639 9571
rect 26065 9537 26099 9571
rect 26433 9537 26467 9571
rect 26985 9537 27019 9571
rect 29029 9537 29063 9571
rect 29285 9537 29319 9571
rect 30389 9537 30423 9571
rect 32321 9537 32355 9571
rect 33517 9537 33551 9571
rect 41337 9537 41371 9571
rect 15577 9469 15611 9503
rect 18153 9469 18187 9503
rect 18245 9469 18279 9503
rect 18337 9469 18371 9503
rect 23305 9469 23339 9503
rect 30573 9469 30607 9503
rect 33609 9469 33643 9503
rect 22201 9401 22235 9435
rect 24685 9401 24719 9435
rect 25145 9401 25179 9435
rect 27169 9401 27203 9435
rect 1685 9333 1719 9367
rect 2237 9333 2271 9367
rect 2881 9333 2915 9367
rect 22845 9333 22879 9367
rect 25329 9333 25363 9367
rect 32137 9333 32171 9367
rect 17969 9129 18003 9163
rect 19901 9129 19935 9163
rect 21649 9129 21683 9163
rect 22477 9129 22511 9163
rect 30205 9129 30239 9163
rect 3065 8993 3099 9027
rect 3249 8993 3283 9027
rect 16497 8993 16531 9027
rect 21281 8993 21315 9027
rect 22109 8993 22143 9027
rect 22937 8993 22971 9027
rect 31493 8993 31527 9027
rect 1409 8925 1443 8959
rect 15485 8925 15519 8959
rect 15669 8925 15703 8959
rect 16129 8925 16163 8959
rect 16313 8925 16347 8959
rect 18153 8925 18187 8959
rect 21465 8925 21499 8959
rect 22293 8925 22327 8959
rect 23121 8925 23155 8959
rect 26341 8925 26375 8959
rect 26525 8925 26559 8959
rect 26985 8925 27019 8959
rect 28365 8925 28399 8959
rect 29561 8925 29595 8959
rect 31760 8925 31794 8959
rect 20085 8857 20119 8891
rect 26157 8857 26191 8891
rect 15577 8789 15611 8823
rect 19717 8789 19751 8823
rect 19885 8789 19919 8823
rect 23305 8789 23339 8823
rect 27169 8789 27203 8823
rect 29009 8789 29043 8823
rect 32873 8789 32907 8823
rect 16129 8585 16163 8619
rect 20913 8585 20947 8619
rect 22201 8585 22235 8619
rect 24409 8585 24443 8619
rect 28641 8585 28675 8619
rect 30481 8585 30515 8619
rect 1961 8517 1995 8551
rect 15016 8517 15050 8551
rect 19901 8517 19935 8551
rect 20545 8517 20579 8551
rect 23274 8517 23308 8551
rect 27506 8517 27540 8551
rect 30941 8517 30975 8551
rect 1777 8449 1811 8483
rect 14749 8449 14783 8483
rect 17509 8449 17543 8483
rect 19533 8449 19567 8483
rect 20729 8449 20763 8483
rect 21005 8449 21039 8483
rect 21833 8449 21867 8483
rect 22017 8449 22051 8483
rect 23029 8449 23063 8483
rect 27261 8449 27295 8483
rect 29101 8449 29135 8483
rect 29357 8449 29391 8483
rect 2789 8381 2823 8415
rect 17233 8381 17267 8415
rect 17417 8381 17451 8415
rect 18245 8381 18279 8415
rect 31401 8381 31435 8415
rect 18521 8313 18555 8347
rect 20085 8313 20119 8347
rect 31309 8313 31343 8347
rect 17325 8245 17359 8279
rect 18705 8245 18739 8279
rect 19901 8245 19935 8279
rect 16037 8041 16071 8075
rect 16129 8041 16163 8075
rect 18245 8041 18279 8075
rect 20637 8041 20671 8075
rect 22477 8041 22511 8075
rect 23121 8041 23155 8075
rect 15945 7905 15979 7939
rect 16865 7905 16899 7939
rect 25329 7905 25363 7939
rect 16221 7837 16255 7871
rect 19257 7837 19291 7871
rect 21097 7837 21131 7871
rect 22937 7837 22971 7871
rect 23765 7837 23799 7871
rect 41705 7837 41739 7871
rect 17132 7769 17166 7803
rect 19502 7769 19536 7803
rect 21342 7769 21376 7803
rect 25596 7769 25630 7803
rect 23581 7701 23615 7735
rect 41613 7701 41647 7735
rect 17325 7497 17359 7531
rect 18797 7497 18831 7531
rect 24409 7497 24443 7531
rect 25513 7497 25547 7531
rect 17141 7429 17175 7463
rect 23296 7429 23330 7463
rect 17417 7361 17451 7395
rect 18613 7361 18647 7395
rect 19993 7361 20027 7395
rect 23029 7361 23063 7395
rect 24869 7361 24903 7395
rect 41889 7361 41923 7395
rect 20269 7293 20303 7327
rect 17141 7225 17175 7259
rect 41705 7225 41739 7259
rect 40969 7157 41003 7191
rect 40325 6817 40359 6851
rect 4261 6749 4295 6783
rect 20269 6749 20303 6783
rect 40509 6681 40543 6715
rect 42165 6681 42199 6715
rect 4169 6613 4203 6647
rect 20453 6613 20487 6647
rect 4169 6341 4203 6375
rect 2881 6273 2915 6307
rect 3985 6205 4019 6239
rect 5089 6205 5123 6239
rect 1409 6069 1443 6103
rect 2053 6069 2087 6103
rect 2789 6069 2823 6103
rect 40969 6069 41003 6103
rect 41797 6069 41831 6103
rect 4445 5865 4479 5899
rect 1409 5729 1443 5763
rect 1869 5729 1903 5763
rect 40877 5729 40911 5763
rect 3985 5661 4019 5695
rect 37841 5661 37875 5695
rect 38577 5661 38611 5695
rect 39865 5661 39899 5695
rect 41337 5661 41371 5695
rect 41981 5661 42015 5695
rect 1593 5593 1627 5627
rect 37933 5525 37967 5559
rect 41429 5525 41463 5559
rect 42073 5525 42107 5559
rect 2145 5253 2179 5287
rect 38669 5253 38703 5287
rect 1961 5185 1995 5219
rect 38485 5185 38519 5219
rect 40969 5185 41003 5219
rect 41429 5185 41463 5219
rect 2789 5117 2823 5151
rect 40325 5117 40359 5151
rect 4261 4981 4295 5015
rect 40877 4981 40911 5015
rect 41521 4981 41555 5015
rect 2145 4777 2179 4811
rect 4629 4641 4663 4675
rect 40325 4641 40359 4675
rect 40509 4641 40543 4675
rect 41889 4641 41923 4675
rect 1409 4573 1443 4607
rect 2237 4573 2271 4607
rect 2881 4573 2915 4607
rect 3985 4573 4019 4607
rect 5089 4573 5123 4607
rect 36737 4573 36771 4607
rect 37841 4573 37875 4607
rect 38669 4573 38703 4607
rect 39129 4573 39163 4607
rect 3893 4437 3927 4471
rect 39221 4437 39255 4471
rect 39773 4165 39807 4199
rect 2145 4097 2179 4131
rect 3157 4097 3191 4131
rect 4997 4097 5031 4131
rect 5641 4097 5675 4131
rect 37841 4097 37875 4131
rect 38761 4097 38795 4131
rect 39589 4097 39623 4131
rect 4813 4029 4847 4063
rect 22661 4029 22695 4063
rect 22845 4029 22879 4063
rect 23213 4029 23247 4063
rect 41337 4029 41371 4063
rect 9413 3961 9447 3995
rect 2053 3893 2087 3927
rect 5549 3893 5583 3927
rect 6377 3893 6411 3927
rect 9873 3893 9907 3927
rect 10977 3893 11011 3927
rect 11529 3893 11563 3927
rect 18153 3893 18187 3927
rect 19625 3893 19659 3927
rect 21925 3893 21959 3927
rect 34713 3893 34747 3927
rect 35633 3893 35667 3927
rect 36737 3893 36771 3927
rect 37933 3893 37967 3927
rect 38669 3893 38703 3927
rect 22477 3689 22511 3723
rect 3065 3553 3099 3587
rect 3249 3553 3283 3587
rect 4721 3553 4755 3587
rect 4905 3553 4939 3587
rect 5181 3553 5215 3587
rect 9045 3553 9079 3587
rect 9229 3553 9263 3587
rect 9689 3553 9723 3587
rect 11345 3553 11379 3587
rect 11805 3553 11839 3587
rect 16865 3553 16899 3587
rect 19533 3553 19567 3587
rect 19993 3553 20027 3587
rect 34713 3553 34747 3587
rect 35173 3553 35207 3587
rect 37013 3553 37047 3587
rect 37473 3553 37507 3587
rect 42165 3553 42199 3587
rect 1409 3485 1443 3519
rect 4261 3485 4295 3519
rect 7297 3485 7331 3519
rect 8217 3485 8251 3519
rect 14841 3485 14875 3519
rect 15669 3485 15703 3519
rect 16129 3485 16163 3519
rect 18613 3485 18647 3519
rect 23121 3485 23155 3519
rect 23581 3485 23615 3519
rect 27813 3485 27847 3519
rect 11529 3417 11563 3451
rect 16313 3417 16347 3451
rect 19717 3417 19751 3451
rect 34897 3417 34931 3451
rect 37197 3417 37231 3451
rect 40325 3417 40359 3451
rect 41981 3417 42015 3451
rect 4169 3349 4203 3383
rect 8125 3349 8159 3383
rect 18521 3349 18555 3383
rect 23673 3349 23707 3383
rect 16773 3145 16807 3179
rect 20545 3145 20579 3179
rect 22753 3145 22787 3179
rect 3709 3077 3743 3111
rect 5365 3077 5399 3111
rect 7389 3077 7423 3111
rect 18337 3077 18371 3111
rect 23673 3077 23707 3111
rect 37749 3077 37783 3111
rect 40049 3077 40083 3111
rect 1409 3009 1443 3043
rect 5549 3009 5583 3043
rect 6377 3009 6411 3043
rect 7205 3009 7239 3043
rect 10241 3009 10275 3043
rect 10977 3009 11011 3043
rect 11529 3009 11563 3043
rect 14289 3009 14323 3043
rect 16865 3009 16899 3043
rect 18153 3009 18187 3043
rect 20637 3009 20671 3043
rect 21925 3009 21959 3043
rect 22661 3009 22695 3043
rect 23489 3009 23523 3043
rect 27813 3009 27847 3043
rect 34897 3009 34931 3043
rect 37565 3009 37599 3043
rect 39865 3009 39899 3043
rect 1593 2941 1627 2975
rect 2789 2941 2823 2975
rect 7665 2941 7699 2975
rect 10885 2941 10919 2975
rect 11713 2941 11747 2975
rect 11989 2941 12023 2975
rect 14473 2941 14507 2975
rect 15485 2941 15519 2975
rect 18705 2941 18739 2975
rect 23949 2941 23983 2975
rect 27997 2941 28031 2975
rect 28365 2941 28399 2975
rect 35081 2941 35115 2975
rect 36093 2941 36127 2975
rect 39313 2941 39347 2975
rect 40601 2941 40635 2975
rect 6469 2805 6503 2839
rect 10149 2805 10183 2839
rect 22017 2805 22051 2839
rect 2053 2601 2087 2635
rect 11621 2601 11655 2635
rect 15209 2601 15243 2635
rect 27905 2601 27939 2635
rect 35817 2601 35851 2635
rect 36461 2601 36495 2635
rect 3801 2465 3835 2499
rect 4261 2465 4295 2499
rect 6377 2465 6411 2499
rect 6561 2465 6595 2499
rect 6929 2465 6963 2499
rect 9137 2465 9171 2499
rect 10793 2465 10827 2499
rect 21833 2465 21867 2499
rect 22017 2465 22051 2499
rect 22569 2465 22603 2499
rect 37473 2465 37507 2499
rect 37657 2465 37691 2499
rect 41337 2465 41371 2499
rect 41705 2465 41739 2499
rect 2145 2397 2179 2431
rect 3065 2397 3099 2431
rect 10977 2397 11011 2431
rect 11713 2397 11747 2431
rect 15301 2397 15335 2431
rect 27813 2397 27847 2431
rect 35909 2397 35943 2431
rect 36369 2397 36403 2431
rect 41889 2397 41923 2431
rect 3157 2329 3191 2363
rect 3985 2329 4019 2363
rect 39313 2329 39347 2363
<< metal1 >>
rect 1104 41370 42872 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 42872 41370
rect 1104 41296 42872 41318
rect 2225 41191 2283 41197
rect 2225 41157 2237 41191
rect 2271 41188 2283 41191
rect 5810 41188 5816 41200
rect 2271 41160 5816 41188
rect 2271 41157 2283 41160
rect 2225 41151 2283 41157
rect 5810 41148 5816 41160
rect 5868 41148 5874 41200
rect 7926 41188 7932 41200
rect 7887 41160 7932 41188
rect 7926 41148 7932 41160
rect 7984 41148 7990 41200
rect 24486 41148 24492 41200
rect 24544 41188 24550 41200
rect 24857 41191 24915 41197
rect 24857 41188 24869 41191
rect 24544 41160 24869 41188
rect 24544 41148 24550 41160
rect 24857 41157 24869 41160
rect 24903 41157 24915 41191
rect 24857 41151 24915 41157
rect 34514 41148 34520 41200
rect 34572 41188 34578 41200
rect 34885 41191 34943 41197
rect 34885 41188 34897 41191
rect 34572 41160 34897 41188
rect 34572 41148 34578 41160
rect 34885 41157 34897 41160
rect 34931 41157 34943 41191
rect 34885 41151 34943 41157
rect 41877 41191 41935 41197
rect 41877 41157 41889 41191
rect 41923 41188 41935 41191
rect 42518 41188 42524 41200
rect 41923 41160 42524 41188
rect 41923 41157 41935 41160
rect 41877 41151 41935 41157
rect 42518 41148 42524 41160
rect 42576 41148 42582 41200
rect 1854 41120 1860 41132
rect 1815 41092 1860 41120
rect 1854 41080 1860 41092
rect 1912 41080 1918 41132
rect 2869 41123 2927 41129
rect 2869 41089 2881 41123
rect 2915 41120 2927 41123
rect 3694 41120 3700 41132
rect 2915 41092 3700 41120
rect 2915 41089 2927 41092
rect 2869 41083 2927 41089
rect 3694 41080 3700 41092
rect 3752 41080 3758 41132
rect 3786 41052 3792 41064
rect 3747 41024 3792 41052
rect 3786 41012 3792 41024
rect 3844 41012 3850 41064
rect 3973 41055 4031 41061
rect 3973 41021 3985 41055
rect 4019 41052 4031 41055
rect 4706 41052 4712 41064
rect 4019 41024 4712 41052
rect 4019 41021 4031 41024
rect 3973 41015 4031 41021
rect 4706 41012 4712 41024
rect 4764 41012 4770 41064
rect 4801 41055 4859 41061
rect 4801 41021 4813 41055
rect 4847 41021 4859 41055
rect 12894 41052 12900 41064
rect 12855 41024 12900 41052
rect 4801 41015 4859 41021
rect 2682 40944 2688 40996
rect 2740 40984 2746 40996
rect 4816 40984 4844 41015
rect 12894 41012 12900 41024
rect 12952 41012 12958 41064
rect 12986 41012 12992 41064
rect 13044 41052 13050 41064
rect 13357 41055 13415 41061
rect 13357 41052 13369 41055
rect 13044 41024 13369 41052
rect 13044 41012 13050 41024
rect 13357 41021 13369 41024
rect 13403 41021 13415 41055
rect 13538 41052 13544 41064
rect 13499 41024 13544 41052
rect 13357 41015 13415 41021
rect 13538 41012 13544 41024
rect 13596 41012 13602 41064
rect 21818 41052 21824 41064
rect 21779 41024 21824 41052
rect 21818 41012 21824 41024
rect 21876 41012 21882 41064
rect 22002 41052 22008 41064
rect 21963 41024 22008 41052
rect 22002 41012 22008 41024
rect 22060 41012 22066 41064
rect 22281 41055 22339 41061
rect 22281 41021 22293 41055
rect 22327 41021 22339 41055
rect 22281 41015 22339 41021
rect 33873 41055 33931 41061
rect 33873 41021 33885 41055
rect 33919 41052 33931 41055
rect 34701 41055 34759 41061
rect 34701 41052 34713 41055
rect 33919 41024 34713 41052
rect 33919 41021 33931 41024
rect 33873 41015 33931 41021
rect 34701 41021 34713 41024
rect 34747 41021 34759 41055
rect 34701 41015 34759 41021
rect 35161 41055 35219 41061
rect 35161 41021 35173 41055
rect 35207 41021 35219 41055
rect 35161 41015 35219 41021
rect 40037 41055 40095 41061
rect 40037 41021 40049 41055
rect 40083 41021 40095 41055
rect 40037 41015 40095 41021
rect 40221 41055 40279 41061
rect 40221 41021 40233 41055
rect 40267 41052 40279 41055
rect 41138 41052 41144 41064
rect 40267 41024 41144 41052
rect 40267 41021 40279 41024
rect 40221 41015 40279 41021
rect 2740 40956 4844 40984
rect 2740 40944 2746 40956
rect 21910 40944 21916 40996
rect 21968 40984 21974 40996
rect 22296 40984 22324 41015
rect 21968 40956 22324 40984
rect 21968 40944 21974 40956
rect 34146 40944 34152 40996
rect 34204 40984 34210 40996
rect 35176 40984 35204 41015
rect 34204 40956 35204 40984
rect 40052 40984 40080 41015
rect 41138 41012 41144 41024
rect 41196 41012 41202 41064
rect 40126 40984 40132 40996
rect 40052 40956 40132 40984
rect 34204 40944 34210 40956
rect 40126 40944 40132 40956
rect 40184 40944 40190 40996
rect 2774 40916 2780 40928
rect 2735 40888 2780 40916
rect 2774 40876 2780 40888
rect 2832 40876 2838 40928
rect 8018 40916 8024 40928
rect 7979 40888 8024 40916
rect 8018 40876 8024 40888
rect 8076 40876 8082 40928
rect 10962 40916 10968 40928
rect 10923 40888 10968 40916
rect 10962 40876 10968 40888
rect 11020 40876 11026 40928
rect 14090 40916 14096 40928
rect 14051 40888 14096 40916
rect 14090 40876 14096 40888
rect 14148 40876 14154 40928
rect 14734 40916 14740 40928
rect 14695 40888 14740 40916
rect 14734 40876 14740 40888
rect 14792 40876 14798 40928
rect 20162 40916 20168 40928
rect 20123 40888 20168 40916
rect 20162 40876 20168 40888
rect 20220 40876 20226 40928
rect 24946 40916 24952 40928
rect 24907 40888 24952 40916
rect 24946 40876 24952 40888
rect 25004 40876 25010 40928
rect 26053 40919 26111 40925
rect 26053 40885 26065 40919
rect 26099 40916 26111 40919
rect 26694 40916 26700 40928
rect 26099 40888 26700 40916
rect 26099 40885 26111 40888
rect 26053 40879 26111 40885
rect 26694 40876 26700 40888
rect 26752 40876 26758 40928
rect 26970 40916 26976 40928
rect 26931 40888 26976 40916
rect 26970 40876 26976 40888
rect 27028 40876 27034 40928
rect 29546 40916 29552 40928
rect 29507 40888 29552 40916
rect 29546 40876 29552 40888
rect 29604 40876 29610 40928
rect 31573 40919 31631 40925
rect 31573 40885 31585 40919
rect 31619 40916 31631 40919
rect 32122 40916 32128 40928
rect 31619 40888 32128 40916
rect 31619 40885 31631 40888
rect 31573 40879 31631 40885
rect 32122 40876 32128 40888
rect 32180 40876 32186 40928
rect 32306 40876 32312 40928
rect 32364 40916 32370 40928
rect 32585 40919 32643 40925
rect 32585 40916 32597 40919
rect 32364 40888 32597 40916
rect 32364 40876 32370 40888
rect 32585 40885 32597 40888
rect 32631 40885 32643 40919
rect 32585 40879 32643 40885
rect 37458 40876 37464 40928
rect 37516 40916 37522 40928
rect 38473 40919 38531 40925
rect 38473 40916 38485 40919
rect 37516 40888 38485 40916
rect 37516 40876 37522 40888
rect 38473 40885 38485 40888
rect 38519 40885 38531 40919
rect 38473 40879 38531 40885
rect 39301 40919 39359 40925
rect 39301 40885 39313 40919
rect 39347 40916 39359 40919
rect 40034 40916 40040 40928
rect 39347 40888 40040 40916
rect 39347 40885 39359 40888
rect 39301 40879 39359 40885
rect 40034 40876 40040 40888
rect 40092 40876 40098 40928
rect 1104 40826 42872 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 42872 40826
rect 1104 40752 42872 40774
rect 21818 40672 21824 40724
rect 21876 40712 21882 40724
rect 22465 40715 22523 40721
rect 22465 40712 22477 40715
rect 21876 40684 22477 40712
rect 21876 40672 21882 40684
rect 22465 40681 22477 40684
rect 22511 40681 22523 40715
rect 22465 40675 22523 40681
rect 9861 40647 9919 40653
rect 9861 40613 9873 40647
rect 9907 40644 9919 40647
rect 13354 40644 13360 40656
rect 9907 40616 13360 40644
rect 9907 40613 9919 40616
rect 9861 40607 9919 40613
rect 13354 40604 13360 40616
rect 13412 40604 13418 40656
rect 26418 40604 26424 40656
rect 26476 40644 26482 40656
rect 26476 40616 27200 40644
rect 26476 40604 26482 40616
rect 2038 40576 2044 40588
rect 1999 40548 2044 40576
rect 2038 40536 2044 40548
rect 2096 40536 2102 40588
rect 4890 40536 4896 40588
rect 4948 40576 4954 40588
rect 5169 40579 5227 40585
rect 5169 40576 5181 40579
rect 4948 40548 5181 40576
rect 4948 40536 4954 40548
rect 5169 40545 5181 40548
rect 5215 40545 5227 40579
rect 10962 40576 10968 40588
rect 10923 40548 10968 40576
rect 5169 40539 5227 40545
rect 10962 40536 10968 40548
rect 11020 40536 11026 40588
rect 11606 40576 11612 40588
rect 11567 40548 11612 40576
rect 11606 40536 11612 40548
rect 11664 40536 11670 40588
rect 14090 40576 14096 40588
rect 14051 40548 14096 40576
rect 14090 40536 14096 40548
rect 14148 40536 14154 40588
rect 14274 40536 14280 40588
rect 14332 40576 14338 40588
rect 14553 40579 14611 40585
rect 14553 40576 14565 40579
rect 14332 40548 14565 40576
rect 14332 40536 14338 40548
rect 14553 40545 14565 40548
rect 14599 40545 14611 40579
rect 20162 40576 20168 40588
rect 20123 40548 20168 40576
rect 14553 40539 14611 40545
rect 20162 40536 20168 40548
rect 20220 40536 20226 40588
rect 20714 40576 20720 40588
rect 20675 40548 20720 40576
rect 20714 40536 20720 40548
rect 20772 40536 20778 40588
rect 23474 40536 23480 40588
rect 23532 40576 23538 40588
rect 24857 40579 24915 40585
rect 24857 40576 24869 40579
rect 23532 40548 24869 40576
rect 23532 40536 23538 40548
rect 24857 40545 24869 40548
rect 24903 40545 24915 40579
rect 26694 40576 26700 40588
rect 26655 40548 26700 40576
rect 24857 40539 24915 40545
rect 26694 40536 26700 40548
rect 26752 40536 26758 40588
rect 27172 40585 27200 40616
rect 27157 40579 27215 40585
rect 27157 40545 27169 40579
rect 27203 40545 27215 40579
rect 29546 40576 29552 40588
rect 29507 40548 29552 40576
rect 27157 40539 27215 40545
rect 29546 40536 29552 40548
rect 29604 40536 29610 40588
rect 30006 40576 30012 40588
rect 29967 40548 30012 40576
rect 30006 40536 30012 40548
rect 30064 40536 30070 40588
rect 32306 40576 32312 40588
rect 32267 40548 32312 40576
rect 32306 40536 32312 40548
rect 32364 40536 32370 40588
rect 32858 40576 32864 40588
rect 32819 40548 32864 40576
rect 32858 40536 32864 40548
rect 32916 40536 32922 40588
rect 36078 40576 36084 40588
rect 36039 40548 36084 40576
rect 36078 40536 36084 40548
rect 36136 40536 36142 40588
rect 37458 40576 37464 40588
rect 37419 40548 37464 40576
rect 37458 40536 37464 40548
rect 37516 40536 37522 40588
rect 39298 40576 39304 40588
rect 39259 40548 39304 40576
rect 39298 40536 39304 40548
rect 39356 40536 39362 40588
rect 41874 40576 41880 40588
rect 41835 40548 41880 40576
rect 41874 40536 41880 40548
rect 41932 40536 41938 40588
rect 3234 40468 3240 40520
rect 3292 40508 3298 40520
rect 4249 40511 4307 40517
rect 3292 40480 3337 40508
rect 3292 40468 3298 40480
rect 4249 40477 4261 40511
rect 4295 40508 4307 40511
rect 4709 40511 4767 40517
rect 4709 40508 4721 40511
rect 4295 40480 4721 40508
rect 4295 40477 4307 40480
rect 4249 40471 4307 40477
rect 4709 40477 4721 40480
rect 4755 40477 4767 40511
rect 4709 40471 4767 40477
rect 9122 40468 9128 40520
rect 9180 40508 9186 40520
rect 9217 40511 9275 40517
rect 9217 40508 9229 40511
rect 9180 40480 9229 40508
rect 9180 40468 9186 40480
rect 9217 40477 9229 40480
rect 9263 40477 9275 40511
rect 9217 40471 9275 40477
rect 10321 40511 10379 40517
rect 10321 40477 10333 40511
rect 10367 40477 10379 40511
rect 10321 40471 10379 40477
rect 3050 40440 3056 40452
rect 3011 40412 3056 40440
rect 3050 40400 3056 40412
rect 3108 40400 3114 40452
rect 4893 40443 4951 40449
rect 4893 40409 4905 40443
rect 4939 40440 4951 40443
rect 5626 40440 5632 40452
rect 4939 40412 5632 40440
rect 4939 40409 4951 40412
rect 4893 40403 4951 40409
rect 5626 40400 5632 40412
rect 5684 40400 5690 40452
rect 10336 40372 10364 40471
rect 13170 40468 13176 40520
rect 13228 40508 13234 40520
rect 13357 40511 13415 40517
rect 13357 40508 13369 40511
rect 13228 40480 13369 40508
rect 13228 40468 13234 40480
rect 13357 40477 13369 40480
rect 13403 40477 13415 40511
rect 13357 40471 13415 40477
rect 23293 40511 23351 40517
rect 23293 40477 23305 40511
rect 23339 40508 23351 40511
rect 24397 40511 24455 40517
rect 24397 40508 24409 40511
rect 23339 40480 24409 40508
rect 23339 40477 23351 40480
rect 23293 40471 23351 40477
rect 24397 40477 24409 40480
rect 24443 40477 24455 40511
rect 24397 40471 24455 40477
rect 36998 40468 37004 40520
rect 37056 40508 37062 40520
rect 40310 40508 40316 40520
rect 37056 40480 37101 40508
rect 40271 40480 40316 40508
rect 37056 40468 37062 40480
rect 40310 40468 40316 40480
rect 40368 40468 40374 40520
rect 10413 40443 10471 40449
rect 10413 40409 10425 40443
rect 10459 40440 10471 40443
rect 11149 40443 11207 40449
rect 11149 40440 11161 40443
rect 10459 40412 11161 40440
rect 10459 40409 10471 40412
rect 10413 40403 10471 40409
rect 11149 40409 11161 40412
rect 11195 40409 11207 40443
rect 14274 40440 14280 40452
rect 14235 40412 14280 40440
rect 11149 40403 11207 40409
rect 14274 40400 14280 40412
rect 14332 40400 14338 40452
rect 20346 40440 20352 40452
rect 20307 40412 20352 40440
rect 20346 40400 20352 40412
rect 20404 40400 20410 40452
rect 24578 40440 24584 40452
rect 24539 40412 24584 40440
rect 24578 40400 24584 40412
rect 24636 40400 24642 40452
rect 26326 40400 26332 40452
rect 26384 40440 26390 40452
rect 26881 40443 26939 40449
rect 26881 40440 26893 40443
rect 26384 40412 26893 40440
rect 26384 40400 26390 40412
rect 26881 40409 26893 40412
rect 26927 40409 26939 40443
rect 29730 40440 29736 40452
rect 29691 40412 29736 40440
rect 26881 40403 26939 40409
rect 29730 40400 29736 40412
rect 29788 40400 29794 40452
rect 32490 40440 32496 40452
rect 32451 40412 32496 40440
rect 32490 40400 32496 40412
rect 32548 40400 32554 40452
rect 35894 40400 35900 40452
rect 35952 40440 35958 40452
rect 36817 40443 36875 40449
rect 36817 40440 36829 40443
rect 35952 40412 36829 40440
rect 35952 40400 35958 40412
rect 36817 40409 36829 40412
rect 36863 40409 36875 40443
rect 37642 40440 37648 40452
rect 37603 40412 37648 40440
rect 36817 40403 36875 40409
rect 37642 40400 37648 40412
rect 37700 40400 37706 40452
rect 40494 40440 40500 40452
rect 40455 40412 40500 40440
rect 40494 40400 40500 40412
rect 40552 40400 40558 40452
rect 13170 40372 13176 40384
rect 10336 40344 13176 40372
rect 13170 40332 13176 40344
rect 13228 40332 13234 40384
rect 13446 40372 13452 40384
rect 13407 40344 13452 40372
rect 13446 40332 13452 40344
rect 13504 40332 13510 40384
rect 1104 40282 42872 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 42872 40282
rect 1104 40208 42872 40230
rect 3050 40128 3056 40180
rect 3108 40168 3114 40180
rect 4065 40171 4123 40177
rect 4065 40168 4077 40171
rect 3108 40140 4077 40168
rect 3108 40128 3114 40140
rect 4065 40137 4077 40140
rect 4111 40137 4123 40171
rect 20346 40168 20352 40180
rect 20307 40140 20352 40168
rect 4065 40131 4123 40137
rect 20346 40128 20352 40140
rect 20404 40128 20410 40180
rect 21913 40171 21971 40177
rect 21913 40137 21925 40171
rect 21959 40168 21971 40171
rect 22002 40168 22008 40180
rect 21959 40140 22008 40168
rect 21959 40137 21971 40140
rect 21913 40131 21971 40137
rect 22002 40128 22008 40140
rect 22060 40128 22066 40180
rect 29365 40171 29423 40177
rect 29365 40137 29377 40171
rect 29411 40168 29423 40171
rect 29730 40168 29736 40180
rect 29411 40140 29736 40168
rect 29411 40137 29423 40140
rect 29365 40131 29423 40137
rect 29730 40128 29736 40140
rect 29788 40128 29794 40180
rect 37642 40128 37648 40180
rect 37700 40168 37706 40180
rect 38289 40171 38347 40177
rect 38289 40168 38301 40171
rect 37700 40140 38301 40168
rect 37700 40128 37706 40140
rect 38289 40137 38301 40140
rect 38335 40137 38347 40171
rect 38289 40131 38347 40137
rect 41322 40128 41328 40180
rect 41380 40128 41386 40180
rect 1857 40103 1915 40109
rect 1857 40069 1869 40103
rect 1903 40100 1915 40103
rect 2774 40100 2780 40112
rect 1903 40072 2780 40100
rect 1903 40069 1915 40072
rect 1857 40063 1915 40069
rect 2774 40060 2780 40072
rect 2832 40060 2838 40112
rect 3510 40100 3516 40112
rect 3471 40072 3516 40100
rect 3510 40060 3516 40072
rect 3568 40060 3574 40112
rect 3694 40060 3700 40112
rect 3752 40100 3758 40112
rect 7190 40100 7196 40112
rect 3752 40072 7196 40100
rect 3752 40060 3758 40072
rect 7190 40060 7196 40072
rect 7248 40100 7254 40112
rect 8202 40100 8208 40112
rect 7248 40072 8208 40100
rect 7248 40060 7254 40072
rect 8202 40060 8208 40072
rect 8260 40060 8266 40112
rect 13446 40060 13452 40112
rect 13504 40100 13510 40112
rect 14277 40103 14335 40109
rect 14277 40100 14289 40103
rect 13504 40072 14289 40100
rect 13504 40060 13510 40072
rect 14277 40069 14289 40072
rect 14323 40069 14335 40103
rect 32309 40103 32367 40109
rect 32309 40100 32321 40103
rect 14277 40063 14335 40069
rect 31726 40072 32321 40100
rect 4157 40035 4215 40041
rect 4157 40001 4169 40035
rect 4203 40001 4215 40035
rect 4706 40032 4712 40044
rect 4667 40004 4712 40032
rect 4157 39995 4215 40001
rect 1578 39924 1584 39976
rect 1636 39964 1642 39976
rect 1673 39967 1731 39973
rect 1673 39964 1685 39967
rect 1636 39936 1685 39964
rect 1636 39924 1642 39936
rect 1673 39933 1685 39936
rect 1719 39933 1731 39967
rect 1673 39927 1731 39933
rect 4172 39896 4200 39995
rect 4706 39992 4712 40004
rect 4764 39992 4770 40044
rect 4801 40035 4859 40041
rect 4801 40001 4813 40035
rect 4847 40001 4859 40035
rect 5626 40032 5632 40044
rect 5587 40004 5632 40032
rect 4801 39995 4859 40001
rect 4614 39924 4620 39976
rect 4672 39964 4678 39976
rect 4816 39964 4844 39995
rect 5626 39992 5632 40004
rect 5684 39992 5690 40044
rect 5721 40035 5779 40041
rect 5721 40001 5733 40035
rect 5767 40032 5779 40035
rect 6730 40032 6736 40044
rect 5767 40004 6736 40032
rect 5767 40001 5779 40004
rect 5721 39995 5779 40001
rect 6730 39992 6736 40004
rect 6788 39992 6794 40044
rect 9122 40032 9128 40044
rect 9083 40004 9128 40032
rect 9122 39992 9128 40004
rect 9180 39992 9186 40044
rect 20254 40032 20260 40044
rect 20215 40004 20260 40032
rect 20254 39992 20260 40004
rect 20312 39992 20318 40044
rect 21634 39992 21640 40044
rect 21692 40032 21698 40044
rect 21821 40035 21879 40041
rect 21821 40032 21833 40035
rect 21692 40004 21833 40032
rect 21692 39992 21698 40004
rect 21821 40001 21833 40004
rect 21867 40001 21879 40035
rect 25958 40032 25964 40044
rect 25919 40004 25964 40032
rect 21821 39995 21879 40001
rect 25958 39992 25964 40004
rect 26016 39992 26022 40044
rect 26053 40035 26111 40041
rect 26053 40001 26065 40035
rect 26099 40032 26111 40035
rect 26326 40032 26332 40044
rect 26099 40004 26332 40032
rect 26099 40001 26111 40004
rect 26053 39995 26111 40001
rect 26326 39992 26332 40004
rect 26384 39992 26390 40044
rect 26970 40032 26976 40044
rect 26931 40004 26976 40032
rect 26970 39992 26976 40004
rect 27028 39992 27034 40044
rect 29270 40032 29276 40044
rect 29231 40004 29276 40032
rect 29270 39992 29276 40004
rect 29328 39992 29334 40044
rect 31386 40032 31392 40044
rect 31347 40004 31392 40032
rect 31386 39992 31392 40004
rect 31444 39992 31450 40044
rect 31481 40035 31539 40041
rect 31481 40001 31493 40035
rect 31527 40032 31539 40035
rect 31726 40032 31754 40072
rect 32309 40069 32321 40072
rect 32355 40069 32367 40103
rect 32309 40063 32367 40069
rect 34790 40060 34796 40112
rect 34848 40100 34854 40112
rect 35069 40103 35127 40109
rect 35069 40100 35081 40103
rect 34848 40072 35081 40100
rect 34848 40060 34854 40072
rect 35069 40069 35081 40072
rect 35115 40069 35127 40103
rect 35069 40063 35127 40069
rect 36725 40103 36783 40109
rect 36725 40069 36737 40103
rect 36771 40100 36783 40103
rect 39298 40100 39304 40112
rect 36771 40072 39304 40100
rect 36771 40069 36783 40072
rect 36725 40063 36783 40069
rect 39298 40060 39304 40072
rect 39356 40060 39362 40112
rect 41340 40100 41368 40128
rect 41877 40103 41935 40109
rect 41877 40100 41889 40103
rect 41340 40072 41889 40100
rect 41877 40069 41889 40072
rect 41923 40069 41935 40103
rect 41877 40063 41935 40069
rect 32122 40032 32128 40044
rect 31527 40004 31754 40032
rect 32083 40004 32128 40032
rect 31527 40001 31539 40004
rect 31481 39995 31539 40001
rect 32122 39992 32128 40004
rect 32180 39992 32186 40044
rect 38194 40032 38200 40044
rect 38155 40004 38200 40032
rect 38194 39992 38200 40004
rect 38252 39992 38258 40044
rect 40034 40032 40040 40044
rect 39995 40004 40040 40032
rect 40034 39992 40040 40004
rect 40092 39992 40098 40044
rect 9306 39964 9312 39976
rect 4672 39936 4844 39964
rect 9267 39936 9312 39964
rect 4672 39924 4678 39936
rect 9306 39924 9312 39936
rect 9364 39924 9370 39976
rect 9674 39964 9680 39976
rect 9635 39936 9680 39964
rect 9674 39924 9680 39936
rect 9732 39924 9738 39976
rect 12250 39964 12256 39976
rect 12211 39936 12256 39964
rect 12250 39924 12256 39936
rect 12308 39924 12314 39976
rect 13262 39964 13268 39976
rect 13223 39936 13268 39964
rect 13262 39924 13268 39936
rect 13320 39924 13326 39976
rect 13446 39964 13452 39976
rect 13407 39936 13452 39964
rect 13446 39924 13452 39936
rect 13504 39924 13510 39976
rect 14093 39967 14151 39973
rect 14093 39933 14105 39967
rect 14139 39964 14151 39967
rect 14734 39964 14740 39976
rect 14139 39936 14740 39964
rect 14139 39933 14151 39936
rect 14093 39927 14151 39933
rect 14734 39924 14740 39936
rect 14792 39924 14798 39976
rect 15930 39964 15936 39976
rect 15891 39936 15936 39964
rect 15930 39924 15936 39936
rect 15988 39924 15994 39976
rect 23290 39964 23296 39976
rect 23251 39936 23296 39964
rect 23290 39924 23296 39936
rect 23348 39924 23354 39976
rect 23474 39964 23480 39976
rect 23435 39936 23480 39964
rect 23474 39924 23480 39936
rect 23532 39924 23538 39976
rect 23842 39964 23848 39976
rect 23803 39936 23848 39964
rect 23842 39924 23848 39936
rect 23900 39924 23906 39976
rect 27154 39964 27160 39976
rect 27115 39936 27160 39964
rect 27154 39924 27160 39936
rect 27212 39924 27218 39976
rect 27338 39924 27344 39976
rect 27396 39964 27402 39976
rect 27433 39967 27491 39973
rect 27433 39964 27445 39967
rect 27396 39936 27445 39964
rect 27396 39924 27402 39936
rect 27433 39933 27445 39936
rect 27479 39933 27491 39967
rect 27433 39927 27491 39933
rect 32398 39924 32404 39976
rect 32456 39964 32462 39976
rect 32585 39967 32643 39973
rect 32585 39964 32597 39967
rect 32456 39936 32597 39964
rect 32456 39924 32462 39936
rect 32585 39933 32597 39936
rect 32631 39933 32643 39967
rect 32585 39927 32643 39933
rect 34885 39967 34943 39973
rect 34885 39933 34897 39967
rect 34931 39964 34943 39967
rect 35342 39964 35348 39976
rect 34931 39936 35348 39964
rect 34931 39933 34943 39936
rect 34885 39927 34943 39933
rect 35342 39924 35348 39936
rect 35400 39924 35406 39976
rect 40221 39967 40279 39973
rect 40221 39933 40233 39967
rect 40267 39964 40279 39967
rect 41966 39964 41972 39976
rect 40267 39936 41972 39964
rect 40267 39933 40279 39936
rect 40221 39927 40279 39933
rect 41966 39924 41972 39936
rect 42024 39924 42030 39976
rect 4982 39896 4988 39908
rect 4172 39868 4988 39896
rect 4982 39856 4988 39868
rect 5040 39896 5046 39908
rect 12434 39896 12440 39908
rect 5040 39868 12440 39896
rect 5040 39856 5046 39868
rect 12434 39856 12440 39868
rect 12492 39856 12498 39908
rect 20254 39856 20260 39908
rect 20312 39896 20318 39908
rect 20312 39868 41414 39896
rect 20312 39856 20318 39868
rect 41386 39840 41414 39868
rect 6365 39831 6423 39837
rect 6365 39797 6377 39831
rect 6411 39828 6423 39831
rect 6454 39828 6460 39840
rect 6411 39800 6460 39828
rect 6411 39797 6423 39800
rect 6365 39791 6423 39797
rect 6454 39788 6460 39800
rect 6512 39788 6518 39840
rect 39577 39831 39635 39837
rect 39577 39797 39589 39831
rect 39623 39828 39635 39831
rect 40310 39828 40316 39840
rect 39623 39800 40316 39828
rect 39623 39797 39635 39800
rect 39577 39791 39635 39797
rect 40310 39788 40316 39800
rect 40368 39788 40374 39840
rect 41386 39800 41420 39840
rect 41414 39788 41420 39800
rect 41472 39788 41478 39840
rect 1104 39738 42872 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 42872 39738
rect 1104 39664 42872 39686
rect 3234 39584 3240 39636
rect 3292 39624 3298 39636
rect 3789 39627 3847 39633
rect 3789 39624 3801 39627
rect 3292 39596 3801 39624
rect 3292 39584 3298 39596
rect 3789 39593 3801 39596
rect 3835 39593 3847 39627
rect 9306 39624 9312 39636
rect 9267 39596 9312 39624
rect 3789 39587 3847 39593
rect 9306 39584 9312 39596
rect 9364 39584 9370 39636
rect 12529 39627 12587 39633
rect 12529 39593 12541 39627
rect 12575 39624 12587 39627
rect 12986 39624 12992 39636
rect 12575 39596 12992 39624
rect 12575 39593 12587 39596
rect 12529 39587 12587 39593
rect 12986 39584 12992 39596
rect 13044 39584 13050 39636
rect 13173 39627 13231 39633
rect 13173 39593 13185 39627
rect 13219 39624 13231 39627
rect 13262 39624 13268 39636
rect 13219 39596 13268 39624
rect 13219 39593 13231 39596
rect 13173 39587 13231 39593
rect 13262 39584 13268 39596
rect 13320 39584 13326 39636
rect 14185 39627 14243 39633
rect 14185 39593 14197 39627
rect 14231 39624 14243 39627
rect 14274 39624 14280 39636
rect 14231 39596 14280 39624
rect 14231 39593 14243 39596
rect 14185 39587 14243 39593
rect 14274 39584 14280 39596
rect 14332 39584 14338 39636
rect 23290 39584 23296 39636
rect 23348 39624 23354 39636
rect 23385 39627 23443 39633
rect 23385 39624 23397 39627
rect 23348 39596 23397 39624
rect 23348 39584 23354 39596
rect 23385 39593 23397 39596
rect 23431 39593 23443 39627
rect 23385 39587 23443 39593
rect 26697 39627 26755 39633
rect 26697 39593 26709 39627
rect 26743 39624 26755 39627
rect 27154 39624 27160 39636
rect 26743 39596 27160 39624
rect 26743 39593 26755 39596
rect 26697 39587 26755 39593
rect 27154 39584 27160 39596
rect 27212 39584 27218 39636
rect 32490 39584 32496 39636
rect 32548 39624 32554 39636
rect 32769 39627 32827 39633
rect 32769 39624 32781 39627
rect 32548 39596 32781 39624
rect 32548 39584 32554 39596
rect 32769 39593 32781 39596
rect 32815 39593 32827 39627
rect 32769 39587 32827 39593
rect 33965 39627 34023 39633
rect 33965 39593 33977 39627
rect 34011 39624 34023 39627
rect 34514 39624 34520 39636
rect 34011 39596 34520 39624
rect 34011 39593 34023 39596
rect 33965 39587 34023 39593
rect 34514 39584 34520 39596
rect 34572 39584 34578 39636
rect 34790 39624 34796 39636
rect 34751 39596 34796 39624
rect 34790 39584 34796 39596
rect 34848 39584 34854 39636
rect 35805 39627 35863 39633
rect 35805 39593 35817 39627
rect 35851 39624 35863 39627
rect 35894 39624 35900 39636
rect 35851 39596 35900 39624
rect 35851 39593 35863 39596
rect 35805 39587 35863 39593
rect 35894 39584 35900 39596
rect 35952 39584 35958 39636
rect 36541 39627 36599 39633
rect 36541 39593 36553 39627
rect 36587 39624 36599 39627
rect 36998 39624 37004 39636
rect 36587 39596 37004 39624
rect 36587 39593 36599 39596
rect 36541 39587 36599 39593
rect 36998 39584 37004 39596
rect 37056 39584 37062 39636
rect 40037 39627 40095 39633
rect 40037 39593 40049 39627
rect 40083 39624 40095 39627
rect 40494 39624 40500 39636
rect 40083 39596 40500 39624
rect 40083 39593 40095 39596
rect 40037 39587 40095 39593
rect 40494 39584 40500 39596
rect 40552 39584 40558 39636
rect 41138 39584 41144 39636
rect 41196 39624 41202 39636
rect 41325 39627 41383 39633
rect 41325 39624 41337 39627
rect 41196 39596 41337 39624
rect 41196 39584 41202 39596
rect 41325 39593 41337 39596
rect 41371 39593 41383 39627
rect 41966 39624 41972 39636
rect 41927 39596 41972 39624
rect 41325 39587 41383 39593
rect 41966 39584 41972 39596
rect 42024 39584 42030 39636
rect 4614 39516 4620 39568
rect 4672 39556 4678 39568
rect 14090 39556 14096 39568
rect 4672 39528 14096 39556
rect 4672 39516 4678 39528
rect 14090 39516 14096 39528
rect 14148 39516 14154 39568
rect 15930 39516 15936 39568
rect 15988 39556 15994 39568
rect 36722 39556 36728 39568
rect 15988 39528 36728 39556
rect 15988 39516 15994 39528
rect 36722 39516 36728 39528
rect 36780 39516 36786 39568
rect 39301 39559 39359 39565
rect 39301 39525 39313 39559
rect 39347 39556 39359 39559
rect 40126 39556 40132 39568
rect 39347 39528 40132 39556
rect 39347 39525 39359 39528
rect 39301 39519 39359 39525
rect 40126 39516 40132 39528
rect 40184 39516 40190 39568
rect 2866 39488 2872 39500
rect 2827 39460 2872 39488
rect 2866 39448 2872 39460
rect 2924 39448 2930 39500
rect 5258 39488 5264 39500
rect 5219 39460 5264 39488
rect 5258 39448 5264 39460
rect 5316 39448 5322 39500
rect 6454 39488 6460 39500
rect 6415 39460 6460 39488
rect 6454 39448 6460 39460
rect 6512 39448 6518 39500
rect 6730 39448 6736 39500
rect 6788 39488 6794 39500
rect 6788 39460 33916 39488
rect 6788 39448 6794 39460
rect 1394 39420 1400 39432
rect 1355 39392 1400 39420
rect 1394 39380 1400 39392
rect 1452 39380 1458 39432
rect 9214 39420 9220 39432
rect 9175 39392 9220 39420
rect 9214 39380 9220 39392
rect 9272 39380 9278 39432
rect 10226 39420 10232 39432
rect 10187 39392 10232 39420
rect 10226 39380 10232 39392
rect 10284 39380 10290 39432
rect 10870 39380 10876 39432
rect 10928 39420 10934 39432
rect 11609 39423 11667 39429
rect 11609 39420 11621 39423
rect 10928 39392 11621 39420
rect 10928 39380 10934 39392
rect 11609 39389 11621 39392
rect 11655 39389 11667 39423
rect 11609 39383 11667 39389
rect 12434 39380 12440 39432
rect 12492 39420 12498 39432
rect 13078 39420 13084 39432
rect 12492 39392 12585 39420
rect 12991 39392 13084 39420
rect 12492 39380 12498 39392
rect 13078 39380 13084 39392
rect 13136 39420 13142 39432
rect 14090 39420 14096 39432
rect 13136 39392 13952 39420
rect 14051 39392 14096 39420
rect 13136 39380 13142 39392
rect 1581 39355 1639 39361
rect 1581 39321 1593 39355
rect 1627 39352 1639 39355
rect 2130 39352 2136 39364
rect 1627 39324 2136 39352
rect 1627 39321 1639 39324
rect 1581 39315 1639 39321
rect 2130 39312 2136 39324
rect 2188 39312 2194 39364
rect 4798 39312 4804 39364
rect 4856 39352 4862 39364
rect 6273 39355 6331 39361
rect 6273 39352 6285 39355
rect 4856 39324 6285 39352
rect 4856 39312 4862 39324
rect 6273 39321 6285 39324
rect 6319 39321 6331 39355
rect 6273 39315 6331 39321
rect 8938 39312 8944 39364
rect 8996 39352 9002 39364
rect 11057 39355 11115 39361
rect 11057 39352 11069 39355
rect 8996 39324 11069 39352
rect 8996 39312 9002 39324
rect 11057 39321 11069 39324
rect 11103 39321 11115 39355
rect 11057 39315 11115 39321
rect 10410 39284 10416 39296
rect 10371 39256 10416 39284
rect 10410 39244 10416 39256
rect 10468 39244 10474 39296
rect 12452 39284 12480 39380
rect 13924 39352 13952 39392
rect 14090 39380 14096 39392
rect 14148 39380 14154 39432
rect 22738 39420 22744 39432
rect 22699 39392 22744 39420
rect 22738 39380 22744 39392
rect 22796 39380 22802 39432
rect 22833 39423 22891 39429
rect 22833 39389 22845 39423
rect 22879 39420 22891 39423
rect 24578 39420 24584 39432
rect 22879 39392 24584 39420
rect 22879 39389 22891 39392
rect 22833 39383 22891 39389
rect 24578 39380 24584 39392
rect 24636 39380 24642 39432
rect 26602 39420 26608 39432
rect 26563 39392 26608 39420
rect 26602 39380 26608 39392
rect 26660 39380 26666 39432
rect 32858 39420 32864 39432
rect 32819 39392 32864 39420
rect 32858 39380 32864 39392
rect 32916 39380 32922 39432
rect 33888 39429 33916 39460
rect 33873 39423 33931 39429
rect 33873 39389 33885 39423
rect 33919 39420 33931 39423
rect 34701 39423 34759 39429
rect 34701 39420 34713 39423
rect 33919 39392 34713 39420
rect 33919 39389 33931 39392
rect 33873 39383 33931 39389
rect 34701 39389 34713 39392
rect 34747 39389 34759 39423
rect 35894 39420 35900 39432
rect 35855 39392 35900 39420
rect 34701 39383 34759 39389
rect 35894 39380 35900 39392
rect 35952 39380 35958 39432
rect 39758 39380 39764 39432
rect 39816 39420 39822 39432
rect 39945 39423 40003 39429
rect 39945 39420 39957 39423
rect 39816 39392 39957 39420
rect 39816 39380 39822 39392
rect 39945 39389 39957 39392
rect 39991 39389 40003 39423
rect 39945 39383 40003 39389
rect 40773 39423 40831 39429
rect 40773 39389 40785 39423
rect 40819 39420 40831 39423
rect 41230 39420 41236 39432
rect 40819 39392 41236 39420
rect 40819 39389 40831 39392
rect 40773 39383 40831 39389
rect 41230 39380 41236 39392
rect 41288 39380 41294 39432
rect 41414 39420 41420 39432
rect 41375 39392 41420 39420
rect 41414 39380 41420 39392
rect 41472 39380 41478 39432
rect 41877 39423 41935 39429
rect 41877 39389 41889 39423
rect 41923 39389 41935 39423
rect 41877 39383 41935 39389
rect 31386 39352 31392 39364
rect 13924 39324 31392 39352
rect 31386 39312 31392 39324
rect 31444 39312 31450 39364
rect 41892 39352 41920 39383
rect 42242 39352 42248 39364
rect 31726 39324 42248 39352
rect 21634 39284 21640 39296
rect 12452 39256 21640 39284
rect 21634 39244 21640 39256
rect 21692 39244 21698 39296
rect 29270 39244 29276 39296
rect 29328 39284 29334 39296
rect 31726 39284 31754 39324
rect 42242 39312 42248 39324
rect 42300 39312 42306 39364
rect 29328 39256 31754 39284
rect 29328 39244 29334 39256
rect 40218 39244 40224 39296
rect 40276 39284 40282 39296
rect 40681 39287 40739 39293
rect 40681 39284 40693 39287
rect 40276 39256 40693 39284
rect 40276 39244 40282 39256
rect 40681 39253 40693 39256
rect 40727 39253 40739 39287
rect 40681 39247 40739 39253
rect 1104 39194 42872 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 42872 39194
rect 1104 39120 42872 39142
rect 2130 39080 2136 39092
rect 2091 39052 2136 39080
rect 2130 39040 2136 39052
rect 2188 39040 2194 39092
rect 4798 39080 4804 39092
rect 4759 39052 4804 39080
rect 4798 39040 4804 39052
rect 4856 39040 4862 39092
rect 23385 39083 23443 39089
rect 23385 39049 23397 39083
rect 23431 39080 23443 39083
rect 23474 39080 23480 39092
rect 23431 39052 23480 39080
rect 23431 39049 23443 39052
rect 23385 39043 23443 39049
rect 23474 39040 23480 39052
rect 23532 39040 23538 39092
rect 25958 39040 25964 39092
rect 26016 39080 26022 39092
rect 39758 39080 39764 39092
rect 26016 39052 39764 39080
rect 26016 39040 26022 39052
rect 39758 39040 39764 39052
rect 39816 39040 39822 39092
rect 41230 39080 41236 39092
rect 39868 39052 41236 39080
rect 6886 38984 10364 39012
rect 1578 38944 1584 38956
rect 1539 38916 1584 38944
rect 1578 38904 1584 38916
rect 1636 38904 1642 38956
rect 2225 38947 2283 38953
rect 2225 38913 2237 38947
rect 2271 38913 2283 38947
rect 3786 38944 3792 38956
rect 3747 38916 3792 38944
rect 2225 38907 2283 38913
rect 2240 38876 2268 38907
rect 3786 38904 3792 38916
rect 3844 38904 3850 38956
rect 4706 38944 4712 38956
rect 4667 38916 4712 38944
rect 4706 38904 4712 38916
rect 4764 38944 4770 38956
rect 6886 38944 6914 38984
rect 8846 38944 8852 38956
rect 4764 38916 6914 38944
rect 8759 38916 8852 38944
rect 4764 38904 4770 38916
rect 8846 38904 8852 38916
rect 8904 38944 8910 38956
rect 9582 38944 9588 38956
rect 8904 38916 9444 38944
rect 9543 38916 9588 38944
rect 8904 38904 8910 38916
rect 2406 38876 2412 38888
rect 2240 38848 2412 38876
rect 2406 38836 2412 38848
rect 2464 38876 2470 38888
rect 8938 38876 8944 38888
rect 2464 38848 8944 38876
rect 2464 38836 2470 38848
rect 8938 38836 8944 38848
rect 8996 38836 9002 38888
rect 9416 38808 9444 38916
rect 9582 38904 9588 38916
rect 9640 38904 9646 38956
rect 10336 38888 10364 38984
rect 14090 38972 14096 39024
rect 14148 39012 14154 39024
rect 39868 39012 39896 39052
rect 41230 39040 41236 39052
rect 41288 39040 41294 39092
rect 40218 39012 40224 39024
rect 14148 38984 39896 39012
rect 40179 38984 40224 39012
rect 14148 38972 14154 38984
rect 40218 38972 40224 38984
rect 40276 38972 40282 39024
rect 41874 39012 41880 39024
rect 41835 38984 41880 39012
rect 41874 38972 41880 38984
rect 41932 38972 41938 39024
rect 10410 38904 10416 38956
rect 10468 38944 10474 38956
rect 10870 38944 10876 38956
rect 10468 38916 10876 38944
rect 10468 38904 10474 38916
rect 10870 38904 10876 38916
rect 10928 38944 10934 38956
rect 11517 38947 11575 38953
rect 11517 38944 11529 38947
rect 10928 38916 11529 38944
rect 10928 38904 10934 38916
rect 11517 38913 11529 38916
rect 11563 38913 11575 38947
rect 11517 38907 11575 38913
rect 13173 38947 13231 38953
rect 13173 38913 13185 38947
rect 13219 38944 13231 38947
rect 13538 38944 13544 38956
rect 13219 38916 13544 38944
rect 13219 38913 13231 38916
rect 13173 38907 13231 38913
rect 13538 38904 13544 38916
rect 13596 38904 13602 38956
rect 22922 38904 22928 38956
rect 22980 38944 22986 38956
rect 23293 38947 23351 38953
rect 23293 38944 23305 38947
rect 22980 38916 23305 38944
rect 22980 38904 22986 38916
rect 23293 38913 23305 38916
rect 23339 38913 23351 38947
rect 32674 38944 32680 38956
rect 32635 38916 32680 38944
rect 23293 38907 23351 38913
rect 32674 38904 32680 38916
rect 32732 38904 32738 38956
rect 32858 38944 32864 38956
rect 32819 38916 32864 38944
rect 32858 38904 32864 38916
rect 32916 38904 32922 38956
rect 33502 38944 33508 38956
rect 33463 38916 33508 38944
rect 33502 38904 33508 38916
rect 33560 38904 33566 38956
rect 35253 38947 35311 38953
rect 35253 38913 35265 38947
rect 35299 38944 35311 38947
rect 35342 38944 35348 38956
rect 35299 38916 35348 38944
rect 35299 38913 35311 38916
rect 35253 38907 35311 38913
rect 35342 38904 35348 38916
rect 35400 38904 35406 38956
rect 35989 38947 36047 38953
rect 35989 38913 36001 38947
rect 36035 38944 36047 38947
rect 36078 38944 36084 38956
rect 36035 38916 36084 38944
rect 36035 38913 36047 38916
rect 35989 38907 36047 38913
rect 36078 38904 36084 38916
rect 36136 38904 36142 38956
rect 36173 38947 36231 38953
rect 36173 38913 36185 38947
rect 36219 38913 36231 38947
rect 36173 38907 36231 38913
rect 36265 38947 36323 38953
rect 36265 38913 36277 38947
rect 36311 38944 36323 38947
rect 36446 38944 36452 38956
rect 36311 38916 36452 38944
rect 36311 38913 36323 38916
rect 36265 38907 36323 38913
rect 10318 38876 10324 38888
rect 10279 38848 10324 38876
rect 10318 38836 10324 38848
rect 10376 38836 10382 38888
rect 12342 38876 12348 38888
rect 12303 38848 12348 38876
rect 12342 38836 12348 38848
rect 12400 38836 12406 38888
rect 36188 38876 36216 38907
rect 36446 38904 36452 38916
rect 36504 38944 36510 38956
rect 37921 38947 37979 38953
rect 37921 38944 37933 38947
rect 36504 38916 37933 38944
rect 36504 38904 36510 38916
rect 37921 38913 37933 38916
rect 37967 38913 37979 38947
rect 38102 38944 38108 38956
rect 38063 38916 38108 38944
rect 37921 38907 37979 38913
rect 38102 38904 38108 38916
rect 38160 38904 38166 38956
rect 36906 38876 36912 38888
rect 36188 38848 36912 38876
rect 36906 38836 36912 38848
rect 36964 38836 36970 38888
rect 39577 38879 39635 38885
rect 39577 38845 39589 38879
rect 39623 38876 39635 38879
rect 40037 38879 40095 38885
rect 40037 38876 40049 38879
rect 39623 38848 40049 38876
rect 39623 38845 39635 38848
rect 39577 38839 39635 38845
rect 40037 38845 40049 38848
rect 40083 38845 40095 38879
rect 40037 38839 40095 38845
rect 38194 38808 38200 38820
rect 9416 38780 38200 38808
rect 38194 38768 38200 38780
rect 38252 38768 38258 38820
rect 9214 38700 9220 38752
rect 9272 38740 9278 38752
rect 11974 38740 11980 38752
rect 9272 38712 11980 38740
rect 9272 38700 9278 38712
rect 11974 38700 11980 38712
rect 12032 38700 12038 38752
rect 33045 38743 33103 38749
rect 33045 38709 33057 38743
rect 33091 38740 33103 38743
rect 33318 38740 33324 38752
rect 33091 38712 33324 38740
rect 33091 38709 33103 38712
rect 33045 38703 33103 38709
rect 33318 38700 33324 38712
rect 33376 38700 33382 38752
rect 33689 38743 33747 38749
rect 33689 38709 33701 38743
rect 33735 38740 33747 38743
rect 33778 38740 33784 38752
rect 33735 38712 33784 38740
rect 33735 38709 33747 38712
rect 33689 38703 33747 38709
rect 33778 38700 33784 38712
rect 33836 38700 33842 38752
rect 35986 38740 35992 38752
rect 35947 38712 35992 38740
rect 35986 38700 35992 38712
rect 36044 38700 36050 38752
rect 38105 38743 38163 38749
rect 38105 38709 38117 38743
rect 38151 38740 38163 38743
rect 38654 38740 38660 38752
rect 38151 38712 38660 38740
rect 38151 38709 38163 38712
rect 38105 38703 38163 38709
rect 38654 38700 38660 38712
rect 38712 38700 38718 38752
rect 1104 38650 42872 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 42872 38650
rect 1104 38576 42872 38598
rect 1394 38496 1400 38548
rect 1452 38536 1458 38548
rect 1673 38539 1731 38545
rect 1673 38536 1685 38539
rect 1452 38508 1685 38536
rect 1452 38496 1458 38508
rect 1673 38505 1685 38508
rect 1719 38505 1731 38539
rect 1673 38499 1731 38505
rect 30650 38496 30656 38548
rect 30708 38536 30714 38548
rect 30929 38539 30987 38545
rect 30929 38536 30941 38539
rect 30708 38508 30941 38536
rect 30708 38496 30714 38508
rect 30929 38505 30941 38508
rect 30975 38505 30987 38539
rect 36906 38536 36912 38548
rect 36867 38508 36912 38536
rect 30929 38499 30987 38505
rect 36906 38496 36912 38508
rect 36964 38496 36970 38548
rect 31113 38471 31171 38477
rect 31113 38437 31125 38471
rect 31159 38468 31171 38471
rect 32674 38468 32680 38480
rect 31159 38440 32680 38468
rect 31159 38437 31171 38440
rect 31113 38431 31171 38437
rect 32674 38428 32680 38440
rect 32732 38428 32738 38480
rect 9217 38403 9275 38409
rect 9217 38400 9229 38403
rect 6886 38372 9229 38400
rect 2777 38335 2835 38341
rect 2777 38301 2789 38335
rect 2823 38301 2835 38335
rect 2777 38295 2835 38301
rect 3973 38335 4031 38341
rect 3973 38301 3985 38335
rect 4019 38332 4031 38335
rect 6886 38332 6914 38372
rect 9217 38369 9229 38372
rect 9263 38400 9275 38403
rect 20254 38400 20260 38412
rect 9263 38372 20260 38400
rect 9263 38369 9275 38372
rect 9217 38363 9275 38369
rect 20254 38360 20260 38372
rect 20312 38360 20318 38412
rect 25225 38403 25283 38409
rect 25225 38369 25237 38403
rect 25271 38400 25283 38403
rect 25958 38400 25964 38412
rect 25271 38372 25964 38400
rect 25271 38369 25283 38372
rect 25225 38363 25283 38369
rect 25958 38360 25964 38372
rect 26016 38360 26022 38412
rect 31573 38403 31631 38409
rect 31573 38400 31585 38403
rect 30760 38372 31585 38400
rect 4019 38304 6914 38332
rect 4019 38301 4031 38304
rect 3973 38295 4031 38301
rect 2792 38264 2820 38295
rect 8846 38292 8852 38344
rect 8904 38332 8910 38344
rect 8941 38335 8999 38341
rect 8941 38332 8953 38335
rect 8904 38304 8953 38332
rect 8904 38292 8910 38304
rect 8941 38301 8953 38304
rect 8987 38301 8999 38335
rect 10870 38332 10876 38344
rect 10831 38304 10876 38332
rect 8941 38295 8999 38301
rect 10870 38292 10876 38304
rect 10928 38292 10934 38344
rect 24946 38332 24952 38344
rect 24907 38304 24952 38332
rect 24946 38292 24952 38304
rect 25004 38292 25010 38344
rect 25133 38335 25191 38341
rect 25133 38301 25145 38335
rect 25179 38301 25191 38335
rect 25866 38332 25872 38344
rect 25827 38304 25872 38332
rect 25133 38295 25191 38301
rect 4430 38264 4436 38276
rect 2792 38236 4436 38264
rect 4430 38224 4436 38236
rect 4488 38224 4494 38276
rect 11701 38267 11759 38273
rect 11701 38233 11713 38267
rect 11747 38233 11759 38267
rect 25148 38264 25176 38295
rect 25866 38292 25872 38304
rect 25924 38292 25930 38344
rect 26050 38332 26056 38344
rect 26011 38304 26056 38332
rect 26050 38292 26056 38304
rect 26108 38292 26114 38344
rect 30190 38332 30196 38344
rect 30151 38304 30196 38332
rect 30190 38292 30196 38304
rect 30248 38292 30254 38344
rect 25222 38264 25228 38276
rect 25148 38236 25228 38264
rect 11701 38227 11759 38233
rect 3881 38199 3939 38205
rect 3881 38165 3893 38199
rect 3927 38196 3939 38199
rect 4246 38196 4252 38208
rect 3927 38168 4252 38196
rect 3927 38165 3939 38168
rect 3881 38159 3939 38165
rect 4246 38156 4252 38168
rect 4304 38156 4310 38208
rect 11422 38156 11428 38208
rect 11480 38196 11486 38208
rect 11716 38196 11744 38227
rect 25222 38224 25228 38236
rect 25280 38224 25286 38276
rect 30282 38224 30288 38276
rect 30340 38264 30346 38276
rect 30760 38273 30788 38372
rect 31573 38369 31585 38372
rect 31619 38369 31631 38403
rect 41322 38400 41328 38412
rect 41283 38372 41328 38400
rect 31573 38363 31631 38369
rect 41322 38360 41328 38372
rect 41380 38360 41386 38412
rect 31849 38335 31907 38341
rect 31312 38304 31754 38332
rect 30745 38267 30803 38273
rect 30745 38264 30757 38267
rect 30340 38236 30757 38264
rect 30340 38224 30346 38236
rect 30745 38233 30757 38236
rect 30791 38233 30803 38267
rect 30745 38227 30803 38233
rect 30961 38267 31019 38273
rect 30961 38233 30973 38267
rect 31007 38264 31019 38267
rect 31312 38264 31340 38304
rect 31726 38276 31754 38304
rect 31849 38301 31861 38335
rect 31895 38332 31907 38335
rect 32858 38332 32864 38344
rect 31895 38304 32864 38332
rect 31895 38301 31907 38304
rect 31849 38295 31907 38301
rect 32858 38292 32864 38304
rect 32916 38292 32922 38344
rect 33778 38292 33784 38344
rect 33836 38341 33842 38344
rect 33836 38332 33848 38341
rect 34057 38335 34115 38341
rect 33836 38304 33881 38332
rect 33836 38295 33848 38304
rect 34057 38301 34069 38335
rect 34103 38332 34115 38335
rect 34790 38332 34796 38344
rect 34103 38304 34796 38332
rect 34103 38301 34115 38304
rect 34057 38295 34115 38301
rect 33836 38292 33842 38295
rect 34790 38292 34796 38304
rect 34848 38332 34854 38344
rect 35529 38335 35587 38341
rect 35529 38332 35541 38335
rect 34848 38304 35541 38332
rect 34848 38292 34854 38304
rect 35529 38301 35541 38304
rect 35575 38301 35587 38335
rect 35529 38295 35587 38301
rect 38654 38292 38660 38344
rect 38712 38341 38718 38344
rect 38712 38332 38724 38341
rect 38930 38332 38936 38344
rect 38712 38304 38757 38332
rect 38891 38304 38936 38332
rect 38712 38295 38724 38304
rect 38712 38292 38718 38295
rect 38930 38292 38936 38304
rect 38988 38292 38994 38344
rect 42150 38292 42156 38344
rect 42208 38332 42214 38344
rect 42208 38304 42253 38332
rect 42208 38292 42214 38304
rect 31007 38236 31340 38264
rect 31007 38233 31019 38236
rect 30961 38227 31019 38233
rect 31662 38224 31668 38276
rect 31720 38264 31754 38276
rect 31941 38267 31999 38273
rect 31941 38264 31953 38267
rect 31720 38236 31953 38264
rect 31720 38224 31726 38236
rect 31941 38233 31953 38236
rect 31987 38264 31999 38267
rect 35796 38267 35854 38273
rect 31987 38236 32720 38264
rect 31987 38233 31999 38236
rect 31941 38227 31999 38233
rect 22738 38196 22744 38208
rect 11480 38168 22744 38196
rect 11480 38156 11486 38168
rect 22738 38156 22744 38168
rect 22796 38196 22802 38208
rect 23382 38196 23388 38208
rect 22796 38168 23388 38196
rect 22796 38156 22802 38168
rect 23382 38156 23388 38168
rect 23440 38156 23446 38208
rect 24762 38196 24768 38208
rect 24723 38168 24768 38196
rect 24762 38156 24768 38168
rect 24820 38156 24826 38208
rect 26237 38199 26295 38205
rect 26237 38165 26249 38199
rect 26283 38196 26295 38199
rect 26418 38196 26424 38208
rect 26283 38168 26424 38196
rect 26283 38165 26295 38168
rect 26237 38159 26295 38165
rect 26418 38156 26424 38168
rect 26476 38156 26482 38208
rect 30009 38199 30067 38205
rect 30009 38165 30021 38199
rect 30055 38196 30067 38199
rect 30098 38196 30104 38208
rect 30055 38168 30104 38196
rect 30055 38165 30067 38168
rect 30009 38159 30067 38165
rect 30098 38156 30104 38168
rect 30156 38156 30162 38208
rect 31202 38156 31208 38208
rect 31260 38196 31266 38208
rect 31757 38199 31815 38205
rect 31757 38196 31769 38199
rect 31260 38168 31769 38196
rect 31260 38156 31266 38168
rect 31757 38165 31769 38168
rect 31803 38165 31815 38199
rect 32122 38196 32128 38208
rect 32083 38168 32128 38196
rect 31757 38159 31815 38165
rect 32122 38156 32128 38168
rect 32180 38156 32186 38208
rect 32692 38205 32720 38236
rect 35796 38233 35808 38267
rect 35842 38264 35854 38267
rect 35986 38264 35992 38276
rect 35842 38236 35992 38264
rect 35842 38233 35854 38236
rect 35796 38227 35854 38233
rect 35986 38224 35992 38236
rect 36044 38224 36050 38276
rect 41690 38224 41696 38276
rect 41748 38264 41754 38276
rect 41969 38267 42027 38273
rect 41969 38264 41981 38267
rect 41748 38236 41981 38264
rect 41748 38224 41754 38236
rect 41969 38233 41981 38236
rect 42015 38233 42027 38267
rect 41969 38227 42027 38233
rect 32677 38199 32735 38205
rect 32677 38165 32689 38199
rect 32723 38165 32735 38199
rect 37550 38196 37556 38208
rect 37511 38168 37556 38196
rect 32677 38159 32735 38165
rect 37550 38156 37556 38168
rect 37608 38156 37614 38208
rect 1104 38106 42872 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 42872 38106
rect 1104 38032 42872 38054
rect 23937 37995 23995 38001
rect 23937 37961 23949 37995
rect 23983 37992 23995 37995
rect 24946 37992 24952 38004
rect 23983 37964 24952 37992
rect 23983 37961 23995 37964
rect 23937 37955 23995 37961
rect 24946 37952 24952 37964
rect 25004 37952 25010 38004
rect 29365 37995 29423 38001
rect 29365 37961 29377 37995
rect 29411 37992 29423 37995
rect 30282 37992 30288 38004
rect 29411 37964 30288 37992
rect 29411 37961 29423 37964
rect 29365 37955 29423 37961
rect 30282 37952 30288 37964
rect 30340 37952 30346 38004
rect 31202 37992 31208 38004
rect 31163 37964 31208 37992
rect 31202 37952 31208 37964
rect 31260 37952 31266 38004
rect 32677 37995 32735 38001
rect 32677 37961 32689 37995
rect 32723 37992 32735 37995
rect 33502 37992 33508 38004
rect 32723 37964 33508 37992
rect 32723 37961 32735 37964
rect 32677 37955 32735 37961
rect 33502 37952 33508 37964
rect 33560 37952 33566 38004
rect 36078 37952 36084 38004
rect 36136 37992 36142 38004
rect 36265 37995 36323 38001
rect 36265 37992 36277 37995
rect 36136 37964 36277 37992
rect 36136 37952 36142 37964
rect 36265 37961 36277 37964
rect 36311 37961 36323 37995
rect 38102 37992 38108 38004
rect 38063 37964 38108 37992
rect 36265 37955 36323 37961
rect 38102 37952 38108 37964
rect 38160 37952 38166 38004
rect 38838 37952 38844 38004
rect 38896 37992 38902 38004
rect 38933 37995 38991 38001
rect 38933 37992 38945 37995
rect 38896 37964 38945 37992
rect 38896 37952 38902 37964
rect 38933 37961 38945 37964
rect 38979 37961 38991 37995
rect 38933 37955 38991 37961
rect 39114 37952 39120 38004
rect 39172 37992 39178 38004
rect 41141 37995 41199 38001
rect 41141 37992 41153 37995
rect 39172 37964 41153 37992
rect 39172 37952 39178 37964
rect 41141 37961 41153 37964
rect 41187 37961 41199 37995
rect 41690 37992 41696 38004
rect 41651 37964 41696 37992
rect 41141 37955 41199 37961
rect 41690 37952 41696 37964
rect 41748 37952 41754 38004
rect 4246 37924 4252 37936
rect 4207 37896 4252 37924
rect 4246 37884 4252 37896
rect 4304 37884 4310 37936
rect 11974 37924 11980 37936
rect 11935 37896 11980 37924
rect 11974 37884 11980 37896
rect 12032 37884 12038 37936
rect 26326 37924 26332 37936
rect 21836 37896 26332 37924
rect 21836 37868 21864 37896
rect 4430 37816 4436 37868
rect 4488 37856 4494 37868
rect 4488 37828 4533 37856
rect 4488 37816 4494 37828
rect 10870 37816 10876 37868
rect 10928 37856 10934 37868
rect 17494 37865 17500 37868
rect 11609 37859 11667 37865
rect 11609 37856 11621 37859
rect 10928 37828 11621 37856
rect 10928 37816 10934 37828
rect 11609 37825 11621 37828
rect 11655 37825 11667 37859
rect 11609 37819 11667 37825
rect 17488 37819 17500 37865
rect 17552 37856 17558 37868
rect 21818 37856 21824 37868
rect 17552 37828 17588 37856
rect 21731 37828 21824 37856
rect 17494 37816 17500 37819
rect 17552 37816 17558 37828
rect 21818 37816 21824 37828
rect 21876 37816 21882 37868
rect 21910 37816 21916 37868
rect 21968 37856 21974 37868
rect 22077 37859 22135 37865
rect 22077 37856 22089 37859
rect 21968 37828 22089 37856
rect 21968 37816 21974 37828
rect 22077 37825 22089 37828
rect 22123 37825 22135 37859
rect 23842 37856 23848 37868
rect 23803 37828 23848 37856
rect 22077 37819 22135 37825
rect 23842 37816 23848 37828
rect 23900 37816 23906 37868
rect 24118 37856 24124 37868
rect 24079 37828 24124 37856
rect 24118 37816 24124 37828
rect 24176 37816 24182 37868
rect 25056 37865 25084 37896
rect 26326 37884 26332 37896
rect 26384 37884 26390 37936
rect 28442 37924 28448 37936
rect 28000 37896 28448 37924
rect 25041 37859 25099 37865
rect 25041 37825 25053 37859
rect 25087 37825 25099 37859
rect 25041 37819 25099 37825
rect 25130 37816 25136 37868
rect 25188 37856 25194 37868
rect 28000 37865 28028 37896
rect 28442 37884 28448 37896
rect 28500 37924 28506 37936
rect 32493 37927 32551 37933
rect 28500 37896 29868 37924
rect 28500 37884 28506 37896
rect 28258 37865 28264 37868
rect 25297 37859 25355 37865
rect 25297 37856 25309 37859
rect 25188 37828 25309 37856
rect 25188 37816 25194 37828
rect 25297 37825 25309 37828
rect 25343 37825 25355 37859
rect 25297 37819 25355 37825
rect 27985 37859 28043 37865
rect 27985 37825 27997 37859
rect 28031 37825 28043 37859
rect 27985 37819 28043 37825
rect 28252 37819 28264 37865
rect 28316 37856 28322 37868
rect 29840 37865 29868 37896
rect 32493 37893 32505 37927
rect 32539 37924 32551 37927
rect 32766 37924 32772 37936
rect 32539 37896 32772 37924
rect 32539 37893 32551 37896
rect 32493 37887 32551 37893
rect 32766 37884 32772 37896
rect 32824 37884 32830 37936
rect 33796 37896 41414 37924
rect 30098 37865 30104 37868
rect 29825 37859 29883 37865
rect 28316 37828 28352 37856
rect 28258 37816 28264 37819
rect 28316 37816 28322 37828
rect 29825 37825 29837 37859
rect 29871 37825 29883 37859
rect 30092 37856 30104 37865
rect 30059 37828 30104 37856
rect 29825 37819 29883 37825
rect 30092 37819 30104 37828
rect 30098 37816 30104 37819
rect 30156 37816 30162 37868
rect 32125 37859 32183 37865
rect 32125 37825 32137 37859
rect 32171 37856 32183 37859
rect 32674 37856 32680 37868
rect 32171 37828 32680 37856
rect 32171 37825 32183 37828
rect 32125 37819 32183 37825
rect 32674 37816 32680 37828
rect 32732 37816 32738 37868
rect 2774 37788 2780 37800
rect 2735 37760 2780 37788
rect 2774 37748 2780 37760
rect 2832 37748 2838 37800
rect 16574 37748 16580 37800
rect 16632 37788 16638 37800
rect 17221 37791 17279 37797
rect 17221 37788 17233 37791
rect 16632 37760 17233 37788
rect 16632 37748 16638 37760
rect 17221 37757 17233 37760
rect 17267 37757 17279 37791
rect 17221 37751 17279 37757
rect 33796 37720 33824 37896
rect 34514 37856 34520 37868
rect 34572 37865 34578 37868
rect 34484 37828 34520 37856
rect 34514 37816 34520 37828
rect 34572 37819 34584 37865
rect 36541 37859 36599 37865
rect 36541 37825 36553 37859
rect 36587 37856 36599 37859
rect 36906 37856 36912 37868
rect 36587 37828 36912 37856
rect 36587 37825 36599 37828
rect 36541 37819 36599 37825
rect 34572 37816 34578 37819
rect 36906 37816 36912 37828
rect 36964 37816 36970 37868
rect 37550 37816 37556 37868
rect 37608 37856 37614 37868
rect 38381 37859 38439 37865
rect 38381 37856 38393 37859
rect 37608 37828 38393 37856
rect 37608 37816 37614 37828
rect 38381 37825 38393 37828
rect 38427 37825 38439 37859
rect 38381 37819 38439 37825
rect 38654 37816 38660 37868
rect 38712 37856 38718 37868
rect 38841 37859 38899 37865
rect 38841 37856 38853 37859
rect 38712 37828 38853 37856
rect 38712 37816 38718 37828
rect 38841 37825 38853 37828
rect 38887 37825 38899 37859
rect 39114 37856 39120 37868
rect 39075 37828 39120 37856
rect 38841 37819 38899 37825
rect 39114 37816 39120 37828
rect 39172 37816 39178 37868
rect 40034 37865 40040 37868
rect 40028 37819 40040 37865
rect 40092 37856 40098 37868
rect 41386 37856 41414 37896
rect 41601 37859 41659 37865
rect 41601 37856 41613 37859
rect 40092 37828 40128 37856
rect 41386 37828 41613 37856
rect 40034 37816 40040 37819
rect 40092 37816 40098 37828
rect 41601 37825 41613 37828
rect 41647 37856 41659 37859
rect 42334 37856 42340 37868
rect 41647 37828 42340 37856
rect 41647 37825 41659 37828
rect 41601 37819 41659 37825
rect 42334 37816 42340 37828
rect 42392 37816 42398 37868
rect 34790 37788 34796 37800
rect 34751 37760 34796 37788
rect 34790 37748 34796 37760
rect 34848 37748 34854 37800
rect 36265 37791 36323 37797
rect 36265 37757 36277 37791
rect 36311 37757 36323 37791
rect 36446 37788 36452 37800
rect 36407 37760 36452 37788
rect 36265 37751 36323 37757
rect 30760 37692 33824 37720
rect 36280 37720 36308 37751
rect 36446 37748 36452 37760
rect 36504 37748 36510 37800
rect 38102 37788 38108 37800
rect 38063 37760 38108 37788
rect 38102 37748 38108 37760
rect 38160 37748 38166 37800
rect 39761 37791 39819 37797
rect 39761 37788 39773 37791
rect 38948 37760 39773 37788
rect 38948 37732 38976 37760
rect 39761 37757 39773 37760
rect 39807 37757 39819 37791
rect 39761 37751 39819 37757
rect 36354 37720 36360 37732
rect 36280 37692 36360 37720
rect 1670 37652 1676 37664
rect 1631 37624 1676 37652
rect 1670 37612 1676 37624
rect 1728 37612 1734 37664
rect 17862 37612 17868 37664
rect 17920 37652 17926 37664
rect 18322 37652 18328 37664
rect 17920 37624 18328 37652
rect 17920 37612 17926 37624
rect 18322 37612 18328 37624
rect 18380 37652 18386 37664
rect 18601 37655 18659 37661
rect 18601 37652 18613 37655
rect 18380 37624 18613 37652
rect 18380 37612 18386 37624
rect 18601 37621 18613 37624
rect 18647 37621 18659 37655
rect 18601 37615 18659 37621
rect 23201 37655 23259 37661
rect 23201 37621 23213 37655
rect 23247 37652 23259 37655
rect 23290 37652 23296 37664
rect 23247 37624 23296 37652
rect 23247 37621 23259 37624
rect 23201 37615 23259 37621
rect 23290 37612 23296 37624
rect 23348 37612 23354 37664
rect 24302 37652 24308 37664
rect 24263 37624 24308 37652
rect 24302 37612 24308 37624
rect 24360 37612 24366 37664
rect 25958 37612 25964 37664
rect 26016 37652 26022 37664
rect 26421 37655 26479 37661
rect 26421 37652 26433 37655
rect 26016 37624 26433 37652
rect 26016 37612 26022 37624
rect 26421 37621 26433 37624
rect 26467 37621 26479 37655
rect 26421 37615 26479 37621
rect 26602 37612 26608 37664
rect 26660 37652 26666 37664
rect 30760 37652 30788 37692
rect 36354 37680 36360 37692
rect 36412 37720 36418 37732
rect 36412 37692 38884 37720
rect 36412 37680 36418 37692
rect 26660 37624 30788 37652
rect 26660 37612 26666 37624
rect 31294 37612 31300 37664
rect 31352 37652 31358 37664
rect 32493 37655 32551 37661
rect 32493 37652 32505 37655
rect 31352 37624 32505 37652
rect 31352 37612 31358 37624
rect 32493 37621 32505 37624
rect 32539 37621 32551 37655
rect 32493 37615 32551 37621
rect 32858 37612 32864 37664
rect 32916 37652 32922 37664
rect 33413 37655 33471 37661
rect 33413 37652 33425 37655
rect 32916 37624 33425 37652
rect 32916 37612 32922 37624
rect 33413 37621 33425 37624
rect 33459 37621 33471 37655
rect 33413 37615 33471 37621
rect 38289 37655 38347 37661
rect 38289 37621 38301 37655
rect 38335 37652 38347 37655
rect 38746 37652 38752 37664
rect 38335 37624 38752 37652
rect 38335 37621 38347 37624
rect 38289 37615 38347 37621
rect 38746 37612 38752 37624
rect 38804 37612 38810 37664
rect 38856 37652 38884 37692
rect 38930 37680 38936 37732
rect 38988 37680 38994 37732
rect 39022 37652 39028 37664
rect 38856 37624 39028 37652
rect 39022 37612 39028 37624
rect 39080 37612 39086 37664
rect 39114 37612 39120 37664
rect 39172 37652 39178 37664
rect 39301 37655 39359 37661
rect 39301 37652 39313 37655
rect 39172 37624 39313 37652
rect 39172 37612 39178 37624
rect 39301 37621 39313 37624
rect 39347 37621 39359 37655
rect 39301 37615 39359 37621
rect 1104 37562 42872 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 42872 37562
rect 1104 37488 42872 37510
rect 17405 37451 17463 37457
rect 17405 37417 17417 37451
rect 17451 37448 17463 37451
rect 17494 37448 17500 37460
rect 17451 37420 17500 37448
rect 17451 37417 17463 37420
rect 17405 37411 17463 37417
rect 17494 37408 17500 37420
rect 17552 37408 17558 37460
rect 20806 37408 20812 37460
rect 20864 37448 20870 37460
rect 22925 37451 22983 37457
rect 22925 37448 22937 37451
rect 20864 37420 22937 37448
rect 20864 37408 20870 37420
rect 22925 37417 22937 37420
rect 22971 37417 22983 37451
rect 25130 37448 25136 37460
rect 25091 37420 25136 37448
rect 22925 37411 22983 37417
rect 25130 37408 25136 37420
rect 25188 37408 25194 37460
rect 28813 37451 28871 37457
rect 28813 37417 28825 37451
rect 28859 37448 28871 37451
rect 29730 37448 29736 37460
rect 28859 37420 29736 37448
rect 28859 37417 28871 37420
rect 28813 37411 28871 37417
rect 29730 37408 29736 37420
rect 29788 37408 29794 37460
rect 30101 37451 30159 37457
rect 30101 37417 30113 37451
rect 30147 37448 30159 37451
rect 30190 37448 30196 37460
rect 30147 37420 30196 37448
rect 30147 37417 30159 37420
rect 30101 37411 30159 37417
rect 30190 37408 30196 37420
rect 30248 37408 30254 37460
rect 31113 37451 31171 37457
rect 31113 37417 31125 37451
rect 31159 37448 31171 37451
rect 31294 37448 31300 37460
rect 31159 37420 31300 37448
rect 31159 37417 31171 37420
rect 31113 37411 31171 37417
rect 31294 37408 31300 37420
rect 31352 37408 31358 37460
rect 31662 37448 31668 37460
rect 31623 37420 31668 37448
rect 31662 37408 31668 37420
rect 31720 37408 31726 37460
rect 33318 37448 33324 37460
rect 33279 37420 33324 37448
rect 33318 37408 33324 37420
rect 33376 37408 33382 37460
rect 39117 37451 39175 37457
rect 39117 37448 39129 37451
rect 33888 37420 39129 37448
rect 29914 37380 29920 37392
rect 29875 37352 29920 37380
rect 29914 37340 29920 37352
rect 29972 37340 29978 37392
rect 1397 37315 1455 37321
rect 1397 37281 1409 37315
rect 1443 37312 1455 37315
rect 1670 37312 1676 37324
rect 1443 37284 1676 37312
rect 1443 37281 1455 37284
rect 1397 37275 1455 37281
rect 1670 37272 1676 37284
rect 1728 37272 1734 37324
rect 17681 37315 17739 37321
rect 17681 37281 17693 37315
rect 17727 37312 17739 37315
rect 17862 37312 17868 37324
rect 17727 37284 17868 37312
rect 17727 37281 17739 37284
rect 17681 37275 17739 37281
rect 17862 37272 17868 37284
rect 17920 37272 17926 37324
rect 23109 37315 23167 37321
rect 23109 37281 23121 37315
rect 23155 37312 23167 37315
rect 24302 37312 24308 37324
rect 23155 37284 24308 37312
rect 23155 37281 23167 37284
rect 23109 37275 23167 37281
rect 24302 37272 24308 37284
rect 24360 37272 24366 37324
rect 33888 37312 33916 37420
rect 39117 37417 39129 37420
rect 39163 37448 39175 37451
rect 39298 37448 39304 37460
rect 39163 37420 39304 37448
rect 39163 37417 39175 37420
rect 39117 37411 39175 37417
rect 39298 37408 39304 37420
rect 39356 37408 39362 37460
rect 40034 37448 40040 37460
rect 39995 37420 40040 37448
rect 40034 37408 40040 37420
rect 40092 37408 40098 37460
rect 41785 37451 41843 37457
rect 41785 37417 41797 37451
rect 41831 37448 41843 37451
rect 42150 37448 42156 37460
rect 41831 37420 42156 37448
rect 41831 37417 41843 37420
rect 41785 37411 41843 37417
rect 42150 37408 42156 37420
rect 42208 37408 42214 37460
rect 38746 37380 38752 37392
rect 38707 37352 38752 37380
rect 38746 37340 38752 37352
rect 38804 37340 38810 37392
rect 37550 37312 37556 37324
rect 33428 37284 33916 37312
rect 37511 37284 37556 37312
rect 2958 37204 2964 37256
rect 3016 37244 3022 37256
rect 3237 37247 3295 37253
rect 3237 37244 3249 37247
rect 3016 37216 3249 37244
rect 3016 37204 3022 37216
rect 3237 37213 3249 37216
rect 3283 37213 3295 37247
rect 3237 37207 3295 37213
rect 4614 37204 4620 37256
rect 4672 37244 4678 37256
rect 4985 37247 5043 37253
rect 4985 37244 4997 37247
rect 4672 37216 4997 37244
rect 4672 37204 4678 37216
rect 4985 37213 4997 37216
rect 5031 37213 5043 37247
rect 4985 37207 5043 37213
rect 14090 37204 14096 37256
rect 14148 37244 14154 37256
rect 15473 37247 15531 37253
rect 15473 37244 15485 37247
rect 14148 37216 15485 37244
rect 14148 37204 14154 37216
rect 15473 37213 15485 37216
rect 15519 37244 15531 37247
rect 16574 37244 16580 37256
rect 15519 37216 16580 37244
rect 15519 37213 15531 37216
rect 15473 37207 15531 37213
rect 16574 37204 16580 37216
rect 16632 37204 16638 37256
rect 17218 37204 17224 37256
rect 17276 37244 17282 37256
rect 17589 37247 17647 37253
rect 17589 37244 17601 37247
rect 17276 37216 17601 37244
rect 17276 37204 17282 37216
rect 17589 37213 17601 37216
rect 17635 37213 17647 37247
rect 17589 37207 17647 37213
rect 18509 37247 18567 37253
rect 18509 37213 18521 37247
rect 18555 37244 18567 37247
rect 18598 37244 18604 37256
rect 18555 37216 18604 37244
rect 18555 37213 18567 37216
rect 18509 37207 18567 37213
rect 18598 37204 18604 37216
rect 18656 37204 18662 37256
rect 20625 37247 20683 37253
rect 20625 37213 20637 37247
rect 20671 37244 20683 37247
rect 20714 37244 20720 37256
rect 20671 37216 20720 37244
rect 20671 37213 20683 37216
rect 20625 37207 20683 37213
rect 20714 37204 20720 37216
rect 20772 37244 20778 37256
rect 21085 37247 21143 37253
rect 21085 37244 21097 37247
rect 20772 37216 21097 37244
rect 20772 37204 20778 37216
rect 21085 37213 21097 37216
rect 21131 37213 21143 37247
rect 23198 37244 23204 37256
rect 23159 37216 23204 37244
rect 21085 37207 21143 37213
rect 23198 37204 23204 37216
rect 23256 37204 23262 37256
rect 23290 37204 23296 37256
rect 23348 37244 23354 37256
rect 24397 37247 24455 37253
rect 24397 37244 24409 37247
rect 23348 37216 24409 37244
rect 23348 37204 23354 37216
rect 24397 37213 24409 37216
rect 24443 37213 24455 37247
rect 25314 37244 25320 37256
rect 25275 37216 25320 37244
rect 24397 37207 24455 37213
rect 25314 37204 25320 37216
rect 25372 37204 25378 37256
rect 25409 37247 25467 37253
rect 25409 37213 25421 37247
rect 25455 37244 25467 37247
rect 25958 37244 25964 37256
rect 25455 37216 25964 37244
rect 25455 37213 25467 37216
rect 25409 37207 25467 37213
rect 25958 37204 25964 37216
rect 26016 37204 26022 37256
rect 26326 37244 26332 37256
rect 26287 37216 26332 37244
rect 26326 37204 26332 37216
rect 26384 37204 26390 37256
rect 29641 37247 29699 37253
rect 29641 37213 29653 37247
rect 29687 37244 29699 37247
rect 30650 37244 30656 37256
rect 29687 37216 30656 37244
rect 29687 37213 29699 37216
rect 29641 37207 29699 37213
rect 30650 37204 30656 37216
rect 30708 37204 30714 37256
rect 30929 37247 30987 37253
rect 30929 37213 30941 37247
rect 30975 37244 30987 37247
rect 31662 37244 31668 37256
rect 30975 37216 31668 37244
rect 30975 37213 30987 37216
rect 30929 37207 30987 37213
rect 31662 37204 31668 37216
rect 31720 37204 31726 37256
rect 31849 37247 31907 37253
rect 31849 37213 31861 37247
rect 31895 37213 31907 37247
rect 31849 37207 31907 37213
rect 32033 37247 32091 37253
rect 32033 37213 32045 37247
rect 32079 37244 32091 37247
rect 32858 37244 32864 37256
rect 32079 37216 32864 37244
rect 32079 37213 32091 37216
rect 32033 37207 32091 37213
rect 1581 37179 1639 37185
rect 1581 37145 1593 37179
rect 1627 37176 1639 37179
rect 2038 37176 2044 37188
rect 1627 37148 2044 37176
rect 1627 37145 1639 37148
rect 1581 37139 1639 37145
rect 2038 37136 2044 37148
rect 2096 37136 2102 37188
rect 4341 37179 4399 37185
rect 4341 37145 4353 37179
rect 4387 37176 4399 37179
rect 4890 37176 4896 37188
rect 4387 37148 4896 37176
rect 4387 37145 4399 37148
rect 4341 37139 4399 37145
rect 4890 37136 4896 37148
rect 4948 37136 4954 37188
rect 15562 37136 15568 37188
rect 15620 37176 15626 37188
rect 15718 37179 15776 37185
rect 15718 37176 15730 37179
rect 15620 37148 15730 37176
rect 15620 37136 15626 37148
rect 15718 37145 15730 37148
rect 15764 37145 15776 37179
rect 20358 37179 20416 37185
rect 20358 37176 20370 37179
rect 15718 37139 15776 37145
rect 18708 37148 20370 37176
rect 16850 37108 16856 37120
rect 16811 37080 16856 37108
rect 16850 37068 16856 37080
rect 16908 37068 16914 37120
rect 18046 37108 18052 37120
rect 18007 37080 18052 37108
rect 18046 37068 18052 37080
rect 18104 37068 18110 37120
rect 18708 37117 18736 37148
rect 20358 37145 20370 37148
rect 20404 37145 20416 37179
rect 20358 37139 20416 37145
rect 20530 37136 20536 37188
rect 20588 37176 20594 37188
rect 21330 37179 21388 37185
rect 21330 37176 21342 37179
rect 20588 37148 21342 37176
rect 20588 37136 20594 37148
rect 21330 37145 21342 37148
rect 21376 37145 21388 37179
rect 21330 37139 21388 37145
rect 24489 37179 24547 37185
rect 24489 37145 24501 37179
rect 24535 37176 24547 37179
rect 25130 37176 25136 37188
rect 24535 37148 25136 37176
rect 24535 37145 24547 37148
rect 24489 37139 24547 37145
rect 25130 37136 25136 37148
rect 25188 37136 25194 37188
rect 25866 37136 25872 37188
rect 25924 37176 25930 37188
rect 26602 37185 26608 37188
rect 25924 37148 26556 37176
rect 25924 37136 25930 37148
rect 18693 37111 18751 37117
rect 18693 37077 18705 37111
rect 18739 37077 18751 37111
rect 19242 37108 19248 37120
rect 19203 37080 19248 37108
rect 18693 37071 18751 37077
rect 19242 37068 19248 37080
rect 19300 37068 19306 37120
rect 22462 37108 22468 37120
rect 22423 37080 22468 37108
rect 22462 37068 22468 37080
rect 22520 37068 22526 37120
rect 23198 37068 23204 37120
rect 23256 37108 23262 37120
rect 23569 37111 23627 37117
rect 23569 37108 23581 37111
rect 23256 37080 23581 37108
rect 23256 37068 23262 37080
rect 23569 37077 23581 37080
rect 23615 37077 23627 37111
rect 23569 37071 23627 37077
rect 24854 37068 24860 37120
rect 24912 37108 24918 37120
rect 25777 37111 25835 37117
rect 25777 37108 25789 37111
rect 24912 37080 25789 37108
rect 24912 37068 24918 37080
rect 25777 37077 25789 37080
rect 25823 37108 25835 37111
rect 26050 37108 26056 37120
rect 25823 37080 26056 37108
rect 25823 37077 25835 37080
rect 25777 37071 25835 37077
rect 26050 37068 26056 37080
rect 26108 37068 26114 37120
rect 26528 37108 26556 37148
rect 26596 37139 26608 37185
rect 26660 37176 26666 37188
rect 28994 37176 29000 37188
rect 26660 37148 26696 37176
rect 28955 37148 29000 37176
rect 26602 37136 26608 37139
rect 26660 37136 26666 37148
rect 28994 37136 29000 37148
rect 29052 37136 29058 37188
rect 29730 37136 29736 37188
rect 29788 37176 29794 37188
rect 31573 37179 31631 37185
rect 29788 37148 30880 37176
rect 29788 37136 29794 37148
rect 27709 37111 27767 37117
rect 27709 37108 27721 37111
rect 26528 37080 27721 37108
rect 27709 37077 27721 37080
rect 27755 37077 27767 37111
rect 28626 37108 28632 37120
rect 28587 37080 28632 37108
rect 27709 37071 27767 37077
rect 28626 37068 28632 37080
rect 28684 37068 28690 37120
rect 28797 37111 28855 37117
rect 28797 37077 28809 37111
rect 28843 37108 28855 37111
rect 28902 37108 28908 37120
rect 28843 37080 28908 37108
rect 28843 37077 28855 37080
rect 28797 37071 28855 37077
rect 28902 37068 28908 37080
rect 28960 37068 28966 37120
rect 30282 37068 30288 37120
rect 30340 37108 30346 37120
rect 30745 37111 30803 37117
rect 30745 37108 30757 37111
rect 30340 37080 30757 37108
rect 30340 37068 30346 37080
rect 30745 37077 30757 37080
rect 30791 37077 30803 37111
rect 30852 37108 30880 37148
rect 31573 37145 31585 37179
rect 31619 37176 31631 37179
rect 31754 37176 31760 37188
rect 31619 37148 31760 37176
rect 31619 37145 31631 37148
rect 31573 37139 31631 37145
rect 31754 37136 31760 37148
rect 31812 37136 31818 37188
rect 31864 37108 31892 37207
rect 32858 37204 32864 37216
rect 32916 37204 32922 37256
rect 32950 37204 32956 37256
rect 33008 37244 33014 37256
rect 33008 37216 33053 37244
rect 33008 37204 33014 37216
rect 33321 37179 33379 37185
rect 33321 37145 33333 37179
rect 33367 37176 33379 37179
rect 33428 37176 33456 37284
rect 37550 37272 37556 37284
rect 37608 37272 37614 37324
rect 33965 37247 34023 37253
rect 33965 37244 33977 37247
rect 33367 37148 33456 37176
rect 33520 37216 33977 37244
rect 33367 37145 33379 37148
rect 33321 37139 33379 37145
rect 32214 37108 32220 37120
rect 30852 37080 31892 37108
rect 32175 37080 32220 37108
rect 30745 37071 30803 37077
rect 32214 37068 32220 37080
rect 32272 37068 32278 37120
rect 32858 37068 32864 37120
rect 32916 37108 32922 37120
rect 33336 37108 33364 37139
rect 33520 37117 33548 37216
rect 33965 37213 33977 37216
rect 34011 37213 34023 37247
rect 33965 37207 34023 37213
rect 36081 37247 36139 37253
rect 36081 37213 36093 37247
rect 36127 37213 36139 37247
rect 36081 37207 36139 37213
rect 36357 37247 36415 37253
rect 36357 37213 36369 37247
rect 36403 37244 36415 37247
rect 36446 37244 36452 37256
rect 36403 37216 36452 37244
rect 36403 37213 36415 37216
rect 36357 37207 36415 37213
rect 36096 37176 36124 37207
rect 36446 37204 36452 37216
rect 36504 37204 36510 37256
rect 37185 37247 37243 37253
rect 37185 37213 37197 37247
rect 37231 37213 37243 37247
rect 37185 37207 37243 37213
rect 37670 37247 37728 37253
rect 37670 37213 37682 37247
rect 37716 37244 37728 37247
rect 39206 37244 39212 37256
rect 37716 37216 39212 37244
rect 37716 37213 37728 37216
rect 37670 37207 37728 37213
rect 36538 37176 36544 37188
rect 36096 37148 36544 37176
rect 36538 37136 36544 37148
rect 36596 37176 36602 37188
rect 37200 37176 37228 37207
rect 39206 37204 39212 37216
rect 39264 37204 39270 37256
rect 39853 37247 39911 37253
rect 39853 37244 39865 37247
rect 39316 37216 39865 37244
rect 39114 37176 39120 37188
rect 36596 37148 37228 37176
rect 39075 37148 39120 37176
rect 36596 37136 36602 37148
rect 39114 37136 39120 37148
rect 39172 37136 39178 37188
rect 32916 37080 33364 37108
rect 33505 37111 33563 37117
rect 32916 37068 32922 37080
rect 33505 37077 33517 37111
rect 33551 37077 33563 37111
rect 33505 37071 33563 37077
rect 34149 37111 34207 37117
rect 34149 37077 34161 37111
rect 34195 37108 34207 37111
rect 34514 37108 34520 37120
rect 34195 37080 34520 37108
rect 34195 37077 34207 37080
rect 34149 37071 34207 37077
rect 34514 37068 34520 37080
rect 34572 37068 34578 37120
rect 35894 37108 35900 37120
rect 35855 37080 35900 37108
rect 35894 37068 35900 37080
rect 35952 37068 35958 37120
rect 36265 37111 36323 37117
rect 36265 37077 36277 37111
rect 36311 37108 36323 37111
rect 36630 37108 36636 37120
rect 36311 37080 36636 37108
rect 36311 37077 36323 37080
rect 36265 37071 36323 37077
rect 36630 37068 36636 37080
rect 36688 37108 36694 37120
rect 36906 37108 36912 37120
rect 36688 37080 36912 37108
rect 36688 37068 36694 37080
rect 36906 37068 36912 37080
rect 36964 37108 36970 37120
rect 37461 37111 37519 37117
rect 37461 37108 37473 37111
rect 36964 37080 37473 37108
rect 36964 37068 36970 37080
rect 37461 37077 37473 37080
rect 37507 37077 37519 37111
rect 37826 37108 37832 37120
rect 37787 37080 37832 37108
rect 37461 37071 37519 37077
rect 37826 37068 37832 37080
rect 37884 37068 37890 37120
rect 39316 37117 39344 37216
rect 39853 37213 39865 37216
rect 39899 37213 39911 37247
rect 39853 37207 39911 37213
rect 39301 37111 39359 37117
rect 39301 37077 39313 37111
rect 39347 37077 39359 37111
rect 39301 37071 39359 37077
rect 1104 37018 42872 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 42872 37018
rect 1104 36944 42872 36966
rect 2038 36904 2044 36916
rect 1999 36876 2044 36904
rect 2038 36864 2044 36876
rect 2096 36864 2102 36916
rect 15562 36904 15568 36916
rect 15523 36876 15568 36904
rect 15562 36864 15568 36876
rect 15620 36864 15626 36916
rect 18598 36904 18604 36916
rect 18559 36876 18604 36904
rect 18598 36864 18604 36876
rect 18656 36864 18662 36916
rect 20349 36907 20407 36913
rect 20349 36873 20361 36907
rect 20395 36904 20407 36907
rect 20530 36904 20536 36916
rect 20395 36876 20536 36904
rect 20395 36873 20407 36876
rect 20349 36867 20407 36873
rect 20530 36864 20536 36876
rect 20588 36864 20594 36916
rect 21082 36904 21088 36916
rect 20640 36876 21088 36904
rect 2222 36836 2228 36848
rect 2135 36808 2228 36836
rect 2148 36777 2176 36808
rect 2222 36796 2228 36808
rect 2280 36836 2286 36848
rect 4890 36836 4896 36848
rect 2280 36808 4896 36836
rect 2280 36796 2286 36808
rect 4890 36796 4896 36808
rect 4948 36796 4954 36848
rect 14550 36796 14556 36848
rect 14608 36836 14614 36848
rect 20640 36836 20668 36876
rect 21082 36864 21088 36876
rect 21140 36864 21146 36916
rect 23198 36904 23204 36916
rect 23159 36876 23204 36904
rect 23198 36864 23204 36876
rect 23256 36864 23262 36916
rect 25222 36904 25228 36916
rect 23584 36876 25228 36904
rect 14608 36808 20668 36836
rect 14608 36796 14614 36808
rect 22462 36796 22468 36848
rect 22520 36836 22526 36848
rect 23584 36836 23612 36876
rect 25222 36864 25228 36876
rect 25280 36864 25286 36916
rect 25314 36864 25320 36916
rect 25372 36904 25378 36916
rect 25777 36907 25835 36913
rect 25777 36904 25789 36907
rect 25372 36876 25789 36904
rect 25372 36864 25378 36876
rect 25777 36873 25789 36876
rect 25823 36873 25835 36907
rect 28258 36904 28264 36916
rect 28219 36876 28264 36904
rect 25777 36867 25835 36873
rect 28258 36864 28264 36876
rect 28316 36864 28322 36916
rect 28902 36904 28908 36916
rect 28863 36876 28908 36904
rect 28902 36864 28908 36876
rect 28960 36864 28966 36916
rect 29549 36907 29607 36913
rect 29549 36873 29561 36907
rect 29595 36904 29607 36907
rect 29730 36904 29736 36916
rect 29595 36876 29736 36904
rect 29595 36873 29607 36876
rect 29549 36867 29607 36873
rect 29730 36864 29736 36876
rect 29788 36864 29794 36916
rect 30650 36904 30656 36916
rect 29932 36876 30656 36904
rect 22520 36808 23612 36836
rect 23661 36839 23719 36845
rect 22520 36796 22526 36808
rect 23661 36805 23673 36839
rect 23707 36836 23719 36839
rect 23842 36836 23848 36848
rect 23707 36808 23848 36836
rect 23707 36805 23719 36808
rect 23661 36799 23719 36805
rect 23842 36796 23848 36808
rect 23900 36836 23906 36848
rect 29932 36845 29960 36876
rect 30650 36864 30656 36876
rect 30708 36904 30714 36916
rect 31297 36907 31355 36913
rect 31297 36904 31309 36907
rect 30708 36876 31309 36904
rect 30708 36864 30714 36876
rect 31297 36873 31309 36876
rect 31343 36873 31355 36907
rect 36538 36904 36544 36916
rect 36499 36876 36544 36904
rect 31297 36867 31355 36873
rect 36538 36864 36544 36876
rect 36596 36864 36602 36916
rect 37550 36864 37556 36916
rect 37608 36904 37614 36916
rect 38565 36907 38623 36913
rect 38565 36904 38577 36907
rect 37608 36876 38577 36904
rect 37608 36864 37614 36876
rect 38565 36873 38577 36876
rect 38611 36873 38623 36907
rect 38565 36867 38623 36873
rect 38746 36864 38752 36916
rect 38804 36904 38810 36916
rect 39209 36907 39267 36913
rect 39209 36904 39221 36907
rect 38804 36876 39221 36904
rect 38804 36864 38810 36876
rect 39209 36873 39221 36876
rect 39255 36873 39267 36907
rect 39209 36867 39267 36873
rect 29917 36839 29975 36845
rect 29917 36836 29929 36839
rect 23900 36808 25452 36836
rect 23900 36796 23906 36808
rect 2133 36771 2191 36777
rect 2133 36737 2145 36771
rect 2179 36737 2191 36771
rect 2133 36731 2191 36737
rect 3513 36771 3571 36777
rect 3513 36737 3525 36771
rect 3559 36768 3571 36771
rect 4249 36771 4307 36777
rect 4249 36768 4261 36771
rect 3559 36740 4261 36768
rect 3559 36737 3571 36740
rect 3513 36731 3571 36737
rect 4249 36737 4261 36740
rect 4295 36768 4307 36771
rect 4614 36768 4620 36780
rect 4295 36740 4620 36768
rect 4295 36737 4307 36740
rect 4249 36731 4307 36737
rect 4614 36728 4620 36740
rect 4672 36728 4678 36780
rect 5534 36728 5540 36780
rect 5592 36768 5598 36780
rect 5810 36768 5816 36780
rect 5592 36740 5816 36768
rect 5592 36728 5598 36740
rect 5810 36728 5816 36740
rect 5868 36768 5874 36780
rect 10226 36768 10232 36780
rect 5868 36740 10232 36768
rect 5868 36728 5874 36740
rect 10226 36728 10232 36740
rect 10284 36728 10290 36780
rect 14185 36771 14243 36777
rect 14185 36737 14197 36771
rect 14231 36737 14243 36771
rect 14185 36731 14243 36737
rect 3237 36703 3295 36709
rect 3237 36669 3249 36703
rect 3283 36700 3295 36703
rect 4522 36700 4528 36712
rect 3283 36672 4528 36700
rect 3283 36669 3295 36672
rect 3237 36663 3295 36669
rect 4522 36660 4528 36672
rect 4580 36660 4586 36712
rect 4893 36703 4951 36709
rect 4893 36669 4905 36703
rect 4939 36700 4951 36703
rect 4982 36700 4988 36712
rect 4939 36672 4988 36700
rect 4939 36669 4951 36672
rect 4893 36663 4951 36669
rect 4982 36660 4988 36672
rect 5040 36660 5046 36712
rect 14200 36700 14228 36731
rect 14274 36728 14280 36780
rect 14332 36768 14338 36780
rect 14461 36771 14519 36777
rect 14332 36740 14377 36768
rect 14332 36728 14338 36740
rect 14461 36737 14473 36771
rect 14507 36768 14519 36771
rect 15654 36768 15660 36780
rect 14507 36740 15660 36768
rect 14507 36737 14519 36740
rect 14461 36731 14519 36737
rect 15654 36728 15660 36740
rect 15712 36728 15718 36780
rect 15841 36771 15899 36777
rect 15841 36737 15853 36771
rect 15887 36768 15899 36771
rect 15930 36768 15936 36780
rect 15887 36740 15936 36768
rect 15887 36737 15899 36740
rect 15841 36731 15899 36737
rect 15930 36728 15936 36740
rect 15988 36728 15994 36780
rect 17494 36768 17500 36780
rect 17455 36740 17500 36768
rect 17494 36728 17500 36740
rect 17552 36728 17558 36780
rect 17681 36771 17739 36777
rect 17681 36737 17693 36771
rect 17727 36768 17739 36771
rect 18046 36768 18052 36780
rect 17727 36740 18052 36768
rect 17727 36737 17739 36740
rect 17681 36731 17739 36737
rect 18046 36728 18052 36740
rect 18104 36768 18110 36780
rect 18417 36771 18475 36777
rect 18417 36768 18429 36771
rect 18104 36740 18429 36768
rect 18104 36728 18110 36740
rect 18417 36737 18429 36740
rect 18463 36737 18475 36771
rect 18417 36731 18475 36737
rect 20257 36771 20315 36777
rect 20257 36737 20269 36771
rect 20303 36768 20315 36771
rect 20346 36768 20352 36780
rect 20303 36740 20352 36768
rect 20303 36737 20315 36740
rect 20257 36731 20315 36737
rect 14550 36700 14556 36712
rect 14200 36672 14556 36700
rect 14550 36660 14556 36672
rect 14608 36660 14614 36712
rect 15565 36703 15623 36709
rect 15565 36669 15577 36703
rect 15611 36669 15623 36703
rect 15672 36700 15700 36728
rect 17126 36700 17132 36712
rect 15672 36672 17132 36700
rect 15565 36663 15623 36669
rect 15580 36632 15608 36663
rect 17126 36660 17132 36672
rect 17184 36700 17190 36712
rect 17221 36703 17279 36709
rect 17221 36700 17233 36703
rect 17184 36672 17233 36700
rect 17184 36660 17190 36672
rect 17221 36669 17233 36672
rect 17267 36669 17279 36703
rect 17221 36663 17279 36669
rect 18138 36660 18144 36712
rect 18196 36700 18202 36712
rect 18233 36703 18291 36709
rect 18233 36700 18245 36703
rect 18196 36672 18245 36700
rect 18196 36660 18202 36672
rect 18233 36669 18245 36672
rect 18279 36700 18291 36703
rect 19242 36700 19248 36712
rect 18279 36672 19248 36700
rect 18279 36669 18291 36672
rect 18233 36663 18291 36669
rect 19242 36660 19248 36672
rect 19300 36660 19306 36712
rect 20272 36632 20300 36731
rect 20346 36728 20352 36740
rect 20404 36728 20410 36780
rect 20441 36771 20499 36777
rect 20441 36737 20453 36771
rect 20487 36768 20499 36771
rect 20806 36768 20812 36780
rect 20487 36740 20812 36768
rect 20487 36737 20499 36740
rect 20441 36731 20499 36737
rect 20806 36728 20812 36740
rect 20864 36728 20870 36780
rect 20901 36771 20959 36777
rect 20901 36737 20913 36771
rect 20947 36768 20959 36771
rect 22094 36768 22100 36780
rect 20947 36740 22100 36768
rect 20947 36737 20959 36740
rect 20901 36731 20959 36737
rect 22094 36728 22100 36740
rect 22152 36728 22158 36780
rect 22646 36728 22652 36780
rect 22704 36768 22710 36780
rect 22741 36771 22799 36777
rect 22741 36768 22753 36771
rect 22704 36740 22753 36768
rect 22704 36728 22710 36740
rect 22741 36737 22753 36740
rect 22787 36737 22799 36771
rect 22741 36731 22799 36737
rect 23106 36728 23112 36780
rect 23164 36768 23170 36780
rect 23385 36771 23443 36777
rect 23385 36768 23397 36771
rect 23164 36740 23397 36768
rect 23164 36728 23170 36740
rect 23385 36737 23397 36740
rect 23431 36768 23443 36771
rect 25314 36768 25320 36780
rect 23431 36740 25320 36768
rect 23431 36737 23443 36740
rect 23385 36731 23443 36737
rect 25314 36728 25320 36740
rect 25372 36728 25378 36780
rect 25424 36777 25452 36808
rect 29104 36808 29929 36836
rect 25409 36771 25467 36777
rect 25409 36737 25421 36771
rect 25455 36737 25467 36771
rect 26421 36771 26479 36777
rect 26421 36768 26433 36771
rect 25409 36731 25467 36737
rect 25700 36740 26433 36768
rect 25700 36712 25728 36740
rect 26421 36737 26433 36740
rect 26467 36768 26479 36771
rect 26878 36768 26884 36780
rect 26467 36740 26884 36768
rect 26467 36737 26479 36740
rect 26421 36731 26479 36737
rect 26878 36728 26884 36740
rect 26936 36728 26942 36780
rect 28445 36771 28503 36777
rect 28445 36737 28457 36771
rect 28491 36768 28503 36771
rect 28626 36768 28632 36780
rect 28491 36740 28632 36768
rect 28491 36737 28503 36740
rect 28445 36731 28503 36737
rect 28626 36728 28632 36740
rect 28684 36728 28690 36780
rect 29104 36777 29132 36808
rect 29917 36805 29929 36808
rect 29963 36805 29975 36839
rect 29917 36799 29975 36805
rect 36446 36796 36452 36848
rect 36504 36836 36510 36848
rect 36814 36836 36820 36848
rect 36504 36808 36820 36836
rect 36504 36796 36510 36808
rect 36814 36796 36820 36808
rect 36872 36836 36878 36848
rect 38197 36839 38255 36845
rect 38197 36836 38209 36839
rect 36872 36808 38209 36836
rect 36872 36796 36878 36808
rect 38197 36805 38209 36808
rect 38243 36805 38255 36839
rect 38197 36799 38255 36805
rect 38838 36796 38844 36848
rect 38896 36836 38902 36848
rect 39114 36836 39120 36848
rect 38896 36808 39120 36836
rect 38896 36796 38902 36808
rect 39114 36796 39120 36808
rect 39172 36836 39178 36848
rect 39390 36845 39396 36848
rect 39377 36839 39396 36845
rect 39172 36808 39344 36836
rect 39172 36796 39178 36808
rect 28905 36771 28963 36777
rect 28905 36737 28917 36771
rect 28951 36737 28963 36771
rect 28905 36731 28963 36737
rect 29089 36771 29147 36777
rect 29089 36737 29101 36771
rect 29135 36737 29147 36771
rect 29089 36731 29147 36737
rect 29733 36771 29791 36777
rect 29733 36737 29745 36771
rect 29779 36768 29791 36771
rect 30282 36768 30288 36780
rect 29779 36740 30288 36768
rect 29779 36737 29791 36740
rect 29733 36731 29791 36737
rect 22465 36703 22523 36709
rect 22465 36669 22477 36703
rect 22511 36700 22523 36703
rect 23290 36700 23296 36712
rect 22511 36672 23296 36700
rect 22511 36669 22523 36672
rect 22465 36663 22523 36669
rect 23290 36660 23296 36672
rect 23348 36660 23354 36712
rect 23477 36703 23535 36709
rect 23477 36669 23489 36703
rect 23523 36669 23535 36703
rect 24118 36700 24124 36712
rect 24079 36672 24124 36700
rect 23477 36663 23535 36669
rect 23492 36632 23520 36663
rect 24118 36660 24124 36672
rect 24176 36660 24182 36712
rect 24397 36703 24455 36709
rect 24397 36669 24409 36703
rect 24443 36669 24455 36703
rect 24397 36663 24455 36669
rect 24412 36632 24440 36663
rect 25222 36660 25228 36712
rect 25280 36700 25286 36712
rect 25501 36703 25559 36709
rect 25501 36700 25513 36703
rect 25280 36672 25513 36700
rect 25280 36660 25286 36672
rect 25501 36669 25513 36672
rect 25547 36700 25559 36703
rect 25682 36700 25688 36712
rect 25547 36672 25688 36700
rect 25547 36669 25559 36672
rect 25501 36663 25559 36669
rect 25682 36660 25688 36672
rect 25740 36660 25746 36712
rect 28920 36700 28948 36731
rect 29748 36700 29776 36731
rect 30282 36728 30288 36740
rect 30340 36728 30346 36780
rect 31202 36728 31208 36780
rect 31260 36768 31266 36780
rect 31481 36771 31539 36777
rect 31481 36768 31493 36771
rect 31260 36740 31493 36768
rect 31260 36728 31266 36740
rect 31481 36737 31493 36740
rect 31527 36737 31539 36771
rect 31481 36731 31539 36737
rect 32122 36728 32128 36780
rect 32180 36768 32186 36780
rect 35434 36777 35440 36780
rect 32401 36771 32459 36777
rect 32401 36768 32413 36771
rect 32180 36740 32413 36768
rect 32180 36728 32186 36740
rect 32401 36737 32413 36740
rect 32447 36737 32459 36771
rect 32401 36731 32459 36737
rect 35428 36731 35440 36777
rect 35492 36768 35498 36780
rect 35492 36740 35528 36768
rect 35434 36728 35440 36731
rect 35492 36728 35498 36740
rect 38286 36728 38292 36780
rect 38344 36768 38350 36780
rect 38381 36771 38439 36777
rect 38381 36768 38393 36771
rect 38344 36740 38393 36768
rect 38344 36728 38350 36740
rect 38381 36737 38393 36740
rect 38427 36737 38439 36771
rect 38381 36731 38439 36737
rect 38473 36771 38531 36777
rect 38473 36737 38485 36771
rect 38519 36768 38531 36771
rect 39206 36768 39212 36780
rect 38519 36740 39212 36768
rect 38519 36737 38531 36740
rect 38473 36731 38531 36737
rect 39206 36728 39212 36740
rect 39264 36728 39270 36780
rect 39316 36768 39344 36808
rect 39377 36805 39389 36839
rect 39377 36799 39396 36805
rect 39390 36796 39396 36799
rect 39448 36796 39454 36848
rect 39577 36839 39635 36845
rect 39577 36805 39589 36839
rect 39623 36805 39635 36839
rect 39577 36799 39635 36805
rect 39592 36768 39620 36799
rect 41598 36768 41604 36780
rect 39316 36740 39620 36768
rect 41386 36740 41604 36768
rect 28920 36672 29776 36700
rect 32677 36703 32735 36709
rect 32677 36669 32689 36703
rect 32723 36700 32735 36703
rect 32950 36700 32956 36712
rect 32723 36672 32956 36700
rect 32723 36669 32735 36672
rect 32677 36663 32735 36669
rect 32950 36660 32956 36672
rect 33008 36660 33014 36712
rect 34790 36660 34796 36712
rect 34848 36700 34854 36712
rect 35161 36703 35219 36709
rect 35161 36700 35173 36703
rect 34848 36672 35173 36700
rect 34848 36660 34854 36672
rect 35161 36669 35173 36672
rect 35207 36669 35219 36703
rect 41386 36700 41414 36740
rect 41598 36728 41604 36740
rect 41656 36728 41662 36780
rect 35161 36663 35219 36669
rect 36280 36672 41414 36700
rect 15580 36604 20300 36632
rect 22848 36604 25452 36632
rect 22848 36576 22876 36604
rect 5074 36524 5080 36576
rect 5132 36564 5138 36576
rect 5629 36567 5687 36573
rect 5629 36564 5641 36567
rect 5132 36536 5641 36564
rect 5132 36524 5138 36536
rect 5629 36533 5641 36536
rect 5675 36533 5687 36567
rect 14366 36564 14372 36576
rect 14327 36536 14372 36564
rect 5629 36527 5687 36533
rect 14366 36524 14372 36536
rect 14424 36524 14430 36576
rect 15746 36564 15752 36576
rect 15707 36536 15752 36564
rect 15746 36524 15752 36536
rect 15804 36524 15810 36576
rect 17310 36564 17316 36576
rect 17271 36536 17316 36564
rect 17310 36524 17316 36536
rect 17368 36524 17374 36576
rect 17494 36524 17500 36576
rect 17552 36564 17558 36576
rect 18506 36564 18512 36576
rect 17552 36536 18512 36564
rect 17552 36524 17558 36536
rect 18506 36524 18512 36536
rect 18564 36524 18570 36576
rect 21726 36524 21732 36576
rect 21784 36564 21790 36576
rect 22557 36567 22615 36573
rect 22557 36564 22569 36567
rect 21784 36536 22569 36564
rect 21784 36524 21790 36536
rect 22557 36533 22569 36536
rect 22603 36533 22615 36567
rect 22557 36527 22615 36533
rect 22649 36567 22707 36573
rect 22649 36533 22661 36567
rect 22695 36564 22707 36567
rect 22830 36564 22836 36576
rect 22695 36536 22836 36564
rect 22695 36533 22707 36536
rect 22649 36527 22707 36533
rect 22830 36524 22836 36536
rect 22888 36524 22894 36576
rect 23474 36564 23480 36576
rect 23435 36536 23480 36564
rect 23474 36524 23480 36536
rect 23532 36524 23538 36576
rect 25424 36573 25452 36604
rect 25409 36567 25467 36573
rect 25409 36533 25421 36567
rect 25455 36533 25467 36567
rect 25409 36527 25467 36533
rect 25590 36524 25596 36576
rect 25648 36564 25654 36576
rect 26329 36567 26387 36573
rect 26329 36564 26341 36567
rect 25648 36536 26341 36564
rect 25648 36524 25654 36536
rect 26329 36533 26341 36536
rect 26375 36533 26387 36567
rect 26329 36527 26387 36533
rect 33778 36524 33784 36576
rect 33836 36564 33842 36576
rect 36280 36564 36308 36672
rect 38749 36635 38807 36641
rect 38749 36601 38761 36635
rect 38795 36632 38807 36635
rect 38838 36632 38844 36644
rect 38795 36604 38844 36632
rect 38795 36601 38807 36604
rect 38749 36595 38807 36601
rect 38838 36592 38844 36604
rect 38896 36592 38902 36644
rect 33836 36536 36308 36564
rect 33836 36524 33842 36536
rect 39206 36524 39212 36576
rect 39264 36564 39270 36576
rect 39393 36567 39451 36573
rect 39393 36564 39405 36567
rect 39264 36536 39405 36564
rect 39264 36524 39270 36536
rect 39393 36533 39405 36536
rect 39439 36533 39451 36567
rect 39393 36527 39451 36533
rect 41693 36567 41751 36573
rect 41693 36533 41705 36567
rect 41739 36564 41751 36567
rect 41966 36564 41972 36576
rect 41739 36536 41972 36564
rect 41739 36533 41751 36536
rect 41693 36527 41751 36533
rect 41966 36524 41972 36536
rect 42024 36524 42030 36576
rect 1104 36474 42872 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 42872 36474
rect 1104 36400 42872 36422
rect 4890 36320 4896 36372
rect 4948 36360 4954 36372
rect 14458 36360 14464 36372
rect 4948 36332 14464 36360
rect 4948 36320 4954 36332
rect 14458 36320 14464 36332
rect 14516 36320 14522 36372
rect 15930 36360 15936 36372
rect 15891 36332 15936 36360
rect 15930 36320 15936 36332
rect 15988 36320 15994 36372
rect 16942 36360 16948 36372
rect 16903 36332 16948 36360
rect 16942 36320 16948 36332
rect 17000 36320 17006 36372
rect 17218 36360 17224 36372
rect 17179 36332 17224 36360
rect 17218 36320 17224 36332
rect 17276 36320 17282 36372
rect 17310 36320 17316 36372
rect 17368 36360 17374 36372
rect 17681 36363 17739 36369
rect 17681 36360 17693 36363
rect 17368 36332 17693 36360
rect 17368 36320 17374 36332
rect 17681 36329 17693 36332
rect 17727 36329 17739 36363
rect 21910 36360 21916 36372
rect 17681 36323 17739 36329
rect 17788 36332 18092 36360
rect 21871 36332 21916 36360
rect 4522 36252 4528 36304
rect 4580 36292 4586 36304
rect 4982 36292 4988 36304
rect 4580 36264 4988 36292
rect 4580 36252 4586 36264
rect 4982 36252 4988 36264
rect 5040 36252 5046 36304
rect 16850 36252 16856 36304
rect 16908 36292 16914 36304
rect 17788 36292 17816 36332
rect 16908 36264 17816 36292
rect 16908 36252 16914 36264
rect 16960 36233 16988 36264
rect 16945 36227 17003 36233
rect 16945 36193 16957 36227
rect 16991 36193 17003 36227
rect 16945 36187 17003 36193
rect 1946 36116 1952 36168
rect 2004 36156 2010 36168
rect 2041 36159 2099 36165
rect 2041 36156 2053 36159
rect 2004 36128 2053 36156
rect 2004 36116 2010 36128
rect 2041 36125 2053 36128
rect 2087 36125 2099 36159
rect 2041 36119 2099 36125
rect 2869 36159 2927 36165
rect 2869 36125 2881 36159
rect 2915 36125 2927 36159
rect 2869 36119 2927 36125
rect 4341 36159 4399 36165
rect 4341 36125 4353 36159
rect 4387 36156 4399 36159
rect 4614 36156 4620 36168
rect 4387 36128 4620 36156
rect 4387 36125 4399 36128
rect 4341 36119 4399 36125
rect 2774 36020 2780 36032
rect 2735 35992 2780 36020
rect 2774 35980 2780 35992
rect 2832 35980 2838 36032
rect 2884 36020 2912 36119
rect 4614 36116 4620 36128
rect 4672 36156 4678 36168
rect 5074 36156 5080 36168
rect 4672 36128 5080 36156
rect 4672 36116 4678 36128
rect 5074 36116 5080 36128
rect 5132 36116 5138 36168
rect 14090 36156 14096 36168
rect 14051 36128 14096 36156
rect 14090 36116 14096 36128
rect 14148 36116 14154 36168
rect 14366 36165 14372 36168
rect 14360 36156 14372 36165
rect 14327 36128 14372 36156
rect 14360 36119 14372 36128
rect 14366 36116 14372 36119
rect 14424 36116 14430 36168
rect 15654 36116 15660 36168
rect 15712 36156 15718 36168
rect 16117 36159 16175 36165
rect 16117 36156 16129 36159
rect 15712 36128 16129 36156
rect 15712 36116 15718 36128
rect 16117 36125 16129 36128
rect 16163 36125 16175 36159
rect 16117 36119 16175 36125
rect 16206 36116 16212 36168
rect 16264 36156 16270 36168
rect 16264 36128 16309 36156
rect 16264 36116 16270 36128
rect 16666 36116 16672 36168
rect 16724 36156 16730 36168
rect 16853 36159 16911 36165
rect 16853 36156 16865 36159
rect 16724 36128 16865 36156
rect 16724 36116 16730 36128
rect 16853 36125 16865 36128
rect 16899 36125 16911 36159
rect 16853 36119 16911 36125
rect 17865 36159 17923 36165
rect 17865 36125 17877 36159
rect 17911 36150 17923 36159
rect 17954 36150 17960 36168
rect 17911 36125 17960 36150
rect 17865 36122 17960 36125
rect 17865 36119 17923 36122
rect 17954 36116 17960 36122
rect 18012 36116 18018 36168
rect 18064 36165 18092 36332
rect 21910 36320 21916 36332
rect 21968 36320 21974 36372
rect 23753 36363 23811 36369
rect 23753 36329 23765 36363
rect 23799 36360 23811 36363
rect 23842 36360 23848 36372
rect 23799 36332 23848 36360
rect 23799 36329 23811 36332
rect 23753 36323 23811 36329
rect 23842 36320 23848 36332
rect 23900 36320 23906 36372
rect 24489 36363 24547 36369
rect 24489 36329 24501 36363
rect 24535 36360 24547 36363
rect 24762 36360 24768 36372
rect 24535 36332 24768 36360
rect 24535 36329 24547 36332
rect 24489 36323 24547 36329
rect 24762 36320 24768 36332
rect 24820 36320 24826 36372
rect 24854 36320 24860 36372
rect 24912 36360 24918 36372
rect 26602 36360 26608 36372
rect 24912 36332 24957 36360
rect 26563 36332 26608 36360
rect 24912 36320 24918 36332
rect 26602 36320 26608 36332
rect 26660 36320 26666 36372
rect 35894 36360 35900 36372
rect 35855 36332 35900 36360
rect 35894 36320 35900 36332
rect 35952 36320 35958 36372
rect 38838 36320 38844 36372
rect 38896 36360 38902 36372
rect 39025 36363 39083 36369
rect 39025 36360 39037 36363
rect 38896 36332 39037 36360
rect 38896 36320 38902 36332
rect 39025 36329 39037 36332
rect 39071 36360 39083 36363
rect 39390 36360 39396 36372
rect 39071 36332 39396 36360
rect 39071 36329 39083 36332
rect 39025 36323 39083 36329
rect 39390 36320 39396 36332
rect 39448 36320 39454 36372
rect 18230 36252 18236 36304
rect 18288 36292 18294 36304
rect 33778 36292 33784 36304
rect 18288 36264 33784 36292
rect 18288 36252 18294 36264
rect 33778 36252 33784 36264
rect 33836 36252 33842 36304
rect 33873 36295 33931 36301
rect 33873 36261 33885 36295
rect 33919 36292 33931 36295
rect 34514 36292 34520 36304
rect 33919 36264 34520 36292
rect 33919 36261 33931 36264
rect 33873 36255 33931 36261
rect 34514 36252 34520 36264
rect 34572 36252 34578 36304
rect 38381 36295 38439 36301
rect 38381 36261 38393 36295
rect 38427 36292 38439 36295
rect 39942 36292 39948 36304
rect 38427 36264 39948 36292
rect 38427 36261 38439 36264
rect 38381 36255 38439 36261
rect 39942 36252 39948 36264
rect 40000 36252 40006 36304
rect 18141 36227 18199 36233
rect 18141 36193 18153 36227
rect 18187 36224 18199 36227
rect 18322 36224 18328 36236
rect 18187 36196 18328 36224
rect 18187 36193 18199 36196
rect 18141 36187 18199 36193
rect 18322 36184 18328 36196
rect 18380 36184 18386 36236
rect 21726 36184 21732 36236
rect 21784 36224 21790 36236
rect 24302 36224 24308 36236
rect 21784 36196 22048 36224
rect 21784 36184 21790 36196
rect 18049 36159 18107 36165
rect 18049 36125 18061 36159
rect 18095 36156 18107 36159
rect 19242 36156 19248 36168
rect 18095 36128 19248 36156
rect 18095 36125 18107 36128
rect 18049 36119 18107 36125
rect 19242 36116 19248 36128
rect 19300 36116 19306 36168
rect 21082 36116 21088 36168
rect 21140 36156 21146 36168
rect 22020 36165 22048 36196
rect 22204 36196 24308 36224
rect 22204 36165 22232 36196
rect 24302 36184 24308 36196
rect 24360 36224 24366 36236
rect 24397 36227 24455 36233
rect 24397 36224 24409 36227
rect 24360 36196 24409 36224
rect 24360 36184 24366 36196
rect 24397 36193 24409 36196
rect 24443 36193 24455 36227
rect 24397 36187 24455 36193
rect 25866 36184 25872 36236
rect 25924 36224 25930 36236
rect 25961 36227 26019 36233
rect 25961 36224 25973 36227
rect 25924 36196 25973 36224
rect 25924 36184 25930 36196
rect 25961 36193 25973 36196
rect 26007 36193 26019 36227
rect 25961 36187 26019 36193
rect 32950 36184 32956 36236
rect 33008 36224 33014 36236
rect 33229 36227 33287 36233
rect 33229 36224 33241 36227
rect 33008 36196 33241 36224
rect 33008 36184 33014 36196
rect 33229 36193 33241 36196
rect 33275 36193 33287 36227
rect 33229 36187 33287 36193
rect 33413 36227 33471 36233
rect 33413 36193 33425 36227
rect 33459 36224 33471 36227
rect 35342 36224 35348 36236
rect 33459 36196 35348 36224
rect 33459 36193 33471 36196
rect 33413 36187 33471 36193
rect 21913 36159 21971 36165
rect 21913 36156 21925 36159
rect 21140 36128 21925 36156
rect 21140 36116 21146 36128
rect 21913 36125 21925 36128
rect 21959 36125 21971 36159
rect 21913 36119 21971 36125
rect 22005 36159 22063 36165
rect 22005 36125 22017 36159
rect 22051 36125 22063 36159
rect 22005 36119 22063 36125
rect 22189 36159 22247 36165
rect 22189 36125 22201 36159
rect 22235 36125 22247 36159
rect 22189 36119 22247 36125
rect 23290 36116 23296 36168
rect 23348 36156 23354 36168
rect 23569 36159 23627 36165
rect 23569 36156 23581 36159
rect 23348 36128 23581 36156
rect 23348 36116 23354 36128
rect 23569 36125 23581 36128
rect 23615 36125 23627 36159
rect 23569 36119 23627 36125
rect 24673 36159 24731 36165
rect 24673 36125 24685 36159
rect 24719 36156 24731 36159
rect 25314 36156 25320 36168
rect 24719 36128 25320 36156
rect 24719 36125 24731 36128
rect 24673 36119 24731 36125
rect 4985 36091 5043 36097
rect 4985 36057 4997 36091
rect 5031 36088 5043 36091
rect 5166 36088 5172 36100
rect 5031 36060 5172 36088
rect 5031 36057 5043 36060
rect 4985 36051 5043 36057
rect 5166 36048 5172 36060
rect 5224 36088 5230 36100
rect 13078 36088 13084 36100
rect 5224 36060 13084 36088
rect 5224 36048 5230 36060
rect 13078 36048 13084 36060
rect 13136 36048 13142 36100
rect 18506 36048 18512 36100
rect 18564 36088 18570 36100
rect 18564 36060 22094 36088
rect 18564 36048 18570 36060
rect 7466 36020 7472 36032
rect 2884 35992 7472 36020
rect 7466 35980 7472 35992
rect 7524 35980 7530 36032
rect 15470 36020 15476 36032
rect 15431 35992 15476 36020
rect 15470 35980 15476 35992
rect 15528 35980 15534 36032
rect 16206 35980 16212 36032
rect 16264 36020 16270 36032
rect 19337 36023 19395 36029
rect 19337 36020 19349 36023
rect 16264 35992 19349 36020
rect 16264 35980 16270 35992
rect 19337 35989 19349 35992
rect 19383 36020 19395 36023
rect 19426 36020 19432 36032
rect 19383 35992 19432 36020
rect 19383 35989 19395 35992
rect 19337 35983 19395 35989
rect 19426 35980 19432 35992
rect 19484 35980 19490 36032
rect 22066 36020 22094 36060
rect 22646 36048 22652 36100
rect 22704 36088 22710 36100
rect 23385 36091 23443 36097
rect 23385 36088 23397 36091
rect 22704 36060 23397 36088
rect 22704 36048 22710 36060
rect 23385 36057 23397 36060
rect 23431 36057 23443 36091
rect 23385 36051 23443 36057
rect 24688 36020 24716 36119
rect 25314 36116 25320 36128
rect 25372 36116 25378 36168
rect 25682 36156 25688 36168
rect 25643 36128 25688 36156
rect 25682 36116 25688 36128
rect 25740 36116 25746 36168
rect 25777 36159 25835 36165
rect 25777 36125 25789 36159
rect 25823 36156 25835 36159
rect 26050 36156 26056 36168
rect 25823 36128 26056 36156
rect 25823 36125 25835 36128
rect 25777 36119 25835 36125
rect 26050 36116 26056 36128
rect 26108 36116 26114 36168
rect 26418 36156 26424 36168
rect 26379 36128 26424 36156
rect 26418 36116 26424 36128
rect 26476 36116 26482 36168
rect 29730 36156 29736 36168
rect 29691 36128 29736 36156
rect 29730 36116 29736 36128
rect 29788 36116 29794 36168
rect 30650 36156 30656 36168
rect 30611 36128 30656 36156
rect 30650 36116 30656 36128
rect 30708 36116 30714 36168
rect 30742 36116 30748 36168
rect 30800 36156 30806 36168
rect 33134 36156 33140 36168
rect 30800 36128 30845 36156
rect 33095 36128 33140 36156
rect 30800 36116 30806 36128
rect 33134 36116 33140 36128
rect 33192 36116 33198 36168
rect 33244 36156 33272 36187
rect 35342 36184 35348 36196
rect 35400 36184 35406 36236
rect 38470 36224 38476 36236
rect 37476 36196 38476 36224
rect 34149 36159 34207 36165
rect 34149 36156 34161 36159
rect 33244 36128 34161 36156
rect 34149 36125 34161 36128
rect 34195 36125 34207 36159
rect 36538 36156 36544 36168
rect 36499 36128 36544 36156
rect 34149 36119 34207 36125
rect 36538 36116 36544 36128
rect 36596 36116 36602 36168
rect 36630 36116 36636 36168
rect 36688 36156 36694 36168
rect 36688 36128 36733 36156
rect 36688 36116 36694 36128
rect 36814 36116 36820 36168
rect 36872 36156 36878 36168
rect 37476 36165 37504 36196
rect 38470 36184 38476 36196
rect 38528 36184 38534 36236
rect 38841 36227 38899 36233
rect 38841 36193 38853 36227
rect 38887 36224 38899 36227
rect 39022 36224 39028 36236
rect 38887 36196 39028 36224
rect 38887 36193 38899 36196
rect 38841 36187 38899 36193
rect 39022 36184 39028 36196
rect 39080 36184 39086 36236
rect 41322 36224 41328 36236
rect 41283 36196 41328 36224
rect 41322 36184 41328 36196
rect 41380 36184 41386 36236
rect 41966 36224 41972 36236
rect 41927 36196 41972 36224
rect 41966 36184 41972 36196
rect 42024 36184 42030 36236
rect 37461 36159 37519 36165
rect 36872 36128 36917 36156
rect 36872 36116 36878 36128
rect 37461 36125 37473 36159
rect 37507 36125 37519 36159
rect 37461 36119 37519 36125
rect 38105 36159 38163 36165
rect 38105 36125 38117 36159
rect 38151 36156 38163 36159
rect 38746 36156 38752 36168
rect 38151 36128 38752 36156
rect 38151 36125 38163 36128
rect 38105 36119 38163 36125
rect 38746 36116 38752 36128
rect 38804 36116 38810 36168
rect 39114 36116 39120 36168
rect 39172 36156 39178 36168
rect 39172 36128 39217 36156
rect 39172 36116 39178 36128
rect 42150 36116 42156 36168
rect 42208 36156 42214 36168
rect 42208 36128 42253 36156
rect 42208 36116 42214 36128
rect 33413 36091 33471 36097
rect 33413 36057 33425 36091
rect 33459 36088 33471 36091
rect 33873 36091 33931 36097
rect 33873 36088 33885 36091
rect 33459 36060 33885 36088
rect 33459 36057 33471 36060
rect 33413 36051 33471 36057
rect 33873 36057 33885 36060
rect 33919 36057 33931 36091
rect 36078 36088 36084 36100
rect 36039 36060 36084 36088
rect 33873 36051 33931 36057
rect 36078 36048 36084 36060
rect 36136 36048 36142 36100
rect 38381 36091 38439 36097
rect 38381 36057 38393 36091
rect 38427 36088 38439 36091
rect 38841 36091 38899 36097
rect 38841 36088 38853 36091
rect 38427 36060 38853 36088
rect 38427 36057 38439 36060
rect 38381 36051 38439 36057
rect 38841 36057 38853 36060
rect 38887 36057 38899 36091
rect 38841 36051 38899 36057
rect 25682 36020 25688 36032
rect 22066 35992 24716 36020
rect 25643 35992 25688 36020
rect 25682 35980 25688 35992
rect 25740 35980 25746 36032
rect 29546 36020 29552 36032
rect 29507 35992 29552 36020
rect 29546 35980 29552 35992
rect 29604 35980 29610 36032
rect 30929 36023 30987 36029
rect 30929 35989 30941 36023
rect 30975 36020 30987 36023
rect 31754 36020 31760 36032
rect 30975 35992 31760 36020
rect 30975 35989 30987 35992
rect 30929 35983 30987 35989
rect 31754 35980 31760 35992
rect 31812 36020 31818 36032
rect 32398 36020 32404 36032
rect 31812 35992 32404 36020
rect 31812 35980 31818 35992
rect 32398 35980 32404 35992
rect 32456 35980 32462 36032
rect 33134 35980 33140 36032
rect 33192 36020 33198 36032
rect 34057 36023 34115 36029
rect 34057 36020 34069 36023
rect 33192 35992 34069 36020
rect 33192 35980 33198 35992
rect 34057 35989 34069 35992
rect 34103 35989 34115 36023
rect 35710 36020 35716 36032
rect 35671 35992 35716 36020
rect 34057 35983 34115 35989
rect 35710 35980 35716 35992
rect 35768 35980 35774 36032
rect 35881 36023 35939 36029
rect 35881 35989 35893 36023
rect 35927 36020 35939 36023
rect 36541 36023 36599 36029
rect 36541 36020 36553 36023
rect 35927 35992 36553 36020
rect 35927 35989 35939 35992
rect 35881 35983 35939 35989
rect 36541 35989 36553 35992
rect 36587 35989 36599 36023
rect 36541 35983 36599 35989
rect 37645 36023 37703 36029
rect 37645 35989 37657 36023
rect 37691 36020 37703 36023
rect 38197 36023 38255 36029
rect 38197 36020 38209 36023
rect 37691 35992 38209 36020
rect 37691 35989 37703 35992
rect 37645 35983 37703 35989
rect 38197 35989 38209 35992
rect 38243 36020 38255 36023
rect 39132 36020 39160 36116
rect 38243 35992 39160 36020
rect 38243 35989 38255 35992
rect 38197 35983 38255 35989
rect 1104 35930 42872 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 42872 35930
rect 1104 35856 42872 35878
rect 14274 35776 14280 35828
rect 14332 35816 14338 35828
rect 14553 35819 14611 35825
rect 14553 35816 14565 35819
rect 14332 35788 14565 35816
rect 14332 35776 14338 35788
rect 14553 35785 14565 35788
rect 14599 35785 14611 35819
rect 17126 35816 17132 35828
rect 17087 35788 17132 35816
rect 14553 35779 14611 35785
rect 17126 35776 17132 35788
rect 17184 35776 17190 35828
rect 24118 35776 24124 35828
rect 24176 35816 24182 35828
rect 24397 35819 24455 35825
rect 24397 35816 24409 35819
rect 24176 35788 24409 35816
rect 24176 35776 24182 35788
rect 24397 35785 24409 35788
rect 24443 35785 24455 35819
rect 24397 35779 24455 35785
rect 25498 35776 25504 35828
rect 25556 35816 25562 35828
rect 25556 35788 27384 35816
rect 25556 35776 25562 35788
rect 2133 35751 2191 35757
rect 2133 35717 2145 35751
rect 2179 35748 2191 35751
rect 2774 35748 2780 35760
rect 2179 35720 2780 35748
rect 2179 35717 2191 35720
rect 2133 35711 2191 35717
rect 2774 35708 2780 35720
rect 2832 35708 2838 35760
rect 15470 35708 15476 35760
rect 15528 35748 15534 35760
rect 15933 35751 15991 35757
rect 15933 35748 15945 35751
rect 15528 35720 15945 35748
rect 15528 35708 15534 35720
rect 15933 35717 15945 35720
rect 15979 35748 15991 35751
rect 24946 35748 24952 35760
rect 15979 35720 17632 35748
rect 15979 35717 15991 35720
rect 15933 35711 15991 35717
rect 1946 35680 1952 35692
rect 1907 35652 1952 35680
rect 1946 35640 1952 35652
rect 2004 35640 2010 35692
rect 5074 35680 5080 35692
rect 5035 35652 5080 35680
rect 5074 35640 5080 35652
rect 5132 35640 5138 35692
rect 14829 35683 14887 35689
rect 14829 35649 14841 35683
rect 14875 35680 14887 35683
rect 15286 35680 15292 35692
rect 14875 35652 15292 35680
rect 14875 35649 14887 35652
rect 14829 35643 14887 35649
rect 15286 35640 15292 35652
rect 15344 35640 15350 35692
rect 2866 35612 2872 35624
rect 2827 35584 2872 35612
rect 2866 35572 2872 35584
rect 2924 35572 2930 35624
rect 4798 35612 4804 35624
rect 4759 35584 4804 35612
rect 4798 35572 4804 35584
rect 4856 35572 4862 35624
rect 14553 35615 14611 35621
rect 14553 35581 14565 35615
rect 14599 35612 14611 35615
rect 15488 35612 15516 35708
rect 16117 35683 16175 35689
rect 16117 35680 16129 35683
rect 14599 35584 15516 35612
rect 15580 35652 16129 35680
rect 14599 35581 14611 35584
rect 14553 35575 14611 35581
rect 15286 35504 15292 35556
rect 15344 35544 15350 35556
rect 15580 35544 15608 35652
rect 16117 35649 16129 35652
rect 16163 35649 16175 35683
rect 16666 35680 16672 35692
rect 16627 35652 16672 35680
rect 16117 35643 16175 35649
rect 16666 35640 16672 35652
rect 16724 35640 16730 35692
rect 16761 35683 16819 35689
rect 16761 35649 16773 35683
rect 16807 35680 16819 35683
rect 16850 35680 16856 35692
rect 16807 35652 16856 35680
rect 16807 35649 16819 35652
rect 16761 35643 16819 35649
rect 16850 35640 16856 35652
rect 16908 35640 16914 35692
rect 16945 35683 17003 35689
rect 16945 35649 16957 35683
rect 16991 35680 17003 35683
rect 17218 35680 17224 35692
rect 16991 35652 17224 35680
rect 16991 35649 17003 35652
rect 16945 35643 17003 35649
rect 17218 35640 17224 35652
rect 17276 35640 17282 35692
rect 17604 35689 17632 35720
rect 19306 35720 19840 35748
rect 17589 35683 17647 35689
rect 17589 35649 17601 35683
rect 17635 35649 17647 35683
rect 17589 35643 17647 35649
rect 15749 35615 15807 35621
rect 15749 35581 15761 35615
rect 15795 35612 15807 35615
rect 16684 35612 16712 35640
rect 15795 35584 16712 35612
rect 16868 35612 16896 35640
rect 17954 35612 17960 35624
rect 16868 35584 17960 35612
rect 15795 35581 15807 35584
rect 15749 35575 15807 35581
rect 17954 35572 17960 35584
rect 18012 35612 18018 35624
rect 19306 35612 19334 35720
rect 19610 35680 19616 35692
rect 19571 35652 19616 35680
rect 19610 35640 19616 35652
rect 19668 35640 19674 35692
rect 19812 35689 19840 35720
rect 23952 35720 24952 35748
rect 19705 35683 19763 35689
rect 19705 35649 19717 35683
rect 19751 35649 19763 35683
rect 19705 35643 19763 35649
rect 19797 35683 19855 35689
rect 19797 35649 19809 35683
rect 19843 35649 19855 35683
rect 19797 35643 19855 35649
rect 19981 35683 20039 35689
rect 19981 35649 19993 35683
rect 20027 35680 20039 35683
rect 22925 35683 22983 35689
rect 20027 35652 22876 35680
rect 20027 35649 20039 35652
rect 19981 35643 20039 35649
rect 18012 35584 19334 35612
rect 18012 35572 18018 35584
rect 15344 35516 15608 35544
rect 19720 35544 19748 35643
rect 19812 35612 19840 35643
rect 22278 35612 22284 35624
rect 19812 35584 22284 35612
rect 22278 35572 22284 35584
rect 22336 35572 22342 35624
rect 22646 35612 22652 35624
rect 22607 35584 22652 35612
rect 22646 35572 22652 35584
rect 22704 35572 22710 35624
rect 22848 35612 22876 35652
rect 22925 35649 22937 35683
rect 22971 35680 22983 35683
rect 23474 35680 23480 35692
rect 22971 35652 23480 35680
rect 22971 35649 22983 35652
rect 22925 35643 22983 35649
rect 23474 35640 23480 35652
rect 23532 35680 23538 35692
rect 23952 35689 23980 35720
rect 24946 35708 24952 35720
rect 25004 35708 25010 35760
rect 25130 35708 25136 35760
rect 25188 35748 25194 35760
rect 25866 35748 25872 35760
rect 25188 35720 25872 35748
rect 25188 35708 25194 35720
rect 23937 35683 23995 35689
rect 23532 35652 23888 35680
rect 23532 35640 23538 35652
rect 23750 35612 23756 35624
rect 22848 35584 23756 35612
rect 23750 35572 23756 35584
rect 23808 35572 23814 35624
rect 20162 35544 20168 35556
rect 19720 35516 20168 35544
rect 15344 35504 15350 35516
rect 20162 35504 20168 35516
rect 20220 35504 20226 35556
rect 22554 35504 22560 35556
rect 22612 35544 22618 35556
rect 22830 35544 22836 35556
rect 22612 35516 22836 35544
rect 22612 35504 22618 35516
rect 22830 35504 22836 35516
rect 22888 35504 22894 35556
rect 14734 35476 14740 35488
rect 14695 35448 14740 35476
rect 14734 35436 14740 35448
rect 14792 35436 14798 35488
rect 17681 35479 17739 35485
rect 17681 35445 17693 35479
rect 17727 35476 17739 35479
rect 18322 35476 18328 35488
rect 17727 35448 18328 35476
rect 17727 35445 17739 35448
rect 17681 35439 17739 35445
rect 18322 35436 18328 35448
rect 18380 35436 18386 35488
rect 19058 35436 19064 35488
rect 19116 35476 19122 35488
rect 19337 35479 19395 35485
rect 19337 35476 19349 35479
rect 19116 35448 19349 35476
rect 19116 35436 19122 35448
rect 19337 35445 19349 35448
rect 19383 35445 19395 35479
rect 19337 35439 19395 35445
rect 22370 35436 22376 35488
rect 22428 35476 22434 35488
rect 23860 35485 23888 35652
rect 23937 35649 23949 35683
rect 23983 35649 23995 35683
rect 24394 35680 24400 35692
rect 24355 35652 24400 35680
rect 23937 35643 23995 35649
rect 24394 35640 24400 35652
rect 24452 35640 24458 35692
rect 24581 35683 24639 35689
rect 24581 35649 24593 35683
rect 24627 35680 24639 35683
rect 24762 35680 24768 35692
rect 24627 35652 24768 35680
rect 24627 35649 24639 35652
rect 24581 35643 24639 35649
rect 24762 35640 24768 35652
rect 24820 35640 24826 35692
rect 25222 35680 25228 35692
rect 25183 35652 25228 35680
rect 25222 35640 25228 35652
rect 25280 35640 25286 35692
rect 25424 35689 25452 35720
rect 25866 35708 25872 35720
rect 25924 35708 25930 35760
rect 25409 35683 25467 35689
rect 25409 35649 25421 35683
rect 25455 35649 25467 35683
rect 25409 35643 25467 35649
rect 25501 35683 25559 35689
rect 25501 35649 25513 35683
rect 25547 35649 25559 35683
rect 25501 35643 25559 35649
rect 25777 35683 25835 35689
rect 25777 35649 25789 35683
rect 25823 35680 25835 35683
rect 26970 35680 26976 35692
rect 25823 35652 26976 35680
rect 25823 35649 25835 35652
rect 25777 35643 25835 35649
rect 25516 35612 25544 35643
rect 26970 35640 26976 35652
rect 27028 35640 27034 35692
rect 27356 35689 27384 35788
rect 29730 35776 29736 35828
rect 29788 35816 29794 35828
rect 30285 35819 30343 35825
rect 30285 35816 30297 35819
rect 29788 35788 30297 35816
rect 29788 35776 29794 35788
rect 30285 35785 30297 35788
rect 30331 35785 30343 35819
rect 30285 35779 30343 35785
rect 32122 35776 32128 35828
rect 32180 35816 32186 35828
rect 32309 35819 32367 35825
rect 32309 35816 32321 35819
rect 32180 35788 32321 35816
rect 32180 35776 32186 35788
rect 32309 35785 32321 35788
rect 32355 35785 32367 35819
rect 32309 35779 32367 35785
rect 32398 35776 32404 35828
rect 32456 35816 32462 35828
rect 32456 35788 32501 35816
rect 32456 35776 32462 35788
rect 35434 35776 35440 35828
rect 35492 35816 35498 35828
rect 35621 35819 35679 35825
rect 35621 35816 35633 35819
rect 35492 35788 35633 35816
rect 35492 35776 35498 35788
rect 35621 35785 35633 35788
rect 35667 35785 35679 35819
rect 35621 35779 35679 35785
rect 28712 35751 28770 35757
rect 28712 35717 28724 35751
rect 28758 35748 28770 35751
rect 29546 35748 29552 35760
rect 28758 35720 29552 35748
rect 28758 35717 28770 35720
rect 28712 35711 28770 35717
rect 29546 35708 29552 35720
rect 29604 35708 29610 35760
rect 30469 35751 30527 35757
rect 30469 35717 30481 35751
rect 30515 35748 30527 35751
rect 30834 35748 30840 35760
rect 30515 35720 30840 35748
rect 30515 35717 30527 35720
rect 30469 35711 30527 35717
rect 30834 35708 30840 35720
rect 30892 35708 30898 35760
rect 34514 35708 34520 35760
rect 34572 35757 34578 35760
rect 34572 35748 34584 35757
rect 34572 35720 34617 35748
rect 34572 35711 34584 35720
rect 34572 35708 34578 35711
rect 39942 35708 39948 35760
rect 40000 35748 40006 35760
rect 40098 35751 40156 35757
rect 40098 35748 40110 35751
rect 40000 35720 40110 35748
rect 40000 35708 40006 35720
rect 40098 35717 40110 35720
rect 40144 35717 40156 35751
rect 40098 35711 40156 35717
rect 27341 35683 27399 35689
rect 27341 35649 27353 35683
rect 27387 35649 27399 35683
rect 28442 35680 28448 35692
rect 28403 35652 28448 35680
rect 27341 35643 27399 35649
rect 28442 35640 28448 35652
rect 28500 35640 28506 35692
rect 32030 35640 32036 35692
rect 32088 35680 32094 35692
rect 32493 35683 32551 35689
rect 32493 35680 32505 35683
rect 32088 35652 32505 35680
rect 32088 35640 32094 35652
rect 32493 35649 32505 35652
rect 32539 35649 32551 35683
rect 32493 35643 32551 35649
rect 35710 35640 35716 35692
rect 35768 35680 35774 35692
rect 35805 35683 35863 35689
rect 35805 35680 35817 35683
rect 35768 35652 35817 35680
rect 35768 35640 35774 35652
rect 35805 35649 35817 35652
rect 35851 35649 35863 35683
rect 35805 35643 35863 35649
rect 41877 35683 41935 35689
rect 41877 35649 41889 35683
rect 41923 35680 41935 35683
rect 42150 35680 42156 35692
rect 41923 35652 42156 35680
rect 41923 35649 41935 35652
rect 41877 35643 41935 35649
rect 42150 35640 42156 35652
rect 42208 35640 42214 35692
rect 25958 35612 25964 35624
rect 25516 35584 25964 35612
rect 25958 35572 25964 35584
rect 26016 35572 26022 35624
rect 26050 35572 26056 35624
rect 26108 35612 26114 35624
rect 27249 35615 27307 35621
rect 27249 35612 27261 35615
rect 26108 35584 27261 35612
rect 26108 35572 26114 35584
rect 27249 35581 27261 35584
rect 27295 35581 27307 35615
rect 34790 35612 34796 35624
rect 34751 35584 34796 35612
rect 27249 35575 27307 35581
rect 34790 35572 34796 35584
rect 34848 35572 34854 35624
rect 38286 35572 38292 35624
rect 38344 35612 38350 35624
rect 38565 35615 38623 35621
rect 38565 35612 38577 35615
rect 38344 35584 38577 35612
rect 38344 35572 38350 35584
rect 38565 35581 38577 35584
rect 38611 35581 38623 35615
rect 38838 35612 38844 35624
rect 38799 35584 38844 35612
rect 38565 35575 38623 35581
rect 38838 35572 38844 35584
rect 38896 35572 38902 35624
rect 38930 35572 38936 35624
rect 38988 35612 38994 35624
rect 39853 35615 39911 35621
rect 39853 35612 39865 35615
rect 38988 35584 39865 35612
rect 38988 35572 38994 35584
rect 39853 35581 39865 35584
rect 39899 35581 39911 35615
rect 39853 35575 39911 35581
rect 25593 35547 25651 35553
rect 25593 35513 25605 35547
rect 25639 35544 25651 35547
rect 26602 35544 26608 35556
rect 25639 35516 26608 35544
rect 25639 35513 25651 35516
rect 25593 35507 25651 35513
rect 26602 35504 26608 35516
rect 26660 35504 26666 35556
rect 29825 35547 29883 35553
rect 29825 35513 29837 35547
rect 29871 35544 29883 35547
rect 30650 35544 30656 35556
rect 29871 35516 30656 35544
rect 29871 35513 29883 35516
rect 29825 35507 29883 35513
rect 30650 35504 30656 35516
rect 30708 35504 30714 35556
rect 30837 35547 30895 35553
rect 30837 35513 30849 35547
rect 30883 35544 30895 35547
rect 31386 35544 31392 35556
rect 30883 35516 31392 35544
rect 30883 35513 30895 35516
rect 30837 35507 30895 35513
rect 31386 35504 31392 35516
rect 31444 35544 31450 35556
rect 32125 35547 32183 35553
rect 32125 35544 32137 35547
rect 31444 35516 32137 35544
rect 31444 35504 31450 35516
rect 32125 35513 32137 35516
rect 32171 35513 32183 35547
rect 32125 35507 32183 35513
rect 32677 35547 32735 35553
rect 32677 35513 32689 35547
rect 32723 35544 32735 35547
rect 32766 35544 32772 35556
rect 32723 35516 32772 35544
rect 32723 35513 32735 35516
rect 32677 35507 32735 35513
rect 32766 35504 32772 35516
rect 32824 35544 32830 35556
rect 33413 35547 33471 35553
rect 33413 35544 33425 35547
rect 32824 35516 33425 35544
rect 32824 35504 32830 35516
rect 33413 35513 33425 35516
rect 33459 35513 33471 35547
rect 33413 35507 33471 35513
rect 22741 35479 22799 35485
rect 22741 35476 22753 35479
rect 22428 35448 22753 35476
rect 22428 35436 22434 35448
rect 22741 35445 22753 35448
rect 22787 35445 22799 35479
rect 22741 35439 22799 35445
rect 23845 35479 23903 35485
rect 23845 35445 23857 35479
rect 23891 35476 23903 35479
rect 23934 35476 23940 35488
rect 23891 35448 23940 35476
rect 23891 35445 23903 35448
rect 23845 35439 23903 35445
rect 23934 35436 23940 35448
rect 23992 35436 23998 35488
rect 25685 35479 25743 35485
rect 25685 35445 25697 35479
rect 25731 35476 25743 35479
rect 25774 35476 25780 35488
rect 25731 35448 25780 35476
rect 25731 35445 25743 35448
rect 25685 35439 25743 35445
rect 25774 35436 25780 35448
rect 25832 35436 25838 35488
rect 26142 35436 26148 35488
rect 26200 35476 26206 35488
rect 26973 35479 27031 35485
rect 26973 35476 26985 35479
rect 26200 35448 26985 35476
rect 26200 35436 26206 35448
rect 26973 35445 26985 35448
rect 27019 35445 27031 35479
rect 26973 35439 27031 35445
rect 30469 35479 30527 35485
rect 30469 35445 30481 35479
rect 30515 35476 30527 35479
rect 30926 35476 30932 35488
rect 30515 35448 30932 35476
rect 30515 35445 30527 35448
rect 30469 35439 30527 35445
rect 30926 35436 30932 35448
rect 30984 35476 30990 35488
rect 36078 35476 36084 35488
rect 30984 35448 36084 35476
rect 30984 35436 30990 35448
rect 36078 35436 36084 35448
rect 36136 35436 36142 35488
rect 38470 35436 38476 35488
rect 38528 35476 38534 35488
rect 41233 35479 41291 35485
rect 41233 35476 41245 35479
rect 38528 35448 41245 35476
rect 38528 35436 38534 35448
rect 41233 35445 41245 35448
rect 41279 35445 41291 35479
rect 41233 35439 41291 35445
rect 1104 35386 42872 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 42872 35386
rect 1104 35312 42872 35334
rect 15565 35275 15623 35281
rect 15565 35241 15577 35275
rect 15611 35272 15623 35275
rect 15746 35272 15752 35284
rect 15611 35244 15752 35272
rect 15611 35241 15623 35244
rect 15565 35235 15623 35241
rect 15746 35232 15752 35244
rect 15804 35232 15810 35284
rect 19610 35232 19616 35284
rect 19668 35272 19674 35284
rect 19889 35275 19947 35281
rect 19889 35272 19901 35275
rect 19668 35244 19901 35272
rect 19668 35232 19674 35244
rect 19889 35241 19901 35244
rect 19935 35241 19947 35275
rect 19889 35235 19947 35241
rect 22738 35232 22744 35284
rect 22796 35272 22802 35284
rect 23201 35275 23259 35281
rect 23201 35272 23213 35275
rect 22796 35244 23213 35272
rect 22796 35232 22802 35244
rect 23201 35241 23213 35244
rect 23247 35241 23259 35275
rect 24762 35272 24768 35284
rect 24723 35244 24768 35272
rect 23201 35235 23259 35241
rect 24762 35232 24768 35244
rect 24820 35232 24826 35284
rect 24857 35275 24915 35281
rect 24857 35241 24869 35275
rect 24903 35272 24915 35275
rect 25682 35272 25688 35284
rect 24903 35244 25688 35272
rect 24903 35241 24915 35244
rect 24857 35235 24915 35241
rect 25682 35232 25688 35244
rect 25740 35232 25746 35284
rect 25792 35244 30512 35272
rect 16666 35204 16672 35216
rect 15580 35176 16672 35204
rect 15580 35077 15608 35176
rect 16666 35164 16672 35176
rect 16724 35164 16730 35216
rect 24946 35204 24952 35216
rect 24688 35176 24952 35204
rect 15749 35139 15807 35145
rect 15749 35105 15761 35139
rect 15795 35136 15807 35139
rect 16942 35136 16948 35148
rect 15795 35108 16948 35136
rect 15795 35105 15807 35108
rect 15749 35099 15807 35105
rect 15565 35071 15623 35077
rect 15565 35037 15577 35071
rect 15611 35037 15623 35071
rect 15565 35031 15623 35037
rect 15470 34960 15476 35012
rect 15528 35000 15534 35012
rect 15764 35000 15792 35099
rect 16942 35096 16948 35108
rect 17000 35096 17006 35148
rect 18230 35096 18236 35148
rect 18288 35136 18294 35148
rect 18414 35136 18420 35148
rect 18288 35108 18420 35136
rect 18288 35096 18294 35108
rect 18414 35096 18420 35108
rect 18472 35096 18478 35148
rect 18693 35139 18751 35145
rect 18693 35105 18705 35139
rect 18739 35136 18751 35139
rect 19978 35136 19984 35148
rect 18739 35108 19288 35136
rect 18739 35105 18751 35108
rect 18693 35099 18751 35105
rect 15841 35071 15899 35077
rect 15841 35037 15853 35071
rect 15887 35068 15899 35071
rect 16666 35068 16672 35080
rect 15887 35040 16672 35068
rect 15887 35037 15899 35040
rect 15841 35031 15899 35037
rect 16666 35028 16672 35040
rect 16724 35028 16730 35080
rect 17218 35068 17224 35080
rect 17179 35040 17224 35068
rect 17218 35028 17224 35040
rect 17276 35028 17282 35080
rect 19260 35077 19288 35108
rect 19628 35108 19984 35136
rect 18325 35071 18383 35077
rect 18325 35037 18337 35071
rect 18371 35037 18383 35071
rect 18325 35031 18383 35037
rect 19245 35071 19303 35077
rect 19245 35037 19257 35071
rect 19291 35037 19303 35071
rect 19245 35031 19303 35037
rect 19393 35071 19451 35077
rect 19393 35037 19405 35071
rect 19439 35068 19451 35071
rect 19628 35068 19656 35108
rect 19978 35096 19984 35108
rect 20036 35096 20042 35148
rect 21818 35136 21824 35148
rect 21779 35108 21824 35136
rect 21818 35096 21824 35108
rect 21876 35096 21882 35148
rect 24688 35145 24716 35176
rect 24946 35164 24952 35176
rect 25004 35164 25010 35216
rect 25792 35204 25820 35244
rect 25056 35176 25820 35204
rect 30484 35204 30512 35244
rect 30558 35232 30564 35284
rect 30616 35272 30622 35284
rect 30742 35272 30748 35284
rect 30616 35244 30748 35272
rect 30616 35232 30622 35244
rect 30742 35232 30748 35244
rect 30800 35272 30806 35284
rect 30929 35275 30987 35281
rect 30929 35272 30941 35275
rect 30800 35244 30941 35272
rect 30800 35232 30806 35244
rect 30929 35241 30941 35244
rect 30975 35272 30987 35275
rect 31202 35272 31208 35284
rect 30975 35244 31208 35272
rect 30975 35241 30987 35244
rect 30929 35235 30987 35241
rect 31202 35232 31208 35244
rect 31260 35232 31266 35284
rect 31726 35244 41368 35272
rect 31726 35204 31754 35244
rect 30484 35176 31754 35204
rect 24673 35139 24731 35145
rect 24673 35105 24685 35139
rect 24719 35105 24731 35139
rect 25056 35136 25084 35176
rect 38010 35164 38016 35216
rect 38068 35204 38074 35216
rect 38657 35207 38715 35213
rect 38657 35204 38669 35207
rect 38068 35176 38669 35204
rect 38068 35164 38074 35176
rect 38657 35173 38669 35176
rect 38703 35173 38715 35207
rect 38657 35167 38715 35173
rect 40037 35207 40095 35213
rect 40037 35173 40049 35207
rect 40083 35204 40095 35207
rect 40126 35204 40132 35216
rect 40083 35176 40132 35204
rect 40083 35173 40095 35176
rect 40037 35167 40095 35173
rect 40126 35164 40132 35176
rect 40184 35164 40190 35216
rect 24673 35099 24731 35105
rect 24780 35108 25084 35136
rect 19439 35040 19656 35068
rect 19439 35037 19451 35040
rect 19393 35031 19451 35037
rect 15528 34972 15792 35000
rect 15933 35003 15991 35009
rect 15528 34960 15534 34972
rect 15933 34969 15945 35003
rect 15979 35000 15991 35003
rect 16206 35000 16212 35012
rect 15979 34972 16212 35000
rect 15979 34969 15991 34972
rect 15933 34963 15991 34969
rect 16206 34960 16212 34972
rect 16264 34960 16270 35012
rect 18340 34932 18368 35031
rect 19702 35028 19708 35080
rect 19760 35077 19766 35080
rect 19760 35068 19768 35077
rect 21836 35068 21864 35096
rect 22646 35068 22652 35080
rect 19760 35040 19805 35068
rect 21836 35040 22652 35068
rect 19760 35031 19768 35040
rect 19760 35028 19766 35031
rect 22646 35028 22652 35040
rect 22704 35028 22710 35080
rect 23382 35028 23388 35080
rect 23440 35068 23446 35080
rect 24780 35068 24808 35108
rect 25774 35096 25780 35148
rect 25832 35136 25838 35148
rect 25832 35108 26832 35136
rect 25832 35096 25838 35108
rect 24946 35068 24952 35080
rect 23440 35040 24808 35068
rect 24907 35040 24952 35068
rect 23440 35028 23446 35040
rect 24946 35028 24952 35040
rect 25004 35028 25010 35080
rect 25590 35028 25596 35080
rect 25648 35077 25654 35080
rect 25648 35071 25697 35077
rect 25648 35037 25651 35071
rect 25685 35037 25697 35071
rect 25866 35068 25872 35080
rect 25827 35040 25872 35068
rect 25648 35031 25697 35037
rect 25648 35028 25654 35031
rect 25866 35028 25872 35040
rect 25924 35028 25930 35080
rect 25958 35028 25964 35080
rect 26016 35077 26022 35080
rect 26016 35071 26055 35077
rect 26043 35037 26055 35071
rect 26016 35031 26055 35037
rect 26016 35028 26022 35031
rect 26142 35028 26148 35080
rect 26200 35068 26206 35080
rect 26602 35068 26608 35080
rect 26200 35040 26245 35068
rect 26563 35040 26608 35068
rect 26200 35028 26206 35040
rect 26602 35028 26608 35040
rect 26660 35028 26666 35080
rect 26698 35071 26756 35077
rect 26698 35037 26710 35071
rect 26744 35037 26756 35071
rect 26804 35068 26832 35108
rect 28442 35096 28448 35148
rect 28500 35136 28506 35148
rect 28902 35136 28908 35148
rect 28500 35108 28908 35136
rect 28500 35096 28506 35108
rect 28902 35096 28908 35108
rect 28960 35136 28966 35148
rect 29549 35139 29607 35145
rect 29549 35136 29561 35139
rect 28960 35108 29561 35136
rect 28960 35096 28966 35108
rect 29549 35105 29561 35108
rect 29595 35105 29607 35139
rect 32766 35136 32772 35148
rect 32727 35108 32772 35136
rect 29549 35099 29607 35105
rect 32766 35096 32772 35108
rect 32824 35096 32830 35148
rect 34790 35096 34796 35148
rect 34848 35136 34854 35148
rect 34848 35108 36952 35136
rect 34848 35096 34854 35108
rect 27070 35071 27128 35077
rect 27070 35068 27082 35071
rect 26804 35040 27082 35068
rect 26698 35031 26756 35037
rect 27070 35037 27082 35040
rect 27116 35037 27128 35071
rect 32030 35068 32036 35080
rect 31991 35040 32036 35068
rect 27070 35031 27128 35037
rect 18414 34960 18420 35012
rect 18472 35000 18478 35012
rect 19521 35003 19579 35009
rect 19521 35000 19533 35003
rect 18472 34972 19533 35000
rect 18472 34960 18478 34972
rect 19521 34969 19533 34972
rect 19567 34969 19579 35003
rect 19521 34963 19579 34969
rect 19613 35003 19671 35009
rect 19613 34969 19625 35003
rect 19659 35000 19671 35003
rect 20070 35000 20076 35012
rect 19659 34972 20076 35000
rect 19659 34969 19671 34972
rect 19613 34963 19671 34969
rect 20070 34960 20076 34972
rect 20128 34960 20134 35012
rect 22088 35003 22146 35009
rect 22088 34969 22100 35003
rect 22134 35000 22146 35003
rect 22186 35000 22192 35012
rect 22134 34972 22192 35000
rect 22134 34969 22146 34972
rect 22088 34963 22146 34969
rect 22186 34960 22192 34972
rect 22244 34960 22250 35012
rect 25777 35003 25835 35009
rect 25777 34969 25789 35003
rect 25823 35000 25835 35003
rect 26418 35000 26424 35012
rect 25823 34972 26424 35000
rect 25823 34969 25835 34972
rect 25777 34963 25835 34969
rect 26418 34960 26424 34972
rect 26476 34960 26482 35012
rect 26510 34960 26516 35012
rect 26568 35000 26574 35012
rect 26712 35000 26740 35031
rect 32030 35028 32036 35040
rect 32088 35028 32094 35080
rect 32309 35071 32367 35077
rect 32309 35037 32321 35071
rect 32355 35068 32367 35071
rect 32950 35068 32956 35080
rect 32355 35040 32956 35068
rect 32355 35037 32367 35040
rect 32309 35031 32367 35037
rect 32950 35028 32956 35040
rect 33008 35028 33014 35080
rect 33045 35071 33103 35077
rect 33045 35037 33057 35071
rect 33091 35037 33103 35071
rect 35526 35068 35532 35080
rect 35487 35040 35532 35068
rect 33045 35031 33103 35037
rect 26878 35000 26884 35012
rect 26568 34972 26740 35000
rect 26839 34972 26884 35000
rect 26568 34960 26574 34972
rect 26878 34960 26884 34972
rect 26936 34960 26942 35012
rect 26970 34960 26976 35012
rect 27028 35000 27034 35012
rect 29822 35009 29828 35012
rect 27028 34972 27073 35000
rect 27028 34960 27034 34972
rect 29816 34963 29828 35009
rect 29880 35000 29886 35012
rect 33060 35000 33088 35031
rect 35526 35028 35532 35040
rect 35584 35028 35590 35080
rect 35713 35071 35771 35077
rect 35713 35037 35725 35071
rect 35759 35068 35771 35071
rect 35894 35068 35900 35080
rect 35759 35040 35900 35068
rect 35759 35037 35771 35040
rect 35713 35031 35771 35037
rect 35894 35028 35900 35040
rect 35952 35028 35958 35080
rect 36924 35068 36952 35108
rect 38102 35096 38108 35148
rect 38160 35136 38166 35148
rect 38473 35139 38531 35145
rect 38473 35136 38485 35139
rect 38160 35108 38485 35136
rect 38160 35096 38166 35108
rect 38473 35105 38485 35108
rect 38519 35105 38531 35139
rect 38930 35136 38936 35148
rect 38473 35099 38531 35105
rect 38580 35108 38936 35136
rect 38013 35071 38071 35077
rect 38013 35068 38025 35071
rect 36924 35040 38025 35068
rect 38013 35037 38025 35040
rect 38059 35068 38071 35071
rect 38580 35068 38608 35108
rect 38930 35096 38936 35108
rect 38988 35096 38994 35148
rect 38746 35068 38752 35080
rect 38059 35040 38608 35068
rect 38707 35040 38752 35068
rect 38059 35037 38071 35040
rect 38013 35031 38071 35037
rect 38746 35028 38752 35040
rect 38804 35028 38810 35080
rect 38838 35028 38844 35080
rect 38896 35068 38902 35080
rect 39853 35071 39911 35077
rect 39853 35068 39865 35071
rect 38896 35040 39865 35068
rect 38896 35028 38902 35040
rect 39853 35037 39865 35040
rect 39899 35037 39911 35071
rect 39853 35031 39911 35037
rect 40037 35071 40095 35077
rect 40037 35037 40049 35071
rect 40083 35037 40095 35071
rect 40678 35068 40684 35080
rect 40639 35040 40684 35068
rect 40037 35031 40095 35037
rect 33134 35000 33140 35012
rect 29880 34972 29916 35000
rect 32508 34972 33140 35000
rect 29822 34960 29828 34963
rect 29880 34960 29886 34972
rect 32508 34944 32536 34972
rect 33134 34960 33140 34972
rect 33192 35000 33198 35012
rect 33502 35000 33508 35012
rect 33192 34972 33508 35000
rect 33192 34960 33198 34972
rect 33502 34960 33508 34972
rect 33560 34960 33566 35012
rect 37550 34960 37556 35012
rect 37608 35000 37614 35012
rect 37746 35003 37804 35009
rect 37746 35000 37758 35003
rect 37608 34972 37758 35000
rect 37608 34960 37614 34972
rect 37746 34969 37758 34972
rect 37792 34969 37804 35003
rect 37746 34963 37804 34969
rect 38473 35003 38531 35009
rect 38473 34969 38485 35003
rect 38519 35000 38531 35003
rect 40052 35000 40080 35031
rect 40678 35028 40684 35040
rect 40736 35028 40742 35080
rect 41340 35077 41368 35244
rect 41325 35071 41383 35077
rect 41325 35037 41337 35071
rect 41371 35037 41383 35071
rect 41966 35068 41972 35080
rect 41927 35040 41972 35068
rect 41325 35031 41383 35037
rect 41966 35028 41972 35040
rect 42024 35028 42030 35080
rect 38519 34972 40080 35000
rect 38519 34969 38531 34972
rect 38473 34963 38531 34969
rect 20254 34932 20260 34944
rect 18340 34904 20260 34932
rect 20254 34892 20260 34904
rect 20312 34892 20318 34944
rect 25501 34935 25559 34941
rect 25501 34901 25513 34935
rect 25547 34932 25559 34935
rect 25682 34932 25688 34944
rect 25547 34904 25688 34932
rect 25547 34901 25559 34904
rect 25501 34895 25559 34901
rect 25682 34892 25688 34904
rect 25740 34892 25746 34944
rect 27246 34932 27252 34944
rect 27207 34904 27252 34932
rect 27246 34892 27252 34904
rect 27304 34892 27310 34944
rect 31846 34932 31852 34944
rect 31807 34904 31852 34932
rect 31846 34892 31852 34904
rect 31904 34892 31910 34944
rect 32217 34935 32275 34941
rect 32217 34901 32229 34935
rect 32263 34932 32275 34935
rect 32490 34932 32496 34944
rect 32263 34904 32496 34932
rect 32263 34901 32275 34904
rect 32217 34895 32275 34901
rect 32490 34892 32496 34904
rect 32548 34892 32554 34944
rect 35618 34932 35624 34944
rect 35579 34904 35624 34932
rect 35618 34892 35624 34904
rect 35676 34892 35682 34944
rect 36633 34935 36691 34941
rect 36633 34901 36645 34935
rect 36679 34932 36691 34935
rect 36814 34932 36820 34944
rect 36679 34904 36820 34932
rect 36679 34901 36691 34904
rect 36633 34895 36691 34901
rect 36814 34892 36820 34904
rect 36872 34892 36878 34944
rect 37274 34892 37280 34944
rect 37332 34932 37338 34944
rect 38102 34932 38108 34944
rect 37332 34904 38108 34932
rect 37332 34892 37338 34904
rect 38102 34892 38108 34904
rect 38160 34892 38166 34944
rect 40218 34892 40224 34944
rect 40276 34932 40282 34944
rect 41417 34935 41475 34941
rect 41417 34932 41429 34935
rect 40276 34904 41429 34932
rect 40276 34892 40282 34904
rect 41417 34901 41429 34904
rect 41463 34901 41475 34935
rect 41417 34895 41475 34901
rect 1104 34842 42872 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 42872 34842
rect 1104 34768 42872 34790
rect 4798 34688 4804 34740
rect 4856 34728 4862 34740
rect 16945 34731 17003 34737
rect 4856 34700 6914 34728
rect 4856 34688 4862 34700
rect 6886 34660 6914 34700
rect 16945 34697 16957 34731
rect 16991 34728 17003 34731
rect 17218 34728 17224 34740
rect 16991 34700 17224 34728
rect 16991 34697 17003 34700
rect 16945 34691 17003 34697
rect 17218 34688 17224 34700
rect 17276 34688 17282 34740
rect 22186 34728 22192 34740
rect 17328 34700 21373 34728
rect 22147 34700 22192 34728
rect 17328 34660 17356 34700
rect 6886 34632 17356 34660
rect 18966 34620 18972 34672
rect 19024 34660 19030 34672
rect 19426 34660 19432 34672
rect 19024 34632 19222 34660
rect 19387 34632 19432 34660
rect 19024 34620 19030 34632
rect 14461 34595 14519 34601
rect 14461 34561 14473 34595
rect 14507 34592 14519 34595
rect 14642 34592 14648 34604
rect 14507 34564 14648 34592
rect 14507 34561 14519 34564
rect 14461 34555 14519 34561
rect 14642 34552 14648 34564
rect 14700 34552 14706 34604
rect 14829 34595 14887 34601
rect 14829 34561 14841 34595
rect 14875 34592 14887 34595
rect 15470 34592 15476 34604
rect 14875 34564 15332 34592
rect 15431 34564 15476 34592
rect 14875 34561 14887 34564
rect 14829 34555 14887 34561
rect 15304 34536 15332 34564
rect 15470 34552 15476 34564
rect 15528 34552 15534 34604
rect 15565 34595 15623 34601
rect 15565 34561 15577 34595
rect 15611 34592 15623 34595
rect 16666 34592 16672 34604
rect 15611 34564 16672 34592
rect 15611 34561 15623 34564
rect 15565 34555 15623 34561
rect 16666 34552 16672 34564
rect 16724 34552 16730 34604
rect 18138 34592 18144 34604
rect 18099 34564 18144 34592
rect 18138 34552 18144 34564
rect 18196 34552 18202 34604
rect 18230 34552 18236 34604
rect 18288 34592 18294 34604
rect 18414 34592 18420 34604
rect 18288 34564 18333 34592
rect 18375 34564 18420 34592
rect 18288 34552 18294 34564
rect 18414 34552 18420 34564
rect 18472 34552 18478 34604
rect 18506 34552 18512 34604
rect 18564 34592 18570 34604
rect 19194 34601 19222 34632
rect 19426 34620 19432 34632
rect 19484 34620 19490 34672
rect 21345 34660 21373 34700
rect 22186 34688 22192 34700
rect 22244 34688 22250 34740
rect 30282 34728 30288 34740
rect 30195 34700 30288 34728
rect 30282 34688 30288 34700
rect 30340 34728 30346 34740
rect 30558 34728 30564 34740
rect 30340 34700 30564 34728
rect 30340 34688 30346 34700
rect 30558 34688 30564 34700
rect 30616 34688 30622 34740
rect 30834 34728 30840 34740
rect 30795 34700 30840 34728
rect 30834 34688 30840 34700
rect 30892 34688 30898 34740
rect 31202 34728 31208 34740
rect 31163 34700 31208 34728
rect 31202 34688 31208 34700
rect 31260 34688 31266 34740
rect 33137 34731 33195 34737
rect 33137 34728 33149 34731
rect 32140 34700 33149 34728
rect 22922 34660 22928 34672
rect 21345 34632 22928 34660
rect 22922 34620 22928 34632
rect 22980 34620 22986 34672
rect 25038 34620 25044 34672
rect 25096 34660 25102 34672
rect 27246 34660 27252 34672
rect 25096 34632 25544 34660
rect 25096 34620 25102 34632
rect 19068 34595 19126 34601
rect 19068 34592 19080 34595
rect 18564 34564 19080 34592
rect 18564 34552 18570 34564
rect 19068 34561 19080 34564
rect 19114 34561 19126 34595
rect 19068 34555 19126 34561
rect 19181 34595 19239 34601
rect 19181 34561 19193 34595
rect 19227 34561 19239 34595
rect 19181 34555 19239 34561
rect 19334 34552 19340 34604
rect 19392 34592 19398 34604
rect 19545 34595 19603 34601
rect 19392 34564 19485 34592
rect 19392 34552 19398 34564
rect 19545 34561 19557 34595
rect 19591 34592 19603 34595
rect 20898 34592 20904 34604
rect 19591 34561 19610 34592
rect 20859 34564 20904 34592
rect 19545 34555 19610 34561
rect 14553 34527 14611 34533
rect 14553 34493 14565 34527
rect 14599 34524 14611 34527
rect 14599 34496 15240 34524
rect 14599 34493 14611 34496
rect 14553 34487 14611 34493
rect 15212 34456 15240 34496
rect 15286 34484 15292 34536
rect 15344 34524 15350 34536
rect 15344 34496 15389 34524
rect 15344 34484 15350 34496
rect 15381 34459 15439 34465
rect 15381 34456 15393 34459
rect 15212 34428 15393 34456
rect 15381 34425 15393 34428
rect 15427 34425 15439 34459
rect 15381 34419 15439 34425
rect 14366 34388 14372 34400
rect 14327 34360 14372 34388
rect 14366 34348 14372 34360
rect 14424 34348 14430 34400
rect 14734 34388 14740 34400
rect 14647 34360 14740 34388
rect 14734 34348 14740 34360
rect 14792 34388 14798 34400
rect 15488 34388 15516 34552
rect 16574 34484 16580 34536
rect 16632 34524 16638 34536
rect 16945 34527 17003 34533
rect 16945 34524 16957 34527
rect 16632 34496 16957 34524
rect 16632 34484 16638 34496
rect 16945 34493 16957 34496
rect 16991 34493 17003 34527
rect 16945 34487 17003 34493
rect 18325 34527 18383 34533
rect 18325 34493 18337 34527
rect 18371 34524 18383 34527
rect 19352 34524 19380 34552
rect 19582 34524 19610 34555
rect 20898 34552 20904 34564
rect 20956 34552 20962 34604
rect 22370 34592 22376 34604
rect 22331 34564 22376 34592
rect 22370 34552 22376 34564
rect 22428 34552 22434 34604
rect 22554 34592 22560 34604
rect 22515 34564 22560 34592
rect 22554 34552 22560 34564
rect 22612 34552 22618 34604
rect 22649 34595 22707 34601
rect 22649 34561 22661 34595
rect 22695 34592 22707 34595
rect 22738 34592 22744 34604
rect 22695 34564 22744 34592
rect 22695 34561 22707 34564
rect 22649 34555 22707 34561
rect 22738 34552 22744 34564
rect 22796 34592 22802 34604
rect 23661 34595 23719 34601
rect 22796 34564 23612 34592
rect 22796 34552 22802 34564
rect 18371 34496 19380 34524
rect 19444 34496 19610 34524
rect 22281 34527 22339 34533
rect 18371 34493 18383 34496
rect 18325 34487 18383 34493
rect 16761 34459 16819 34465
rect 16761 34425 16773 34459
rect 16807 34456 16819 34459
rect 17957 34459 18015 34465
rect 17957 34456 17969 34459
rect 16807 34428 17969 34456
rect 16807 34425 16819 34428
rect 16761 34419 16819 34425
rect 17957 34425 17969 34428
rect 18003 34425 18015 34459
rect 17957 34419 18015 34425
rect 18138 34416 18144 34468
rect 18196 34456 18202 34468
rect 19444 34456 19472 34496
rect 22281 34493 22293 34527
rect 22327 34524 22339 34527
rect 22922 34524 22928 34536
rect 22327 34496 22928 34524
rect 22327 34493 22339 34496
rect 22281 34487 22339 34493
rect 22922 34484 22928 34496
rect 22980 34484 22986 34536
rect 23584 34533 23612 34564
rect 23661 34561 23673 34595
rect 23707 34592 23719 34595
rect 25130 34592 25136 34604
rect 23707 34564 25136 34592
rect 23707 34561 23719 34564
rect 23661 34555 23719 34561
rect 25130 34552 25136 34564
rect 25188 34552 25194 34604
rect 25516 34601 25544 34632
rect 25608 34632 27252 34660
rect 25608 34601 25636 34632
rect 27246 34620 27252 34632
rect 27304 34620 27310 34672
rect 30392 34632 31340 34660
rect 30392 34604 30420 34632
rect 25317 34595 25375 34601
rect 25317 34561 25329 34595
rect 25363 34561 25375 34595
rect 25317 34555 25375 34561
rect 25501 34595 25559 34601
rect 25501 34561 25513 34595
rect 25547 34561 25559 34595
rect 25501 34555 25559 34561
rect 25593 34595 25651 34601
rect 25593 34561 25605 34595
rect 25639 34561 25651 34595
rect 25593 34555 25651 34561
rect 23569 34527 23627 34533
rect 23569 34493 23581 34527
rect 23615 34493 23627 34527
rect 23569 34487 23627 34493
rect 23750 34484 23756 34536
rect 23808 34524 23814 34536
rect 24394 34524 24400 34536
rect 23808 34496 24400 34524
rect 23808 34484 23814 34496
rect 24394 34484 24400 34496
rect 24452 34524 24458 34536
rect 25332 34524 25360 34555
rect 25682 34552 25688 34604
rect 25740 34592 25746 34604
rect 25740 34564 25785 34592
rect 25740 34552 25746 34564
rect 26418 34552 26424 34604
rect 26476 34592 26482 34604
rect 27157 34595 27215 34601
rect 27157 34592 27169 34595
rect 26476 34564 27169 34592
rect 26476 34552 26482 34564
rect 27157 34561 27169 34564
rect 27203 34592 27215 34595
rect 27522 34592 27528 34604
rect 27203 34564 27528 34592
rect 27203 34561 27215 34564
rect 27157 34555 27215 34561
rect 27522 34552 27528 34564
rect 27580 34552 27586 34604
rect 29914 34592 29920 34604
rect 29875 34564 29920 34592
rect 29914 34552 29920 34564
rect 29972 34552 29978 34604
rect 30374 34552 30380 34604
rect 30432 34592 30438 34604
rect 30432 34564 30477 34592
rect 30432 34552 30438 34564
rect 30650 34552 30656 34604
rect 30708 34592 30714 34604
rect 31312 34601 31340 34632
rect 32140 34601 32168 34700
rect 33137 34697 33149 34700
rect 33183 34697 33195 34731
rect 33137 34691 33195 34697
rect 37921 34731 37979 34737
rect 37921 34697 37933 34731
rect 37967 34728 37979 34731
rect 38010 34728 38016 34740
rect 37967 34700 38016 34728
rect 37967 34697 37979 34700
rect 37921 34691 37979 34697
rect 38010 34688 38016 34700
rect 38068 34688 38074 34740
rect 39117 34731 39175 34737
rect 39117 34697 39129 34731
rect 39163 34728 39175 34731
rect 39206 34728 39212 34740
rect 39163 34700 39212 34728
rect 39163 34697 39175 34700
rect 39117 34691 39175 34697
rect 39206 34688 39212 34700
rect 39264 34688 39270 34740
rect 32493 34663 32551 34669
rect 32493 34629 32505 34663
rect 32539 34660 32551 34663
rect 32858 34660 32864 34672
rect 32539 34632 32864 34660
rect 32539 34629 32551 34632
rect 32493 34623 32551 34629
rect 32858 34620 32864 34632
rect 32916 34620 32922 34672
rect 32950 34620 32956 34672
rect 33008 34660 33014 34672
rect 33289 34663 33347 34669
rect 33289 34660 33301 34663
rect 33008 34632 33301 34660
rect 33008 34620 33014 34632
rect 33289 34629 33301 34632
rect 33335 34629 33347 34663
rect 33502 34660 33508 34672
rect 33463 34632 33508 34660
rect 33289 34623 33347 34629
rect 33502 34620 33508 34632
rect 33560 34620 33566 34672
rect 35060 34663 35118 34669
rect 35060 34629 35072 34663
rect 35106 34660 35118 34663
rect 35618 34660 35624 34672
rect 35106 34632 35624 34660
rect 35106 34629 35118 34632
rect 35060 34623 35118 34629
rect 35618 34620 35624 34632
rect 35676 34620 35682 34672
rect 36814 34620 36820 34672
rect 36872 34660 36878 34672
rect 37553 34663 37611 34669
rect 37553 34660 37565 34663
rect 36872 34632 37565 34660
rect 36872 34620 36878 34632
rect 37553 34629 37565 34632
rect 37599 34629 37611 34663
rect 37553 34623 37611 34629
rect 37758 34663 37816 34669
rect 37758 34629 37770 34663
rect 37804 34660 37816 34663
rect 38470 34660 38476 34672
rect 37804 34632 37872 34660
rect 38431 34632 38476 34660
rect 37804 34629 37816 34632
rect 37758 34623 37816 34629
rect 31021 34595 31079 34601
rect 31021 34592 31033 34595
rect 30708 34564 31033 34592
rect 30708 34552 30714 34564
rect 31021 34561 31033 34564
rect 31067 34561 31079 34595
rect 31021 34555 31079 34561
rect 31297 34595 31355 34601
rect 31297 34561 31309 34595
rect 31343 34592 31355 34595
rect 32125 34595 32183 34601
rect 32125 34592 32137 34595
rect 31343 34564 32137 34592
rect 31343 34561 31355 34564
rect 31297 34555 31355 34561
rect 32125 34561 32137 34564
rect 32171 34561 32183 34595
rect 34149 34595 34207 34601
rect 34149 34592 34161 34595
rect 32125 34555 32183 34561
rect 32692 34564 34161 34592
rect 24452 34496 25360 34524
rect 24452 34484 24458 34496
rect 25406 34484 25412 34536
rect 25464 34524 25470 34536
rect 25961 34527 26019 34533
rect 25961 34524 25973 34527
rect 25464 34496 25973 34524
rect 25464 34484 25470 34496
rect 25961 34493 25973 34496
rect 26007 34493 26019 34527
rect 25961 34487 26019 34493
rect 18196 34428 19472 34456
rect 19705 34459 19763 34465
rect 18196 34416 18202 34428
rect 19705 34425 19717 34459
rect 19751 34456 19763 34459
rect 20162 34456 20168 34468
rect 19751 34428 20168 34456
rect 19751 34425 19763 34428
rect 19705 34419 19763 34425
rect 20162 34416 20168 34428
rect 20220 34416 20226 34468
rect 24029 34459 24087 34465
rect 24029 34425 24041 34459
rect 24075 34456 24087 34459
rect 25222 34456 25228 34468
rect 24075 34428 25228 34456
rect 24075 34425 24087 34428
rect 24029 34419 24087 34425
rect 25222 34416 25228 34428
rect 25280 34416 25286 34468
rect 32030 34416 32036 34468
rect 32088 34456 32094 34468
rect 32692 34465 32720 34564
rect 34149 34561 34161 34564
rect 34195 34561 34207 34595
rect 34149 34555 34207 34561
rect 34514 34484 34520 34536
rect 34572 34524 34578 34536
rect 34790 34524 34796 34536
rect 34572 34496 34796 34524
rect 34572 34484 34578 34496
rect 34790 34484 34796 34496
rect 34848 34484 34854 34536
rect 37568 34524 37596 34623
rect 37844 34592 37872 34632
rect 38470 34620 38476 34632
rect 38528 34620 38534 34672
rect 40218 34660 40224 34672
rect 40179 34632 40224 34660
rect 40218 34620 40224 34632
rect 40276 34620 40282 34672
rect 41874 34660 41880 34672
rect 41835 34632 41880 34660
rect 41874 34620 41880 34632
rect 41932 34620 41938 34672
rect 38378 34592 38384 34604
rect 37844 34564 38384 34592
rect 38378 34552 38384 34564
rect 38436 34552 38442 34604
rect 38838 34592 38844 34604
rect 38672 34564 38844 34592
rect 38672 34524 38700 34564
rect 38838 34552 38844 34564
rect 38896 34592 38902 34604
rect 38933 34595 38991 34601
rect 38933 34592 38945 34595
rect 38896 34564 38945 34592
rect 38896 34552 38902 34564
rect 38933 34561 38945 34564
rect 38979 34561 38991 34595
rect 38933 34555 38991 34561
rect 37568 34496 38700 34524
rect 38746 34484 38752 34536
rect 38804 34524 38810 34536
rect 40037 34527 40095 34533
rect 38804 34496 38849 34524
rect 38804 34484 38810 34496
rect 40037 34493 40049 34527
rect 40083 34524 40095 34527
rect 40678 34524 40684 34536
rect 40083 34496 40684 34524
rect 40083 34493 40095 34496
rect 40037 34487 40095 34493
rect 40678 34484 40684 34496
rect 40736 34484 40742 34536
rect 32677 34459 32735 34465
rect 32088 34428 32628 34456
rect 32088 34416 32094 34428
rect 21082 34388 21088 34400
rect 14792 34360 15516 34388
rect 21043 34360 21088 34388
rect 14792 34348 14798 34360
rect 21082 34348 21088 34360
rect 21140 34348 21146 34400
rect 26510 34348 26516 34400
rect 26568 34388 26574 34400
rect 27065 34391 27123 34397
rect 27065 34388 27077 34391
rect 26568 34360 27077 34388
rect 26568 34348 26574 34360
rect 27065 34357 27077 34360
rect 27111 34357 27123 34391
rect 27065 34351 27123 34357
rect 30006 34348 30012 34400
rect 30064 34388 30070 34400
rect 30101 34391 30159 34397
rect 30101 34388 30113 34391
rect 30064 34360 30113 34388
rect 30064 34348 30070 34360
rect 30101 34357 30113 34360
rect 30147 34357 30159 34391
rect 30101 34351 30159 34357
rect 31846 34348 31852 34400
rect 31904 34388 31910 34400
rect 32493 34391 32551 34397
rect 32493 34388 32505 34391
rect 31904 34360 32505 34388
rect 31904 34348 31910 34360
rect 32493 34357 32505 34360
rect 32539 34357 32551 34391
rect 32600 34388 32628 34428
rect 32677 34425 32689 34459
rect 32723 34425 32735 34459
rect 32677 34419 32735 34425
rect 33321 34391 33379 34397
rect 33321 34388 33333 34391
rect 32600 34360 33333 34388
rect 32493 34351 32551 34357
rect 33321 34357 33333 34360
rect 33367 34357 33379 34391
rect 33962 34388 33968 34400
rect 33923 34360 33968 34388
rect 33321 34351 33379 34357
rect 33962 34348 33968 34360
rect 34020 34348 34026 34400
rect 36173 34391 36231 34397
rect 36173 34357 36185 34391
rect 36219 34388 36231 34391
rect 36262 34388 36268 34400
rect 36219 34360 36268 34388
rect 36219 34357 36231 34360
rect 36173 34351 36231 34357
rect 36262 34348 36268 34360
rect 36320 34388 36326 34400
rect 37737 34391 37795 34397
rect 37737 34388 37749 34391
rect 36320 34360 37749 34388
rect 36320 34348 36326 34360
rect 37737 34357 37749 34360
rect 37783 34388 37795 34391
rect 38654 34388 38660 34400
rect 37783 34360 38660 34388
rect 37783 34357 37795 34360
rect 37737 34351 37795 34357
rect 38654 34348 38660 34360
rect 38712 34348 38718 34400
rect 1104 34298 42872 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 42872 34298
rect 1104 34224 42872 34246
rect 18506 34184 18512 34196
rect 18467 34156 18512 34184
rect 18506 34144 18512 34156
rect 18564 34144 18570 34196
rect 18966 34144 18972 34196
rect 19024 34184 19030 34196
rect 20162 34184 20168 34196
rect 19024 34156 20168 34184
rect 19024 34144 19030 34156
rect 20162 34144 20168 34156
rect 20220 34144 20226 34196
rect 27154 34184 27160 34196
rect 27115 34156 27160 34184
rect 27154 34144 27160 34156
rect 27212 34144 27218 34196
rect 29822 34184 29828 34196
rect 29783 34156 29828 34184
rect 29822 34144 29828 34156
rect 29880 34144 29886 34196
rect 30193 34187 30251 34193
rect 30193 34153 30205 34187
rect 30239 34184 30251 34187
rect 30374 34184 30380 34196
rect 30239 34156 30380 34184
rect 30239 34153 30251 34156
rect 30193 34147 30251 34153
rect 30374 34144 30380 34156
rect 30432 34144 30438 34196
rect 31941 34187 31999 34193
rect 31941 34153 31953 34187
rect 31987 34184 31999 34187
rect 32030 34184 32036 34196
rect 31987 34156 32036 34184
rect 31987 34153 31999 34156
rect 31941 34147 31999 34153
rect 32030 34144 32036 34156
rect 32088 34144 32094 34196
rect 35253 34187 35311 34193
rect 35253 34153 35265 34187
rect 35299 34184 35311 34187
rect 35526 34184 35532 34196
rect 35299 34156 35532 34184
rect 35299 34153 35311 34156
rect 35253 34147 35311 34153
rect 35526 34144 35532 34156
rect 35584 34144 35590 34196
rect 35894 34184 35900 34196
rect 35855 34156 35900 34184
rect 35894 34144 35900 34156
rect 35952 34184 35958 34196
rect 36909 34187 36967 34193
rect 36909 34184 36921 34187
rect 35952 34156 36921 34184
rect 35952 34144 35958 34156
rect 36909 34153 36921 34156
rect 36955 34153 36967 34187
rect 37550 34184 37556 34196
rect 37511 34156 37556 34184
rect 36909 34147 36967 34153
rect 37550 34144 37556 34156
rect 37608 34144 37614 34196
rect 38286 34184 38292 34196
rect 38247 34156 38292 34184
rect 38286 34144 38292 34156
rect 38344 34144 38350 34196
rect 15286 34076 15292 34128
rect 15344 34116 15350 34128
rect 15473 34119 15531 34125
rect 15473 34116 15485 34119
rect 15344 34088 15485 34116
rect 15344 34076 15350 34088
rect 15473 34085 15485 34088
rect 15519 34085 15531 34119
rect 15473 34079 15531 34085
rect 16945 34119 17003 34125
rect 16945 34085 16957 34119
rect 16991 34085 17003 34119
rect 16945 34079 17003 34085
rect 15488 34048 15516 34079
rect 16485 34051 16543 34057
rect 16485 34048 16497 34051
rect 15488 34020 16497 34048
rect 16485 34017 16497 34020
rect 16531 34017 16543 34051
rect 16485 34011 16543 34017
rect 14090 33980 14096 33992
rect 14051 33952 14096 33980
rect 14090 33940 14096 33952
rect 14148 33940 14154 33992
rect 14366 33989 14372 33992
rect 14360 33980 14372 33989
rect 14327 33952 14372 33980
rect 14360 33943 14372 33952
rect 14366 33940 14372 33943
rect 14424 33940 14430 33992
rect 16577 33983 16635 33989
rect 16577 33949 16589 33983
rect 16623 33949 16635 33983
rect 16960 33980 16988 34079
rect 18138 34076 18144 34128
rect 18196 34116 18202 34128
rect 18601 34119 18659 34125
rect 18601 34116 18613 34119
rect 18196 34088 18613 34116
rect 18196 34076 18202 34088
rect 18601 34085 18613 34088
rect 18647 34085 18659 34119
rect 18601 34079 18659 34085
rect 20070 34076 20076 34128
rect 20128 34116 20134 34128
rect 20622 34116 20628 34128
rect 20128 34088 20628 34116
rect 20128 34076 20134 34088
rect 20622 34076 20628 34088
rect 20680 34116 20686 34128
rect 20717 34119 20775 34125
rect 20717 34116 20729 34119
rect 20680 34088 20729 34116
rect 20680 34076 20686 34088
rect 20717 34085 20729 34088
rect 20763 34085 20775 34119
rect 20717 34079 20775 34085
rect 27341 34119 27399 34125
rect 27341 34085 27353 34119
rect 27387 34085 27399 34119
rect 27341 34079 27399 34085
rect 18141 33983 18199 33989
rect 18141 33980 18153 33983
rect 16960 33952 18153 33980
rect 16577 33943 16635 33949
rect 18141 33949 18153 33952
rect 18187 33949 18199 33983
rect 18322 33980 18328 33992
rect 18283 33952 18328 33980
rect 18141 33943 18199 33949
rect 16592 33912 16620 33943
rect 18322 33940 18328 33952
rect 18380 33940 18386 33992
rect 18417 33983 18475 33989
rect 18417 33949 18429 33983
rect 18463 33949 18475 33983
rect 18690 33980 18696 33992
rect 18651 33952 18696 33980
rect 18417 33943 18475 33949
rect 18230 33912 18236 33924
rect 16592 33884 18236 33912
rect 18230 33872 18236 33884
rect 18288 33872 18294 33924
rect 18432 33912 18460 33943
rect 18690 33940 18696 33952
rect 18748 33980 18754 33992
rect 19426 33980 19432 33992
rect 18748 33952 19432 33980
rect 18748 33940 18754 33952
rect 19426 33940 19432 33952
rect 19484 33940 19490 33992
rect 20070 33980 20076 33992
rect 20031 33952 20076 33980
rect 20070 33940 20076 33952
rect 20128 33940 20134 33992
rect 21082 33940 21088 33992
rect 21140 33980 21146 33992
rect 21830 33983 21888 33989
rect 21830 33980 21842 33983
rect 21140 33952 21842 33980
rect 21140 33940 21146 33952
rect 21830 33949 21842 33952
rect 21876 33949 21888 33983
rect 21830 33943 21888 33949
rect 22097 33983 22155 33989
rect 22097 33949 22109 33983
rect 22143 33980 22155 33983
rect 22646 33980 22652 33992
rect 22143 33952 22652 33980
rect 22143 33949 22155 33952
rect 22097 33943 22155 33949
rect 22646 33940 22652 33952
rect 22704 33940 22710 33992
rect 26142 33940 26148 33992
rect 26200 33980 26206 33992
rect 26329 33983 26387 33989
rect 26329 33980 26341 33983
rect 26200 33952 26341 33980
rect 26200 33940 26206 33952
rect 26329 33949 26341 33952
rect 26375 33949 26387 33983
rect 26510 33980 26516 33992
rect 26471 33952 26516 33980
rect 26329 33943 26387 33949
rect 26510 33940 26516 33952
rect 26568 33940 26574 33992
rect 27356 33980 27384 34079
rect 35342 34076 35348 34128
rect 35400 34116 35406 34128
rect 38838 34116 38844 34128
rect 35400 34088 37136 34116
rect 38799 34088 38844 34116
rect 35400 34076 35406 34088
rect 30282 34048 30288 34060
rect 30243 34020 30288 34048
rect 30282 34008 30288 34020
rect 30340 34008 30346 34060
rect 35161 34051 35219 34057
rect 35161 34017 35173 34051
rect 35207 34048 35219 34051
rect 35618 34048 35624 34060
rect 35207 34020 35624 34048
rect 35207 34017 35219 34020
rect 35161 34011 35219 34017
rect 35618 34008 35624 34020
rect 35676 34008 35682 34060
rect 36262 34048 36268 34060
rect 36004 34020 36268 34048
rect 27801 33983 27859 33989
rect 27801 33980 27813 33983
rect 27356 33952 27813 33980
rect 27801 33949 27813 33952
rect 27847 33949 27859 33983
rect 30006 33980 30012 33992
rect 29967 33952 30012 33980
rect 27801 33943 27859 33949
rect 30006 33940 30012 33952
rect 30064 33940 30070 33992
rect 33321 33983 33379 33989
rect 33321 33949 33333 33983
rect 33367 33980 33379 33983
rect 33870 33980 33876 33992
rect 33367 33952 33876 33980
rect 33367 33949 33379 33952
rect 33321 33943 33379 33949
rect 33870 33940 33876 33952
rect 33928 33940 33934 33992
rect 35345 33983 35403 33989
rect 35345 33949 35357 33983
rect 35391 33949 35403 33983
rect 35345 33943 35403 33949
rect 35437 33983 35495 33989
rect 35437 33949 35449 33983
rect 35483 33980 35495 33983
rect 36004 33980 36032 34020
rect 36262 34008 36268 34020
rect 36320 34008 36326 34060
rect 37108 34057 37136 34088
rect 38838 34076 38844 34088
rect 38896 34076 38902 34128
rect 37093 34051 37151 34057
rect 37093 34017 37105 34051
rect 37139 34048 37151 34051
rect 37182 34048 37188 34060
rect 37139 34020 37188 34048
rect 37139 34017 37151 34020
rect 37093 34011 37151 34017
rect 37182 34008 37188 34020
rect 37240 34008 37246 34060
rect 38930 34008 38936 34060
rect 38988 34048 38994 34060
rect 39850 34048 39856 34060
rect 38988 34020 39856 34048
rect 38988 34008 38994 34020
rect 39850 34008 39856 34020
rect 39908 34008 39914 34060
rect 35483 33952 36032 33980
rect 36081 33983 36139 33989
rect 35483 33949 35495 33952
rect 35437 33943 35495 33949
rect 36081 33949 36093 33983
rect 36127 33949 36139 33983
rect 36814 33980 36820 33992
rect 36775 33952 36820 33980
rect 36081 33943 36139 33949
rect 18782 33912 18788 33924
rect 18432 33884 18788 33912
rect 18782 33872 18788 33884
rect 18840 33912 18846 33924
rect 19978 33912 19984 33924
rect 18840 33884 19984 33912
rect 18840 33872 18846 33884
rect 19978 33872 19984 33884
rect 20036 33872 20042 33924
rect 22186 33872 22192 33924
rect 22244 33912 22250 33924
rect 26973 33915 27031 33921
rect 26973 33912 26985 33915
rect 22244 33884 26985 33912
rect 22244 33872 22250 33884
rect 26973 33881 26985 33884
rect 27019 33912 27031 33915
rect 28442 33912 28448 33924
rect 27019 33884 28448 33912
rect 27019 33881 27031 33884
rect 26973 33875 27031 33881
rect 28442 33872 28448 33884
rect 28500 33912 28506 33924
rect 28994 33912 29000 33924
rect 28500 33884 29000 33912
rect 28500 33872 28506 33884
rect 28994 33872 29000 33884
rect 29052 33872 29058 33924
rect 33076 33915 33134 33921
rect 33076 33881 33088 33915
rect 33122 33912 33134 33915
rect 33962 33912 33968 33924
rect 33122 33884 33968 33912
rect 33122 33881 33134 33884
rect 33076 33875 33134 33881
rect 33962 33872 33968 33884
rect 34020 33872 34026 33924
rect 35360 33912 35388 33943
rect 36096 33912 36124 33943
rect 36814 33940 36820 33952
rect 36872 33940 36878 33992
rect 37553 33983 37611 33989
rect 37553 33980 37565 33983
rect 37108 33952 37565 33980
rect 37108 33921 37136 33952
rect 37553 33949 37565 33952
rect 37599 33949 37611 33983
rect 37553 33943 37611 33949
rect 37737 33983 37795 33989
rect 37737 33949 37749 33983
rect 37783 33980 37795 33983
rect 38010 33980 38016 33992
rect 37783 33952 38016 33980
rect 37783 33949 37795 33952
rect 37737 33943 37795 33949
rect 38010 33940 38016 33952
rect 38068 33940 38074 33992
rect 38654 33980 38660 33992
rect 38615 33952 38660 33980
rect 38654 33940 38660 33952
rect 38712 33940 38718 33992
rect 40126 33989 40132 33992
rect 40120 33980 40132 33989
rect 40087 33952 40132 33980
rect 40120 33943 40132 33952
rect 40126 33940 40132 33943
rect 40184 33940 40190 33992
rect 41598 33940 41604 33992
rect 41656 33980 41662 33992
rect 41693 33983 41751 33989
rect 41693 33980 41705 33983
rect 41656 33952 41705 33980
rect 41656 33940 41662 33952
rect 41693 33949 41705 33952
rect 41739 33949 41751 33983
rect 41693 33943 41751 33949
rect 35360 33884 36124 33912
rect 26513 33847 26571 33853
rect 26513 33813 26525 33847
rect 26559 33844 26571 33847
rect 27173 33847 27231 33853
rect 27173 33844 27185 33847
rect 26559 33816 27185 33844
rect 26559 33813 26571 33816
rect 26513 33807 26571 33813
rect 27173 33813 27185 33816
rect 27219 33813 27231 33847
rect 27982 33844 27988 33856
rect 27943 33816 27988 33844
rect 27173 33807 27231 33813
rect 27982 33804 27988 33816
rect 28040 33804 28046 33856
rect 36096 33844 36124 33884
rect 37093 33915 37151 33921
rect 37093 33881 37105 33915
rect 37139 33881 37151 33915
rect 37093 33875 37151 33881
rect 38565 33915 38623 33921
rect 38565 33881 38577 33915
rect 38611 33912 38623 33915
rect 38746 33912 38752 33924
rect 38611 33884 38752 33912
rect 38611 33881 38623 33884
rect 38565 33875 38623 33881
rect 38746 33872 38752 33884
rect 38804 33912 38810 33924
rect 38804 33884 41276 33912
rect 38804 33872 38810 33884
rect 38470 33844 38476 33856
rect 36096 33816 38476 33844
rect 38470 33804 38476 33816
rect 38528 33804 38534 33856
rect 41248 33853 41276 33884
rect 41233 33847 41291 33853
rect 41233 33813 41245 33847
rect 41279 33813 41291 33847
rect 41233 33807 41291 33813
rect 41690 33804 41696 33856
rect 41748 33844 41754 33856
rect 41785 33847 41843 33853
rect 41785 33844 41797 33847
rect 41748 33816 41797 33844
rect 41748 33804 41754 33816
rect 41785 33813 41797 33816
rect 41831 33813 41843 33847
rect 41785 33807 41843 33813
rect 1104 33754 42872 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 42872 33754
rect 1104 33680 42872 33702
rect 16666 33600 16672 33652
rect 16724 33640 16730 33652
rect 16761 33643 16819 33649
rect 16761 33640 16773 33643
rect 16724 33612 16773 33640
rect 16724 33600 16730 33612
rect 16761 33609 16773 33612
rect 16807 33609 16819 33643
rect 19058 33640 19064 33652
rect 16761 33603 16819 33609
rect 18984 33612 19064 33640
rect 18984 33581 19012 33612
rect 19058 33600 19064 33612
rect 19116 33640 19122 33652
rect 19116 33612 19932 33640
rect 19116 33600 19122 33612
rect 18969 33575 19027 33581
rect 18969 33541 18981 33575
rect 19015 33541 19027 33575
rect 18969 33535 19027 33541
rect 19150 33532 19156 33584
rect 19208 33581 19214 33584
rect 19904 33581 19932 33612
rect 20898 33600 20904 33652
rect 20956 33640 20962 33652
rect 21821 33643 21879 33649
rect 21821 33640 21833 33643
rect 20956 33612 21833 33640
rect 20956 33600 20962 33612
rect 21821 33609 21833 33612
rect 21867 33609 21879 33643
rect 25958 33640 25964 33652
rect 21821 33603 21879 33609
rect 24964 33612 25964 33640
rect 19208 33575 19237 33581
rect 19225 33541 19237 33575
rect 19208 33535 19237 33541
rect 19889 33575 19947 33581
rect 19889 33541 19901 33575
rect 19935 33541 19947 33575
rect 19889 33535 19947 33541
rect 19208 33532 19214 33535
rect 20622 33532 20628 33584
rect 20680 33572 20686 33584
rect 20993 33575 21051 33581
rect 20993 33572 21005 33575
rect 20680 33544 21005 33572
rect 20680 33532 20686 33544
rect 20993 33541 21005 33544
rect 21039 33541 21051 33575
rect 20993 33535 21051 33541
rect 21266 33532 21272 33584
rect 21324 33572 21330 33584
rect 21973 33575 22031 33581
rect 21973 33572 21985 33575
rect 21324 33544 21985 33572
rect 21324 33532 21330 33544
rect 21973 33541 21985 33544
rect 22019 33541 22031 33575
rect 22186 33572 22192 33584
rect 22147 33544 22192 33572
rect 21973 33535 22031 33541
rect 22186 33532 22192 33544
rect 22244 33532 22250 33584
rect 16850 33504 16856 33516
rect 16811 33476 16856 33504
rect 16850 33464 16856 33476
rect 16908 33464 16914 33516
rect 18874 33504 18880 33516
rect 18835 33476 18880 33504
rect 18874 33464 18880 33476
rect 18932 33464 18938 33516
rect 19058 33464 19064 33516
rect 19116 33504 19122 33516
rect 20717 33507 20775 33513
rect 19116 33476 19161 33504
rect 19116 33464 19122 33476
rect 20717 33473 20729 33507
rect 20763 33504 20775 33507
rect 20806 33504 20812 33516
rect 20763 33476 20812 33504
rect 20763 33473 20775 33476
rect 20717 33467 20775 33473
rect 20806 33464 20812 33476
rect 20864 33464 20870 33516
rect 20901 33507 20959 33513
rect 20901 33473 20913 33507
rect 20947 33473 20959 33507
rect 21085 33507 21143 33513
rect 21085 33504 21097 33507
rect 20901 33467 20959 33473
rect 21008 33476 21097 33504
rect 19337 33439 19395 33445
rect 19337 33405 19349 33439
rect 19383 33436 19395 33439
rect 19978 33436 19984 33448
rect 19383 33408 19984 33436
rect 19383 33405 19395 33408
rect 19337 33399 19395 33405
rect 19978 33396 19984 33408
rect 20036 33396 20042 33448
rect 20530 33396 20536 33448
rect 20588 33436 20594 33448
rect 20916 33436 20944 33467
rect 20588 33408 20944 33436
rect 21008 33436 21036 33476
rect 21085 33473 21097 33476
rect 21131 33473 21143 33507
rect 23014 33504 23020 33516
rect 22975 33476 23020 33504
rect 21085 33467 21143 33473
rect 23014 33464 23020 33476
rect 23072 33464 23078 33516
rect 23842 33504 23848 33516
rect 23803 33476 23848 33504
rect 23842 33464 23848 33476
rect 23900 33464 23906 33516
rect 24964 33513 24992 33612
rect 24949 33507 25007 33513
rect 24949 33473 24961 33507
rect 24995 33504 25007 33507
rect 25038 33504 25044 33516
rect 24995 33476 25044 33504
rect 24995 33473 25007 33476
rect 24949 33467 25007 33473
rect 25038 33464 25044 33476
rect 25096 33464 25102 33516
rect 25130 33464 25136 33516
rect 25188 33504 25194 33516
rect 25792 33513 25820 33612
rect 25958 33600 25964 33612
rect 26016 33600 26022 33652
rect 27062 33600 27068 33652
rect 27120 33640 27126 33652
rect 27522 33640 27528 33652
rect 27120 33612 27528 33640
rect 27120 33600 27126 33612
rect 27522 33600 27528 33612
rect 27580 33600 27586 33652
rect 27982 33532 27988 33584
rect 28040 33572 28046 33584
rect 28638 33575 28696 33581
rect 28638 33572 28650 33575
rect 28040 33544 28650 33572
rect 28040 33532 28046 33544
rect 28638 33541 28650 33544
rect 28684 33541 28696 33575
rect 28638 33535 28696 33541
rect 32030 33532 32036 33584
rect 32088 33572 32094 33584
rect 33229 33575 33287 33581
rect 32088 33544 32536 33572
rect 32088 33532 32094 33544
rect 25593 33507 25651 33513
rect 25593 33504 25605 33507
rect 25188 33476 25605 33504
rect 25188 33464 25194 33476
rect 25593 33473 25605 33476
rect 25639 33473 25651 33507
rect 25593 33467 25651 33473
rect 25777 33507 25835 33513
rect 25777 33473 25789 33507
rect 25823 33473 25835 33507
rect 25777 33467 25835 33473
rect 26237 33507 26295 33513
rect 26237 33473 26249 33507
rect 26283 33473 26295 33507
rect 26237 33467 26295 33473
rect 26421 33507 26479 33513
rect 26421 33473 26433 33507
rect 26467 33504 26479 33507
rect 26510 33504 26516 33516
rect 26467 33476 26516 33504
rect 26467 33473 26479 33476
rect 26421 33467 26479 33473
rect 24854 33436 24860 33448
rect 21008 33408 24860 33436
rect 20588 33396 20594 33408
rect 17402 33328 17408 33380
rect 17460 33368 17466 33380
rect 19150 33368 19156 33380
rect 17460 33340 19156 33368
rect 17460 33328 17466 33340
rect 19150 33328 19156 33340
rect 19208 33368 19214 33380
rect 21008 33368 21036 33408
rect 24854 33396 24860 33408
rect 24912 33396 24918 33448
rect 26142 33436 26148 33448
rect 25700 33408 26148 33436
rect 19208 33340 21036 33368
rect 21269 33371 21327 33377
rect 19208 33328 19214 33340
rect 21269 33337 21281 33371
rect 21315 33368 21327 33371
rect 21315 33340 22048 33368
rect 21315 33337 21327 33340
rect 21269 33331 21327 33337
rect 17954 33260 17960 33312
rect 18012 33300 18018 33312
rect 18693 33303 18751 33309
rect 18693 33300 18705 33303
rect 18012 33272 18705 33300
rect 18012 33260 18018 33272
rect 18693 33269 18705 33272
rect 18739 33269 18751 33303
rect 18693 33263 18751 33269
rect 19981 33303 20039 33309
rect 19981 33269 19993 33303
rect 20027 33300 20039 33303
rect 20530 33300 20536 33312
rect 20027 33272 20536 33300
rect 20027 33269 20039 33272
rect 19981 33263 20039 33269
rect 20530 33260 20536 33272
rect 20588 33260 20594 33312
rect 22020 33309 22048 33340
rect 25700 33312 25728 33408
rect 26142 33396 26148 33408
rect 26200 33436 26206 33448
rect 26252 33436 26280 33467
rect 26510 33464 26516 33476
rect 26568 33464 26574 33516
rect 28902 33504 28908 33516
rect 28863 33476 28908 33504
rect 28902 33464 28908 33476
rect 28960 33464 28966 33516
rect 32309 33507 32367 33513
rect 32309 33473 32321 33507
rect 32355 33504 32367 33507
rect 32398 33504 32404 33516
rect 32355 33476 32404 33504
rect 32355 33473 32367 33476
rect 32309 33467 32367 33473
rect 32398 33464 32404 33476
rect 32456 33464 32462 33516
rect 32508 33513 32536 33544
rect 33229 33541 33241 33575
rect 33275 33572 33287 33575
rect 35342 33572 35348 33584
rect 33275 33544 35348 33572
rect 33275 33541 33287 33544
rect 33229 33535 33287 33541
rect 35342 33532 35348 33544
rect 35400 33532 35406 33584
rect 39022 33532 39028 33584
rect 39080 33572 39086 33584
rect 39209 33575 39267 33581
rect 39209 33572 39221 33575
rect 39080 33544 39221 33572
rect 39080 33532 39086 33544
rect 39209 33541 39221 33544
rect 39255 33541 39267 33575
rect 41690 33572 41696 33584
rect 41651 33544 41696 33572
rect 39209 33535 39267 33541
rect 41690 33532 41696 33544
rect 41748 33532 41754 33584
rect 32493 33507 32551 33513
rect 32493 33473 32505 33507
rect 32539 33473 32551 33507
rect 32493 33467 32551 33473
rect 32674 33464 32680 33516
rect 32732 33504 32738 33516
rect 33045 33507 33103 33513
rect 33045 33504 33057 33507
rect 32732 33476 33057 33504
rect 32732 33464 32738 33476
rect 33045 33473 33057 33476
rect 33091 33473 33103 33507
rect 33045 33467 33103 33473
rect 38197 33507 38255 33513
rect 38197 33473 38209 33507
rect 38243 33504 38255 33507
rect 38930 33504 38936 33516
rect 38243 33476 38936 33504
rect 38243 33473 38255 33476
rect 38197 33467 38255 33473
rect 38930 33464 38936 33476
rect 38988 33464 38994 33516
rect 41877 33507 41935 33513
rect 41877 33473 41889 33507
rect 41923 33504 41935 33507
rect 41966 33504 41972 33516
rect 41923 33476 41972 33504
rect 41923 33473 41935 33476
rect 41877 33467 41935 33473
rect 41966 33464 41972 33476
rect 42024 33464 42030 33516
rect 38378 33436 38384 33448
rect 26200 33408 26280 33436
rect 38339 33408 38384 33436
rect 26200 33396 26206 33408
rect 38378 33396 38384 33408
rect 38436 33396 38442 33448
rect 41322 33436 41328 33448
rect 41283 33408 41328 33436
rect 41322 33396 41328 33408
rect 41380 33396 41386 33448
rect 32401 33371 32459 33377
rect 32401 33337 32413 33371
rect 32447 33368 32459 33371
rect 33226 33368 33232 33380
rect 32447 33340 33232 33368
rect 32447 33337 32459 33340
rect 32401 33331 32459 33337
rect 33226 33328 33232 33340
rect 33284 33328 33290 33380
rect 38470 33328 38476 33380
rect 38528 33368 38534 33380
rect 38841 33371 38899 33377
rect 38841 33368 38853 33371
rect 38528 33340 38853 33368
rect 38528 33328 38534 33340
rect 38841 33337 38853 33340
rect 38887 33337 38899 33371
rect 38841 33331 38899 33337
rect 22005 33303 22063 33309
rect 22005 33269 22017 33303
rect 22051 33269 22063 33303
rect 22005 33263 22063 33269
rect 22646 33260 22652 33312
rect 22704 33300 22710 33312
rect 23109 33303 23167 33309
rect 23109 33300 23121 33303
rect 22704 33272 23121 33300
rect 22704 33260 22710 33272
rect 23109 33269 23121 33272
rect 23155 33269 23167 33303
rect 23658 33300 23664 33312
rect 23619 33272 23664 33300
rect 23109 33263 23167 33269
rect 23658 33260 23664 33272
rect 23716 33260 23722 33312
rect 24762 33300 24768 33312
rect 24723 33272 24768 33300
rect 24762 33260 24768 33272
rect 24820 33260 24826 33312
rect 25682 33300 25688 33312
rect 25643 33272 25688 33300
rect 25682 33260 25688 33272
rect 25740 33260 25746 33312
rect 26237 33303 26295 33309
rect 26237 33269 26249 33303
rect 26283 33300 26295 33303
rect 26326 33300 26332 33312
rect 26283 33272 26332 33300
rect 26283 33269 26295 33272
rect 26237 33263 26295 33269
rect 26326 33260 26332 33272
rect 26384 33260 26390 33312
rect 38013 33303 38071 33309
rect 38013 33269 38025 33303
rect 38059 33300 38071 33303
rect 38286 33300 38292 33312
rect 38059 33272 38292 33300
rect 38059 33269 38071 33272
rect 38013 33263 38071 33269
rect 38286 33260 38292 33272
rect 38344 33260 38350 33312
rect 39209 33303 39267 33309
rect 39209 33269 39221 33303
rect 39255 33300 39267 33303
rect 39298 33300 39304 33312
rect 39255 33272 39304 33300
rect 39255 33269 39267 33272
rect 39209 33263 39267 33269
rect 39298 33260 39304 33272
rect 39356 33260 39362 33312
rect 39393 33303 39451 33309
rect 39393 33269 39405 33303
rect 39439 33300 39451 33303
rect 39942 33300 39948 33312
rect 39439 33272 39948 33300
rect 39439 33269 39451 33272
rect 39393 33263 39451 33269
rect 39942 33260 39948 33272
rect 40000 33260 40006 33312
rect 1104 33210 42872 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 42872 33210
rect 1104 33136 42872 33158
rect 18601 33099 18659 33105
rect 18601 33065 18613 33099
rect 18647 33096 18659 33099
rect 18874 33096 18880 33108
rect 18647 33068 18880 33096
rect 18647 33065 18659 33068
rect 18601 33059 18659 33065
rect 18874 33056 18880 33068
rect 18932 33096 18938 33108
rect 18932 33068 20760 33096
rect 18932 33056 18938 33068
rect 19337 33031 19395 33037
rect 19337 32997 19349 33031
rect 19383 33028 19395 33031
rect 20254 33028 20260 33040
rect 19383 33000 20260 33028
rect 19383 32997 19395 33000
rect 19337 32991 19395 32997
rect 20254 32988 20260 33000
rect 20312 32988 20318 33040
rect 18414 32920 18420 32972
rect 18472 32960 18478 32972
rect 19797 32963 19855 32969
rect 18472 32932 19748 32960
rect 18472 32920 18478 32932
rect 15289 32895 15347 32901
rect 15289 32861 15301 32895
rect 15335 32892 15347 32895
rect 16669 32895 16727 32901
rect 16669 32892 16681 32895
rect 15335 32864 16681 32892
rect 15335 32861 15347 32864
rect 15289 32855 15347 32861
rect 16669 32861 16681 32864
rect 16715 32861 16727 32895
rect 16850 32892 16856 32904
rect 16811 32864 16856 32892
rect 16669 32855 16727 32861
rect 16850 32852 16856 32864
rect 16908 32852 16914 32904
rect 17037 32895 17095 32901
rect 17037 32861 17049 32895
rect 17083 32892 17095 32895
rect 17773 32895 17831 32901
rect 17773 32892 17785 32895
rect 17083 32864 17785 32892
rect 17083 32861 17095 32864
rect 17037 32855 17095 32861
rect 17773 32861 17785 32864
rect 17819 32861 17831 32895
rect 17773 32855 17831 32861
rect 17865 32895 17923 32901
rect 17865 32861 17877 32895
rect 17911 32892 17923 32895
rect 17954 32892 17960 32904
rect 17911 32864 17960 32892
rect 17911 32861 17923 32864
rect 17865 32855 17923 32861
rect 17788 32824 17816 32855
rect 17954 32852 17960 32864
rect 18012 32852 18018 32904
rect 18230 32852 18236 32904
rect 18288 32892 18294 32904
rect 18506 32892 18512 32904
rect 18288 32864 18512 32892
rect 18288 32852 18294 32864
rect 18506 32852 18512 32864
rect 18564 32852 18570 32904
rect 18693 32895 18751 32901
rect 18693 32861 18705 32895
rect 18739 32892 18751 32895
rect 18782 32892 18788 32904
rect 18739 32864 18788 32892
rect 18739 32861 18751 32864
rect 18693 32855 18751 32861
rect 18782 32852 18788 32864
rect 18840 32852 18846 32904
rect 19720 32892 19748 32932
rect 19797 32929 19809 32963
rect 19843 32960 19855 32963
rect 20162 32960 20168 32972
rect 19843 32932 20168 32960
rect 19843 32929 19855 32932
rect 19797 32923 19855 32929
rect 20162 32920 20168 32932
rect 20220 32960 20226 32972
rect 20346 32960 20352 32972
rect 20220 32932 20352 32960
rect 20220 32920 20226 32932
rect 20346 32920 20352 32932
rect 20404 32960 20410 32972
rect 20404 32932 20576 32960
rect 20404 32920 20410 32932
rect 20070 32892 20076 32904
rect 19720 32864 20076 32892
rect 20070 32852 20076 32864
rect 20128 32852 20134 32904
rect 20548 32901 20576 32932
rect 20732 32901 20760 33068
rect 20806 33056 20812 33108
rect 20864 33096 20870 33108
rect 21269 33099 21327 33105
rect 21269 33096 21281 33099
rect 20864 33068 21281 33096
rect 20864 33056 20870 33068
rect 21269 33065 21281 33068
rect 21315 33065 21327 33099
rect 21269 33059 21327 33065
rect 24854 33056 24860 33108
rect 24912 33096 24918 33108
rect 26142 33096 26148 33108
rect 24912 33068 26148 33096
rect 24912 33056 24918 33068
rect 26142 33056 26148 33068
rect 26200 33056 26206 33108
rect 26789 33099 26847 33105
rect 26789 33065 26801 33099
rect 26835 33096 26847 33099
rect 27154 33096 27160 33108
rect 26835 33068 27160 33096
rect 26835 33065 26847 33068
rect 26789 33059 26847 33065
rect 27154 33056 27160 33068
rect 27212 33056 27218 33108
rect 29914 33056 29920 33108
rect 29972 33096 29978 33108
rect 30101 33099 30159 33105
rect 30101 33096 30113 33099
rect 29972 33068 30113 33096
rect 29972 33056 29978 33068
rect 30101 33065 30113 33068
rect 30147 33096 30159 33099
rect 32306 33096 32312 33108
rect 30147 33068 31754 33096
rect 32267 33068 32312 33096
rect 30147 33065 30159 33068
rect 30101 33059 30159 33065
rect 23845 33031 23903 33037
rect 23845 32997 23857 33031
rect 23891 33028 23903 33031
rect 25038 33028 25044 33040
rect 23891 33000 25044 33028
rect 23891 32997 23903 33000
rect 23845 32991 23903 32997
rect 25038 32988 25044 33000
rect 25096 32988 25102 33040
rect 30926 33028 30932 33040
rect 30887 33000 30932 33028
rect 30926 32988 30932 33000
rect 30984 32988 30990 33040
rect 31726 33028 31754 33068
rect 32306 33056 32312 33068
rect 32364 33056 32370 33108
rect 33229 33099 33287 33105
rect 33229 33065 33241 33099
rect 33275 33096 33287 33099
rect 33275 33068 38332 33096
rect 33275 33065 33287 33068
rect 33229 33059 33287 33065
rect 32950 33028 32956 33040
rect 31726 33000 32956 33028
rect 32950 32988 32956 33000
rect 33008 32988 33014 33040
rect 38304 33028 38332 33068
rect 38378 33056 38384 33108
rect 38436 33096 38442 33108
rect 38565 33099 38623 33105
rect 38565 33096 38577 33099
rect 38436 33068 38577 33096
rect 38436 33056 38442 33068
rect 38565 33065 38577 33068
rect 38611 33096 38623 33099
rect 39666 33096 39672 33108
rect 38611 33068 39672 33096
rect 38611 33065 38623 33068
rect 38565 33059 38623 33065
rect 39666 33056 39672 33068
rect 39724 33056 39730 33108
rect 39482 33028 39488 33040
rect 38304 33000 39488 33028
rect 39482 32988 39488 33000
rect 39540 32988 39546 33040
rect 25682 32960 25688 32972
rect 24596 32932 25688 32960
rect 20533 32895 20591 32901
rect 20533 32861 20545 32895
rect 20579 32861 20591 32895
rect 20533 32855 20591 32861
rect 20717 32895 20775 32901
rect 20717 32861 20729 32895
rect 20763 32861 20775 32895
rect 20717 32855 20775 32861
rect 21361 32895 21419 32901
rect 21361 32861 21373 32895
rect 21407 32861 21419 32895
rect 21361 32855 21419 32861
rect 22465 32895 22523 32901
rect 22465 32861 22477 32895
rect 22511 32892 22523 32895
rect 22554 32892 22560 32904
rect 22511 32864 22560 32892
rect 22511 32861 22523 32864
rect 22465 32855 22523 32861
rect 18322 32824 18328 32836
rect 17788 32796 18328 32824
rect 18322 32784 18328 32796
rect 18380 32784 18386 32836
rect 19058 32784 19064 32836
rect 19116 32824 19122 32836
rect 19337 32827 19395 32833
rect 19337 32824 19349 32827
rect 19116 32796 19349 32824
rect 19116 32784 19122 32796
rect 19337 32793 19349 32796
rect 19383 32793 19395 32827
rect 19337 32787 19395 32793
rect 20625 32827 20683 32833
rect 20625 32793 20637 32827
rect 20671 32824 20683 32827
rect 20806 32824 20812 32836
rect 20671 32796 20812 32824
rect 20671 32793 20683 32796
rect 20625 32787 20683 32793
rect 20806 32784 20812 32796
rect 20864 32824 20870 32836
rect 21376 32824 21404 32855
rect 22554 32852 22560 32864
rect 22612 32852 22618 32904
rect 22732 32895 22790 32901
rect 22732 32861 22744 32895
rect 22778 32892 22790 32895
rect 23658 32892 23664 32904
rect 22778 32864 23664 32892
rect 22778 32861 22790 32864
rect 22732 32855 22790 32861
rect 23658 32852 23664 32864
rect 23716 32852 23722 32904
rect 24596 32901 24624 32932
rect 25682 32920 25688 32932
rect 25740 32920 25746 32972
rect 27893 32963 27951 32969
rect 27893 32960 27905 32963
rect 27356 32932 27905 32960
rect 24581 32895 24639 32901
rect 24581 32861 24593 32895
rect 24627 32861 24639 32895
rect 24762 32892 24768 32904
rect 24723 32864 24768 32892
rect 24581 32855 24639 32861
rect 24762 32852 24768 32864
rect 24820 32852 24826 32904
rect 24854 32852 24860 32904
rect 24912 32901 24918 32904
rect 24912 32895 24941 32901
rect 24929 32861 24941 32895
rect 25038 32892 25044 32904
rect 24999 32864 25044 32892
rect 24912 32855 24941 32861
rect 24912 32852 24918 32855
rect 25038 32852 25044 32864
rect 25096 32852 25102 32904
rect 25406 32852 25412 32904
rect 25464 32892 25470 32904
rect 25501 32895 25559 32901
rect 25501 32892 25513 32895
rect 25464 32864 25513 32892
rect 25464 32852 25470 32864
rect 25501 32861 25513 32864
rect 25547 32861 25559 32895
rect 25501 32855 25559 32861
rect 25777 32895 25835 32901
rect 25777 32861 25789 32895
rect 25823 32861 25835 32895
rect 25777 32855 25835 32861
rect 20864 32796 21404 32824
rect 24673 32827 24731 32833
rect 20864 32784 20870 32796
rect 24673 32793 24685 32827
rect 24719 32793 24731 32827
rect 24673 32787 24731 32793
rect 15102 32756 15108 32768
rect 15063 32728 15108 32756
rect 15102 32716 15108 32728
rect 15160 32716 15166 32768
rect 18049 32759 18107 32765
rect 18049 32725 18061 32759
rect 18095 32756 18107 32759
rect 18414 32756 18420 32768
rect 18095 32728 18420 32756
rect 18095 32725 18107 32728
rect 18049 32719 18107 32725
rect 18414 32716 18420 32728
rect 18472 32716 18478 32768
rect 18690 32716 18696 32768
rect 18748 32756 18754 32768
rect 19889 32759 19947 32765
rect 19889 32756 19901 32759
rect 18748 32728 19901 32756
rect 18748 32716 18754 32728
rect 19889 32725 19901 32728
rect 19935 32756 19947 32759
rect 19978 32756 19984 32768
rect 19935 32728 19984 32756
rect 19935 32725 19947 32728
rect 19889 32719 19947 32725
rect 19978 32716 19984 32728
rect 20036 32716 20042 32768
rect 24394 32756 24400 32768
rect 24355 32728 24400 32756
rect 24394 32716 24400 32728
rect 24452 32716 24458 32768
rect 24688 32756 24716 32787
rect 25424 32756 25452 32852
rect 25792 32824 25820 32855
rect 26142 32852 26148 32904
rect 26200 32892 26206 32904
rect 26927 32895 26985 32901
rect 26927 32892 26939 32895
rect 26200 32864 26939 32892
rect 26200 32852 26206 32864
rect 26927 32861 26939 32864
rect 26973 32861 26985 32895
rect 27062 32892 27068 32904
rect 27023 32864 27068 32892
rect 26927 32855 26985 32861
rect 27062 32852 27068 32864
rect 27120 32852 27126 32904
rect 27356 32901 27384 32932
rect 27893 32929 27905 32932
rect 27939 32929 27951 32963
rect 32214 32960 32220 32972
rect 32175 32932 32220 32960
rect 27893 32923 27951 32929
rect 32214 32920 32220 32932
rect 32272 32920 32278 32972
rect 34054 32960 34060 32972
rect 32324 32932 34060 32960
rect 27341 32895 27399 32901
rect 27341 32861 27353 32895
rect 27387 32861 27399 32895
rect 27801 32895 27859 32901
rect 27801 32892 27813 32895
rect 27341 32855 27399 32861
rect 27448 32864 27813 32892
rect 26234 32824 26240 32836
rect 25792 32796 26240 32824
rect 26234 32784 26240 32796
rect 26292 32824 26298 32836
rect 27157 32827 27215 32833
rect 27157 32824 27169 32827
rect 26292 32796 27169 32824
rect 26292 32784 26298 32796
rect 27157 32793 27169 32796
rect 27203 32793 27215 32827
rect 27157 32787 27215 32793
rect 24688 32728 25452 32756
rect 26326 32716 26332 32768
rect 26384 32756 26390 32768
rect 27448 32756 27476 32864
rect 27801 32861 27813 32864
rect 27847 32861 27859 32895
rect 29914 32892 29920 32904
rect 29875 32864 29920 32892
rect 27801 32855 27859 32861
rect 29914 32852 29920 32864
rect 29972 32892 29978 32904
rect 30745 32895 30803 32901
rect 30745 32892 30757 32895
rect 29972 32864 30757 32892
rect 29972 32852 29978 32864
rect 30745 32861 30757 32864
rect 30791 32892 30803 32895
rect 31481 32895 31539 32901
rect 31481 32892 31493 32895
rect 30791 32864 31493 32892
rect 30791 32861 30803 32864
rect 30745 32855 30803 32861
rect 31481 32861 31493 32864
rect 31527 32892 31539 32895
rect 32125 32895 32183 32901
rect 31527 32864 31754 32892
rect 31527 32861 31539 32864
rect 31481 32855 31539 32861
rect 26384 32728 27476 32756
rect 26384 32716 26390 32728
rect 31202 32716 31208 32768
rect 31260 32756 31266 32768
rect 31573 32759 31631 32765
rect 31573 32756 31585 32759
rect 31260 32728 31585 32756
rect 31260 32716 31266 32728
rect 31573 32725 31585 32728
rect 31619 32725 31631 32759
rect 31726 32756 31754 32864
rect 32125 32861 32137 32895
rect 32171 32892 32183 32895
rect 32324 32892 32352 32932
rect 34054 32920 34060 32932
rect 34112 32920 34118 32972
rect 34977 32963 35035 32969
rect 34977 32929 34989 32963
rect 35023 32960 35035 32963
rect 35342 32960 35348 32972
rect 35023 32932 35348 32960
rect 35023 32929 35035 32932
rect 34977 32923 35035 32929
rect 35342 32920 35348 32932
rect 35400 32920 35406 32972
rect 37826 32920 37832 32972
rect 37884 32960 37890 32972
rect 38105 32963 38163 32969
rect 38105 32960 38117 32963
rect 37884 32932 38117 32960
rect 37884 32920 37890 32932
rect 38105 32929 38117 32932
rect 38151 32929 38163 32963
rect 38105 32923 38163 32929
rect 32171 32864 32352 32892
rect 32401 32895 32459 32901
rect 32171 32861 32183 32864
rect 32125 32855 32183 32861
rect 32401 32861 32413 32895
rect 32447 32892 32459 32895
rect 32490 32892 32496 32904
rect 32447 32864 32496 32892
rect 32447 32861 32459 32864
rect 32401 32855 32459 32861
rect 32490 32852 32496 32864
rect 32548 32852 32554 32904
rect 33045 32895 33103 32901
rect 33045 32892 33057 32895
rect 32600 32864 33057 32892
rect 32490 32756 32496 32768
rect 31726 32728 32496 32756
rect 31573 32719 31631 32725
rect 32490 32716 32496 32728
rect 32548 32716 32554 32768
rect 32600 32765 32628 32864
rect 33045 32861 33057 32864
rect 33091 32861 33103 32895
rect 33226 32892 33232 32904
rect 33187 32864 33232 32892
rect 33045 32855 33103 32861
rect 33226 32852 33232 32864
rect 33284 32852 33290 32904
rect 34698 32892 34704 32904
rect 34659 32864 34704 32892
rect 34698 32852 34704 32864
rect 34756 32852 34762 32904
rect 34793 32895 34851 32901
rect 34793 32861 34805 32895
rect 34839 32892 34851 32895
rect 35802 32892 35808 32904
rect 34839 32864 35808 32892
rect 34839 32861 34851 32864
rect 34793 32855 34851 32861
rect 32950 32784 32956 32836
rect 33008 32824 33014 32836
rect 33008 32796 34100 32824
rect 33008 32784 33014 32796
rect 32585 32759 32643 32765
rect 32585 32725 32597 32759
rect 32631 32725 32643 32759
rect 33410 32756 33416 32768
rect 33371 32728 33416 32756
rect 32585 32719 32643 32725
rect 33410 32716 33416 32728
rect 33468 32716 33474 32768
rect 34072 32756 34100 32796
rect 34146 32784 34152 32836
rect 34204 32824 34210 32836
rect 34808 32824 34836 32855
rect 35802 32852 35808 32864
rect 35860 32852 35866 32904
rect 36817 32895 36875 32901
rect 36817 32861 36829 32895
rect 36863 32892 36875 32895
rect 36998 32892 37004 32904
rect 36863 32864 37004 32892
rect 36863 32861 36875 32864
rect 36817 32855 36875 32861
rect 36998 32852 37004 32864
rect 37056 32852 37062 32904
rect 38194 32852 38200 32904
rect 38252 32892 38258 32904
rect 38565 32895 38623 32901
rect 38252 32864 38297 32892
rect 38252 32852 38258 32864
rect 38565 32861 38577 32895
rect 38611 32892 38623 32895
rect 38654 32892 38660 32904
rect 38611 32864 38660 32892
rect 38611 32861 38623 32864
rect 38565 32855 38623 32861
rect 38654 32852 38660 32864
rect 38712 32852 38718 32904
rect 40310 32892 40316 32904
rect 40271 32864 40316 32892
rect 40310 32852 40316 32864
rect 40368 32852 40374 32904
rect 36354 32824 36360 32836
rect 34204 32796 34836 32824
rect 34900 32796 36360 32824
rect 34204 32784 34210 32796
rect 34900 32756 34928 32796
rect 36354 32784 36360 32796
rect 36412 32784 36418 32836
rect 36446 32784 36452 32836
rect 36504 32824 36510 32836
rect 36541 32827 36599 32833
rect 36541 32824 36553 32827
rect 36504 32796 36553 32824
rect 36504 32784 36510 32796
rect 36541 32793 36553 32796
rect 36587 32793 36599 32827
rect 36722 32824 36728 32836
rect 36683 32796 36728 32824
rect 36541 32787 36599 32793
rect 36722 32784 36728 32796
rect 36780 32824 36786 32836
rect 37918 32824 37924 32836
rect 36780 32796 37924 32824
rect 36780 32784 36786 32796
rect 37918 32784 37924 32796
rect 37976 32784 37982 32836
rect 40497 32827 40555 32833
rect 40497 32793 40509 32827
rect 40543 32824 40555 32827
rect 41506 32824 41512 32836
rect 40543 32796 41512 32824
rect 40543 32793 40555 32796
rect 40497 32787 40555 32793
rect 41506 32784 41512 32796
rect 41564 32784 41570 32836
rect 42150 32824 42156 32836
rect 42111 32796 42156 32824
rect 42150 32784 42156 32796
rect 42208 32784 42214 32836
rect 34072 32728 34928 32756
rect 34977 32759 35035 32765
rect 34977 32725 34989 32759
rect 35023 32756 35035 32759
rect 35710 32756 35716 32768
rect 35023 32728 35716 32756
rect 35023 32725 35035 32728
rect 34977 32719 35035 32725
rect 35710 32716 35716 32728
rect 35768 32716 35774 32768
rect 36630 32756 36636 32768
rect 36688 32765 36694 32768
rect 36597 32728 36636 32756
rect 36630 32716 36636 32728
rect 36688 32719 36697 32765
rect 38749 32759 38807 32765
rect 38749 32725 38761 32759
rect 38795 32756 38807 32759
rect 39114 32756 39120 32768
rect 38795 32728 39120 32756
rect 38795 32725 38807 32728
rect 38749 32719 38807 32725
rect 36688 32716 36694 32719
rect 39114 32716 39120 32728
rect 39172 32716 39178 32768
rect 1104 32666 42872 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 42872 32666
rect 1104 32592 42872 32614
rect 18601 32555 18659 32561
rect 18601 32521 18613 32555
rect 18647 32552 18659 32555
rect 18782 32552 18788 32564
rect 18647 32524 18788 32552
rect 18647 32521 18659 32524
rect 18601 32515 18659 32521
rect 18782 32512 18788 32524
rect 18840 32512 18846 32564
rect 19058 32552 19064 32564
rect 19019 32524 19064 32552
rect 19058 32512 19064 32524
rect 19116 32512 19122 32564
rect 20349 32555 20407 32561
rect 20349 32521 20361 32555
rect 20395 32552 20407 32555
rect 21266 32552 21272 32564
rect 20395 32524 21272 32552
rect 20395 32521 20407 32524
rect 20349 32515 20407 32521
rect 21266 32512 21272 32524
rect 21324 32512 21330 32564
rect 23385 32555 23443 32561
rect 23385 32521 23397 32555
rect 23431 32552 23443 32555
rect 23842 32552 23848 32564
rect 23431 32524 23848 32552
rect 23431 32521 23443 32524
rect 23385 32515 23443 32521
rect 23842 32512 23848 32524
rect 23900 32512 23906 32564
rect 24946 32512 24952 32564
rect 25004 32552 25010 32564
rect 26237 32555 26295 32561
rect 26237 32552 26249 32555
rect 25004 32524 26249 32552
rect 25004 32512 25010 32524
rect 26237 32521 26249 32524
rect 26283 32521 26295 32555
rect 26237 32515 26295 32521
rect 26418 32512 26424 32564
rect 26476 32552 26482 32564
rect 26970 32552 26976 32564
rect 26476 32524 26976 32552
rect 26476 32512 26482 32524
rect 26970 32512 26976 32524
rect 27028 32552 27034 32564
rect 27065 32555 27123 32561
rect 27065 32552 27077 32555
rect 27028 32524 27077 32552
rect 27028 32512 27034 32524
rect 27065 32521 27077 32524
rect 27111 32521 27123 32555
rect 27065 32515 27123 32521
rect 28905 32555 28963 32561
rect 28905 32521 28917 32555
rect 28951 32552 28963 32555
rect 29914 32552 29920 32564
rect 28951 32524 29920 32552
rect 28951 32521 28963 32524
rect 28905 32515 28963 32521
rect 29914 32512 29920 32524
rect 29972 32512 29978 32564
rect 30926 32512 30932 32564
rect 30984 32552 30990 32564
rect 34422 32552 34428 32564
rect 30984 32524 34428 32552
rect 30984 32512 30990 32524
rect 34422 32512 34428 32524
rect 34480 32512 34486 32564
rect 34698 32512 34704 32564
rect 34756 32552 34762 32564
rect 35897 32555 35955 32561
rect 35897 32552 35909 32555
rect 34756 32524 35909 32552
rect 34756 32512 34762 32524
rect 35897 32521 35909 32524
rect 35943 32521 35955 32555
rect 36446 32552 36452 32564
rect 36407 32524 36452 32552
rect 35897 32515 35955 32521
rect 36446 32512 36452 32524
rect 36504 32512 36510 32564
rect 36630 32512 36636 32564
rect 36688 32552 36694 32564
rect 38654 32552 38660 32564
rect 36688 32524 37412 32552
rect 38615 32524 38660 32552
rect 36688 32512 36694 32524
rect 14476 32456 17264 32484
rect 14090 32376 14096 32428
rect 14148 32416 14154 32428
rect 14476 32425 14504 32456
rect 14461 32419 14519 32425
rect 14461 32416 14473 32419
rect 14148 32388 14473 32416
rect 14148 32376 14154 32388
rect 14461 32385 14473 32388
rect 14507 32385 14519 32419
rect 14461 32379 14519 32385
rect 14728 32419 14786 32425
rect 14728 32385 14740 32419
rect 14774 32416 14786 32419
rect 15102 32416 15108 32428
rect 14774 32388 15108 32416
rect 14774 32385 14786 32388
rect 14728 32379 14786 32385
rect 15102 32376 15108 32388
rect 15160 32376 15166 32428
rect 17236 32357 17264 32456
rect 17488 32419 17546 32425
rect 17488 32385 17500 32419
rect 17534 32416 17546 32419
rect 18230 32416 18236 32428
rect 17534 32388 18236 32416
rect 17534 32385 17546 32388
rect 17488 32379 17546 32385
rect 18230 32376 18236 32388
rect 18288 32376 18294 32428
rect 18800 32416 18828 32512
rect 18874 32444 18880 32496
rect 18932 32484 18938 32496
rect 21177 32487 21235 32493
rect 18932 32456 20208 32484
rect 18932 32444 18938 32456
rect 19245 32419 19303 32425
rect 19245 32416 19257 32419
rect 18800 32388 19257 32416
rect 19245 32385 19257 32388
rect 19291 32385 19303 32419
rect 19245 32379 19303 32385
rect 19334 32376 19340 32428
rect 19392 32416 19398 32428
rect 20180 32425 20208 32456
rect 21177 32453 21189 32487
rect 21223 32484 21235 32487
rect 22554 32484 22560 32496
rect 21223 32456 22560 32484
rect 21223 32453 21235 32456
rect 21177 32447 21235 32453
rect 22554 32444 22560 32456
rect 22612 32484 22618 32496
rect 23014 32484 23020 32496
rect 22612 32456 23020 32484
rect 22612 32444 22618 32456
rect 23014 32444 23020 32456
rect 23072 32444 23078 32496
rect 24394 32484 24400 32496
rect 23216 32456 24400 32484
rect 19429 32419 19487 32425
rect 19429 32416 19441 32419
rect 19392 32388 19441 32416
rect 19392 32376 19398 32388
rect 19429 32385 19441 32388
rect 19475 32385 19487 32419
rect 19429 32379 19487 32385
rect 20165 32419 20223 32425
rect 20165 32385 20177 32419
rect 20211 32385 20223 32419
rect 20346 32416 20352 32428
rect 20307 32388 20352 32416
rect 20165 32379 20223 32385
rect 20346 32376 20352 32388
rect 20404 32376 20410 32428
rect 23216 32425 23244 32456
rect 24394 32444 24400 32456
rect 24452 32444 24458 32496
rect 33410 32484 33416 32496
rect 25332 32456 33416 32484
rect 23201 32419 23259 32425
rect 23201 32385 23213 32419
rect 23247 32385 23259 32419
rect 23934 32416 23940 32428
rect 23895 32388 23940 32416
rect 23201 32379 23259 32385
rect 23934 32376 23940 32388
rect 23992 32376 23998 32428
rect 24210 32416 24216 32428
rect 24171 32388 24216 32416
rect 24210 32376 24216 32388
rect 24268 32376 24274 32428
rect 24946 32416 24952 32428
rect 24907 32388 24952 32416
rect 24946 32376 24952 32388
rect 25004 32376 25010 32428
rect 25332 32425 25360 32456
rect 25317 32419 25375 32425
rect 25317 32385 25329 32419
rect 25363 32385 25375 32419
rect 25317 32379 25375 32385
rect 25777 32419 25835 32425
rect 25777 32385 25789 32419
rect 25823 32385 25835 32419
rect 25777 32379 25835 32385
rect 26053 32419 26111 32425
rect 26053 32385 26065 32419
rect 26099 32416 26111 32419
rect 27154 32416 27160 32428
rect 26099 32388 27160 32416
rect 26099 32385 26111 32388
rect 26053 32379 26111 32385
rect 17221 32351 17279 32357
rect 17221 32317 17233 32351
rect 17267 32317 17279 32351
rect 17221 32311 17279 32317
rect 15838 32212 15844 32224
rect 15799 32184 15844 32212
rect 15838 32172 15844 32184
rect 15896 32172 15902 32224
rect 17236 32212 17264 32311
rect 18322 32308 18328 32360
rect 18380 32348 18386 32360
rect 23017 32351 23075 32357
rect 23017 32348 23029 32351
rect 18380 32320 23029 32348
rect 18380 32308 18386 32320
rect 23017 32317 23029 32320
rect 23063 32348 23075 32351
rect 23750 32348 23756 32360
rect 23063 32320 23756 32348
rect 23063 32317 23075 32320
rect 23017 32311 23075 32317
rect 23750 32308 23756 32320
rect 23808 32308 23814 32360
rect 24762 32308 24768 32360
rect 24820 32348 24826 32360
rect 25792 32348 25820 32379
rect 27154 32376 27160 32388
rect 27212 32376 27218 32428
rect 28626 32416 28632 32428
rect 28587 32388 28632 32416
rect 28626 32376 28632 32388
rect 28684 32376 28690 32428
rect 28736 32425 28764 32456
rect 33410 32444 33416 32456
rect 33468 32444 33474 32496
rect 34514 32444 34520 32496
rect 34572 32484 34578 32496
rect 37384 32484 37412 32524
rect 38654 32512 38660 32524
rect 38712 32512 38718 32564
rect 39482 32552 39488 32564
rect 39443 32524 39488 32552
rect 39482 32512 39488 32524
rect 39540 32512 39546 32564
rect 37522 32487 37580 32493
rect 37522 32484 37534 32487
rect 34572 32456 37320 32484
rect 37384 32456 37534 32484
rect 34572 32444 34578 32456
rect 28721 32419 28779 32425
rect 28721 32385 28733 32419
rect 28767 32385 28779 32419
rect 28721 32379 28779 32385
rect 28902 32376 28908 32428
rect 28960 32416 28966 32428
rect 29638 32425 29644 32428
rect 29365 32419 29423 32425
rect 29365 32416 29377 32419
rect 28960 32388 29377 32416
rect 28960 32376 28966 32388
rect 29365 32385 29377 32388
rect 29411 32385 29423 32419
rect 29365 32379 29423 32385
rect 29632 32379 29644 32425
rect 29696 32416 29702 32428
rect 29696 32388 29732 32416
rect 29638 32376 29644 32379
rect 29696 32376 29702 32388
rect 31110 32376 31116 32428
rect 31168 32416 31174 32428
rect 31481 32419 31539 32425
rect 31481 32416 31493 32419
rect 31168 32388 31493 32416
rect 31168 32376 31174 32388
rect 31481 32385 31493 32388
rect 31527 32416 31539 32419
rect 32306 32416 32312 32428
rect 31527 32388 32312 32416
rect 31527 32385 31539 32388
rect 31481 32379 31539 32385
rect 32306 32376 32312 32388
rect 32364 32376 32370 32428
rect 32674 32416 32680 32428
rect 32635 32388 32680 32416
rect 32674 32376 32680 32388
rect 32732 32376 32738 32428
rect 34140 32419 34198 32425
rect 34140 32385 34152 32419
rect 34186 32416 34198 32419
rect 35710 32416 35716 32428
rect 34186 32388 34928 32416
rect 35671 32388 35716 32416
rect 34186 32385 34198 32388
rect 34140 32379 34198 32385
rect 24820 32320 25820 32348
rect 25961 32351 26019 32357
rect 24820 32308 24826 32320
rect 25961 32317 25973 32351
rect 26007 32348 26019 32351
rect 27062 32348 27068 32360
rect 26007 32320 27068 32348
rect 26007 32317 26019 32320
rect 25961 32311 26019 32317
rect 27062 32308 27068 32320
rect 27120 32308 27126 32360
rect 31202 32348 31208 32360
rect 31163 32320 31208 32348
rect 31202 32308 31208 32320
rect 31260 32348 31266 32360
rect 31570 32348 31576 32360
rect 31260 32320 31576 32348
rect 31260 32308 31266 32320
rect 31570 32308 31576 32320
rect 31628 32308 31634 32360
rect 32493 32351 32551 32357
rect 32493 32317 32505 32351
rect 32539 32348 32551 32351
rect 32858 32348 32864 32360
rect 32539 32320 32864 32348
rect 32539 32317 32551 32320
rect 32493 32311 32551 32317
rect 32858 32308 32864 32320
rect 32916 32308 32922 32360
rect 33870 32348 33876 32360
rect 33831 32320 33876 32348
rect 33870 32308 33876 32320
rect 33928 32308 33934 32360
rect 34900 32348 34928 32388
rect 35710 32376 35716 32388
rect 35768 32376 35774 32428
rect 35802 32376 35808 32428
rect 35860 32416 35866 32428
rect 35989 32419 36047 32425
rect 35989 32416 36001 32419
rect 35860 32388 36001 32416
rect 35860 32376 35866 32388
rect 35989 32385 36001 32388
rect 36035 32385 36047 32419
rect 36722 32416 36728 32428
rect 36683 32388 36728 32416
rect 35989 32379 36047 32385
rect 36722 32376 36728 32388
rect 36780 32376 36786 32428
rect 37292 32425 37320 32456
rect 37522 32453 37534 32456
rect 37568 32453 37580 32487
rect 37522 32447 37580 32453
rect 37277 32419 37335 32425
rect 37277 32385 37289 32419
rect 37323 32385 37335 32419
rect 39114 32416 39120 32428
rect 39075 32388 39120 32416
rect 37277 32379 37335 32385
rect 39114 32376 39120 32388
rect 39172 32376 39178 32428
rect 39850 32376 39856 32428
rect 39908 32416 39914 32428
rect 40218 32425 40224 32428
rect 39945 32419 40003 32425
rect 39945 32416 39957 32419
rect 39908 32388 39957 32416
rect 39908 32376 39914 32388
rect 39945 32385 39957 32388
rect 39991 32385 40003 32419
rect 39945 32379 40003 32385
rect 40212 32379 40224 32425
rect 40276 32416 40282 32428
rect 40276 32388 40312 32416
rect 40218 32376 40224 32379
rect 40276 32376 40282 32388
rect 34900 32320 35756 32348
rect 20714 32280 20720 32292
rect 18156 32252 20720 32280
rect 18156 32212 18184 32252
rect 20714 32240 20720 32252
rect 20772 32280 20778 32292
rect 20993 32283 21051 32289
rect 20993 32280 21005 32283
rect 20772 32252 21005 32280
rect 20772 32240 20778 32252
rect 20993 32249 21005 32252
rect 21039 32249 21051 32283
rect 20993 32243 21051 32249
rect 30374 32240 30380 32292
rect 30432 32280 30438 32292
rect 31297 32283 31355 32289
rect 31297 32280 31309 32283
rect 30432 32252 31309 32280
rect 30432 32240 30438 32252
rect 31297 32249 31309 32252
rect 31343 32249 31355 32283
rect 31297 32243 31355 32249
rect 31386 32240 31392 32292
rect 31444 32280 31450 32292
rect 35728 32289 35756 32320
rect 36354 32308 36360 32360
rect 36412 32348 36418 32360
rect 36449 32351 36507 32357
rect 36449 32348 36461 32351
rect 36412 32320 36461 32348
rect 36412 32308 36418 32320
rect 36449 32317 36461 32320
rect 36495 32317 36507 32351
rect 36449 32311 36507 32317
rect 38930 32308 38936 32360
rect 38988 32348 38994 32360
rect 39209 32351 39267 32357
rect 39209 32348 39221 32351
rect 38988 32320 39221 32348
rect 38988 32308 38994 32320
rect 39209 32317 39221 32320
rect 39255 32348 39267 32351
rect 39482 32348 39488 32360
rect 39255 32320 39488 32348
rect 39255 32317 39267 32320
rect 39209 32311 39267 32317
rect 39482 32308 39488 32320
rect 39540 32308 39546 32360
rect 35713 32283 35771 32289
rect 31444 32252 31489 32280
rect 31444 32240 31450 32252
rect 35713 32249 35725 32283
rect 35759 32249 35771 32283
rect 35713 32243 35771 32249
rect 17236 32184 18184 32212
rect 18506 32172 18512 32224
rect 18564 32212 18570 32224
rect 19242 32212 19248 32224
rect 18564 32184 19248 32212
rect 18564 32172 18570 32184
rect 19242 32172 19248 32184
rect 19300 32172 19306 32224
rect 25314 32212 25320 32224
rect 25275 32184 25320 32212
rect 25314 32172 25320 32184
rect 25372 32172 25378 32224
rect 25498 32172 25504 32224
rect 25556 32212 25562 32224
rect 25777 32215 25835 32221
rect 25777 32212 25789 32215
rect 25556 32184 25789 32212
rect 25556 32172 25562 32184
rect 25777 32181 25789 32184
rect 25823 32212 25835 32215
rect 25866 32212 25872 32224
rect 25823 32184 25872 32212
rect 25823 32181 25835 32184
rect 25777 32175 25835 32181
rect 25866 32172 25872 32184
rect 25924 32172 25930 32224
rect 30745 32215 30803 32221
rect 30745 32181 30757 32215
rect 30791 32212 30803 32215
rect 31110 32212 31116 32224
rect 30791 32184 31116 32212
rect 30791 32181 30803 32184
rect 30745 32175 30803 32181
rect 31110 32172 31116 32184
rect 31168 32172 31174 32224
rect 34790 32172 34796 32224
rect 34848 32212 34854 32224
rect 35253 32215 35311 32221
rect 35253 32212 35265 32215
rect 34848 32184 35265 32212
rect 34848 32172 34854 32184
rect 35253 32181 35265 32184
rect 35299 32181 35311 32215
rect 35253 32175 35311 32181
rect 36633 32215 36691 32221
rect 36633 32181 36645 32215
rect 36679 32212 36691 32215
rect 36998 32212 37004 32224
rect 36679 32184 37004 32212
rect 36679 32181 36691 32184
rect 36633 32175 36691 32181
rect 36998 32172 37004 32184
rect 37056 32172 37062 32224
rect 39206 32212 39212 32224
rect 39167 32184 39212 32212
rect 39206 32172 39212 32184
rect 39264 32172 39270 32224
rect 39666 32172 39672 32224
rect 39724 32212 39730 32224
rect 41325 32215 41383 32221
rect 41325 32212 41337 32215
rect 39724 32184 41337 32212
rect 39724 32172 39730 32184
rect 41325 32181 41337 32184
rect 41371 32181 41383 32215
rect 41325 32175 41383 32181
rect 1104 32122 42872 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 42872 32122
rect 1104 32048 42872 32070
rect 16850 31968 16856 32020
rect 16908 32008 16914 32020
rect 17221 32011 17279 32017
rect 17221 32008 17233 32011
rect 16908 31980 17233 32008
rect 16908 31968 16914 31980
rect 17221 31977 17233 31980
rect 17267 31977 17279 32011
rect 18230 32008 18236 32020
rect 18191 31980 18236 32008
rect 17221 31971 17279 31977
rect 18230 31968 18236 31980
rect 18288 31968 18294 32020
rect 20070 31968 20076 32020
rect 20128 32008 20134 32020
rect 22462 32008 22468 32020
rect 20128 31980 22468 32008
rect 20128 31968 20134 31980
rect 22462 31968 22468 31980
rect 22520 31968 22526 32020
rect 24854 31968 24860 32020
rect 24912 32008 24918 32020
rect 24949 32011 25007 32017
rect 24949 32008 24961 32011
rect 24912 31980 24961 32008
rect 24912 31968 24918 31980
rect 24949 31977 24961 31980
rect 24995 31977 25007 32011
rect 27154 32008 27160 32020
rect 27115 31980 27160 32008
rect 24949 31971 25007 31977
rect 27154 31968 27160 31980
rect 27212 31968 27218 32020
rect 33870 32008 33876 32020
rect 30024 31980 33876 32008
rect 15473 31943 15531 31949
rect 15473 31909 15485 31943
rect 15519 31940 15531 31943
rect 15562 31940 15568 31952
rect 15519 31912 15568 31940
rect 15519 31909 15531 31912
rect 15473 31903 15531 31909
rect 15562 31900 15568 31912
rect 15620 31940 15626 31952
rect 15620 31912 15976 31940
rect 15620 31900 15626 31912
rect 14090 31872 14096 31884
rect 14051 31844 14096 31872
rect 14090 31832 14096 31844
rect 14148 31832 14154 31884
rect 15948 31881 15976 31912
rect 20254 31900 20260 31952
rect 20312 31940 20318 31952
rect 20622 31940 20628 31952
rect 20312 31912 20628 31940
rect 20312 31900 20318 31912
rect 20456 31881 20484 31912
rect 20622 31900 20628 31912
rect 20680 31900 20686 31952
rect 15933 31875 15991 31881
rect 15933 31841 15945 31875
rect 15979 31841 15991 31875
rect 15933 31835 15991 31841
rect 20349 31875 20407 31881
rect 20349 31841 20361 31875
rect 20395 31841 20407 31875
rect 20349 31835 20407 31841
rect 20441 31875 20499 31881
rect 20441 31841 20453 31875
rect 20487 31841 20499 31875
rect 20441 31835 20499 31841
rect 16206 31804 16212 31816
rect 16167 31776 16212 31804
rect 16206 31764 16212 31776
rect 16264 31764 16270 31816
rect 17402 31764 17408 31816
rect 17460 31804 17466 31816
rect 17770 31804 17776 31816
rect 17460 31776 17505 31804
rect 17731 31776 17776 31804
rect 17460 31764 17466 31776
rect 17770 31764 17776 31776
rect 17828 31764 17834 31816
rect 18414 31804 18420 31816
rect 18375 31776 18420 31804
rect 18414 31764 18420 31776
rect 18472 31764 18478 31816
rect 14366 31745 14372 31748
rect 14360 31699 14372 31745
rect 14424 31736 14430 31748
rect 14424 31708 14460 31736
rect 14366 31696 14372 31699
rect 14424 31696 14430 31708
rect 16942 31696 16948 31748
rect 17000 31736 17006 31748
rect 17497 31739 17555 31745
rect 17497 31736 17509 31739
rect 17000 31708 17509 31736
rect 17000 31696 17006 31708
rect 17497 31705 17509 31708
rect 17543 31705 17555 31739
rect 17497 31699 17555 31705
rect 17586 31696 17592 31748
rect 17644 31736 17650 31748
rect 20364 31736 20392 31835
rect 25498 31832 25504 31884
rect 25556 31872 25562 31884
rect 26697 31875 26755 31881
rect 25556 31844 26372 31872
rect 25556 31832 25562 31844
rect 20530 31804 20536 31816
rect 20491 31776 20536 31804
rect 20530 31764 20536 31776
rect 20588 31764 20594 31816
rect 20625 31807 20683 31813
rect 20625 31773 20637 31807
rect 20671 31804 20683 31807
rect 20806 31804 20812 31816
rect 20671 31776 20812 31804
rect 20671 31773 20683 31776
rect 20625 31767 20683 31773
rect 20806 31764 20812 31776
rect 20864 31764 20870 31816
rect 22646 31804 22652 31816
rect 22559 31776 22652 31804
rect 22646 31764 22652 31776
rect 22704 31804 22710 31816
rect 24670 31804 24676 31816
rect 22704 31776 24676 31804
rect 22704 31764 22710 31776
rect 24670 31764 24676 31776
rect 24728 31764 24734 31816
rect 24762 31764 24768 31816
rect 24820 31804 24826 31816
rect 24857 31807 24915 31813
rect 24857 31804 24869 31807
rect 24820 31776 24869 31804
rect 24820 31764 24826 31776
rect 24857 31773 24869 31776
rect 24903 31773 24915 31807
rect 24857 31767 24915 31773
rect 25958 31764 25964 31816
rect 26016 31804 26022 31816
rect 26344 31813 26372 31844
rect 26697 31841 26709 31875
rect 26743 31841 26755 31875
rect 26697 31835 26755 31841
rect 26053 31807 26111 31813
rect 26053 31804 26065 31807
rect 26016 31776 26065 31804
rect 26016 31764 26022 31776
rect 26053 31773 26065 31776
rect 26099 31773 26111 31807
rect 26216 31807 26274 31813
rect 26216 31804 26228 31807
rect 26053 31767 26111 31773
rect 26160 31776 26228 31804
rect 17644 31708 17689 31736
rect 20364 31708 21312 31736
rect 17644 31696 17650 31708
rect 20806 31668 20812 31680
rect 20767 31640 20812 31668
rect 20806 31628 20812 31640
rect 20864 31628 20870 31680
rect 21284 31677 21312 31708
rect 22094 31696 22100 31748
rect 22152 31736 22158 31748
rect 22382 31739 22440 31745
rect 22382 31736 22394 31739
rect 22152 31708 22394 31736
rect 22152 31696 22158 31708
rect 22382 31705 22394 31708
rect 22428 31705 22440 31739
rect 26160 31736 26188 31776
rect 26216 31773 26228 31776
rect 26262 31773 26274 31807
rect 26216 31767 26274 31773
rect 26332 31807 26390 31813
rect 26332 31773 26344 31807
rect 26378 31773 26390 31807
rect 26332 31767 26390 31773
rect 26418 31764 26424 31816
rect 26476 31813 26482 31816
rect 26476 31807 26499 31813
rect 26487 31773 26499 31807
rect 26712 31804 26740 31835
rect 28534 31832 28540 31884
rect 28592 31872 28598 31884
rect 28902 31872 28908 31884
rect 28592 31844 28908 31872
rect 28592 31832 28598 31844
rect 28902 31832 28908 31844
rect 28960 31872 28966 31884
rect 30024 31881 30052 31980
rect 33870 31968 33876 31980
rect 33928 31968 33934 32020
rect 32306 31940 32312 31952
rect 32267 31912 32312 31940
rect 32306 31900 32312 31912
rect 32364 31900 32370 31952
rect 30009 31875 30067 31881
rect 30009 31872 30021 31875
rect 28960 31844 30021 31872
rect 28960 31832 28966 31844
rect 30009 31841 30021 31844
rect 30055 31841 30067 31875
rect 31849 31875 31907 31881
rect 31849 31872 31861 31875
rect 30009 31835 30067 31841
rect 30208 31844 31861 31872
rect 30208 31813 30236 31844
rect 31849 31841 31861 31844
rect 31895 31872 31907 31875
rect 33134 31872 33140 31884
rect 31895 31844 33140 31872
rect 31895 31841 31907 31844
rect 31849 31835 31907 31841
rect 33134 31832 33140 31844
rect 33192 31832 33198 31884
rect 33597 31875 33655 31881
rect 33597 31841 33609 31875
rect 33643 31872 33655 31875
rect 34146 31872 34152 31884
rect 33643 31844 34152 31872
rect 33643 31841 33655 31844
rect 33597 31835 33655 31841
rect 34146 31832 34152 31844
rect 34204 31832 34210 31884
rect 34701 31875 34759 31881
rect 34701 31841 34713 31875
rect 34747 31872 34759 31875
rect 34790 31872 34796 31884
rect 34747 31844 34796 31872
rect 34747 31841 34759 31844
rect 34701 31835 34759 31841
rect 34790 31832 34796 31844
rect 34848 31832 34854 31884
rect 34974 31872 34980 31884
rect 34935 31844 34980 31872
rect 34974 31832 34980 31844
rect 35032 31832 35038 31884
rect 37918 31832 37924 31884
rect 37976 31872 37982 31884
rect 38381 31875 38439 31881
rect 38381 31872 38393 31875
rect 37976 31844 38393 31872
rect 37976 31832 37982 31844
rect 38381 31841 38393 31844
rect 38427 31841 38439 31875
rect 38654 31872 38660 31884
rect 38615 31844 38660 31872
rect 38381 31835 38439 31841
rect 38654 31832 38660 31844
rect 38712 31832 38718 31884
rect 41322 31872 41328 31884
rect 41283 31844 41328 31872
rect 41322 31832 41328 31844
rect 41380 31832 41386 31884
rect 28270 31807 28328 31813
rect 28270 31804 28282 31807
rect 26712 31776 28282 31804
rect 26476 31767 26499 31773
rect 28270 31773 28282 31776
rect 28316 31773 28328 31807
rect 28270 31767 28328 31773
rect 30193 31807 30251 31813
rect 30193 31773 30205 31807
rect 30239 31773 30251 31807
rect 30193 31767 30251 31773
rect 30929 31807 30987 31813
rect 30929 31773 30941 31807
rect 30975 31804 30987 31807
rect 31110 31804 31116 31816
rect 30975 31776 31009 31804
rect 31071 31776 31116 31804
rect 30975 31773 30987 31776
rect 30929 31767 30987 31773
rect 26476 31764 26482 31767
rect 26970 31736 26976 31748
rect 26160 31708 26976 31736
rect 22382 31699 22440 31705
rect 26970 31696 26976 31708
rect 27028 31696 27034 31748
rect 30944 31736 30972 31767
rect 31110 31764 31116 31776
rect 31168 31764 31174 31816
rect 31662 31804 31668 31816
rect 31623 31776 31668 31804
rect 31662 31764 31668 31776
rect 31720 31764 31726 31816
rect 32861 31807 32919 31813
rect 32861 31773 32873 31807
rect 32907 31804 32919 31807
rect 33318 31804 33324 31816
rect 32907 31776 33324 31804
rect 32907 31773 32919 31776
rect 32861 31767 32919 31773
rect 33318 31764 33324 31776
rect 33376 31764 33382 31816
rect 36998 31804 37004 31816
rect 36959 31776 37004 31804
rect 36998 31764 37004 31776
rect 37056 31764 37062 31816
rect 37274 31804 37280 31816
rect 37235 31776 37280 31804
rect 37274 31764 37280 31776
rect 37332 31764 37338 31816
rect 42150 31764 42156 31816
rect 42208 31804 42214 31816
rect 42208 31776 42253 31804
rect 42208 31764 42214 31776
rect 31294 31736 31300 31748
rect 30944 31708 31300 31736
rect 31294 31696 31300 31708
rect 31352 31696 31358 31748
rect 31386 31696 31392 31748
rect 31444 31736 31450 31748
rect 32677 31739 32735 31745
rect 32677 31736 32689 31739
rect 31444 31708 32689 31736
rect 31444 31696 31450 31708
rect 32324 31680 32352 31708
rect 32677 31705 32689 31708
rect 32723 31705 32735 31739
rect 41966 31736 41972 31748
rect 41927 31708 41972 31736
rect 32677 31699 32735 31705
rect 41966 31696 41972 31708
rect 42024 31696 42030 31748
rect 21269 31671 21327 31677
rect 21269 31637 21281 31671
rect 21315 31668 21327 31671
rect 22002 31668 22008 31680
rect 21315 31640 22008 31668
rect 21315 31637 21327 31640
rect 21269 31631 21327 31637
rect 22002 31628 22008 31640
rect 22060 31628 22066 31680
rect 25958 31628 25964 31680
rect 26016 31668 26022 31680
rect 29178 31668 29184 31680
rect 26016 31640 29184 31668
rect 26016 31628 26022 31640
rect 29178 31628 29184 31640
rect 29236 31628 29242 31680
rect 30745 31671 30803 31677
rect 30745 31637 30757 31671
rect 30791 31668 30803 31671
rect 30834 31668 30840 31680
rect 30791 31640 30840 31668
rect 30791 31637 30803 31640
rect 30745 31631 30803 31637
rect 30834 31628 30840 31640
rect 30892 31628 30898 31680
rect 32306 31628 32312 31680
rect 32364 31628 32370 31680
rect 32398 31628 32404 31680
rect 32456 31668 32462 31680
rect 32493 31671 32551 31677
rect 32493 31668 32505 31671
rect 32456 31640 32505 31668
rect 32456 31628 32462 31640
rect 32493 31637 32505 31640
rect 32539 31637 32551 31671
rect 32493 31631 32551 31637
rect 32585 31671 32643 31677
rect 32585 31637 32597 31671
rect 32631 31668 32643 31671
rect 33226 31668 33232 31680
rect 32631 31640 33232 31668
rect 32631 31637 32643 31640
rect 32585 31631 32643 31637
rect 33226 31628 33232 31640
rect 33284 31628 33290 31680
rect 33318 31628 33324 31680
rect 33376 31668 33382 31680
rect 34422 31668 34428 31680
rect 33376 31640 34428 31668
rect 33376 31628 33382 31640
rect 34422 31628 34428 31640
rect 34480 31628 34486 31680
rect 1104 31578 42872 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 42872 31578
rect 1104 31504 42872 31526
rect 14277 31467 14335 31473
rect 14277 31433 14289 31467
rect 14323 31464 14335 31467
rect 14366 31464 14372 31476
rect 14323 31436 14372 31464
rect 14323 31433 14335 31436
rect 14277 31427 14335 31433
rect 14366 31424 14372 31436
rect 14424 31424 14430 31476
rect 15930 31464 15936 31476
rect 15843 31436 15936 31464
rect 15930 31424 15936 31436
rect 15988 31464 15994 31476
rect 17770 31464 17776 31476
rect 15988 31436 17776 31464
rect 15988 31424 15994 31436
rect 17770 31424 17776 31436
rect 17828 31424 17834 31476
rect 21269 31467 21327 31473
rect 21269 31433 21281 31467
rect 21315 31464 21327 31467
rect 22094 31464 22100 31476
rect 21315 31436 22100 31464
rect 21315 31433 21327 31436
rect 21269 31427 21327 31433
rect 22094 31424 22100 31436
rect 22152 31424 22158 31476
rect 25038 31424 25044 31476
rect 25096 31464 25102 31476
rect 25958 31464 25964 31476
rect 25096 31436 25964 31464
rect 25096 31424 25102 31436
rect 25958 31424 25964 31436
rect 26016 31424 26022 31476
rect 26145 31467 26203 31473
rect 26145 31433 26157 31467
rect 26191 31464 26203 31467
rect 26234 31464 26240 31476
rect 26191 31436 26240 31464
rect 26191 31433 26203 31436
rect 26145 31427 26203 31433
rect 26234 31424 26240 31436
rect 26292 31424 26298 31476
rect 26970 31464 26976 31476
rect 26931 31436 26976 31464
rect 26970 31424 26976 31436
rect 27028 31424 27034 31476
rect 29638 31424 29644 31476
rect 29696 31464 29702 31476
rect 29825 31467 29883 31473
rect 29825 31464 29837 31467
rect 29696 31436 29837 31464
rect 29696 31424 29702 31436
rect 29825 31433 29837 31436
rect 29871 31433 29883 31467
rect 30834 31464 30840 31476
rect 29825 31427 29883 31433
rect 30484 31436 30840 31464
rect 15194 31396 15200 31408
rect 14568 31368 15200 31396
rect 14568 31337 14596 31368
rect 15194 31356 15200 31368
rect 15252 31356 15258 31408
rect 15562 31396 15568 31408
rect 15523 31368 15568 31396
rect 15562 31356 15568 31368
rect 15620 31356 15626 31408
rect 19978 31356 19984 31408
rect 20036 31396 20042 31408
rect 21913 31399 21971 31405
rect 21913 31396 21925 31399
rect 20036 31368 21925 31396
rect 20036 31356 20042 31368
rect 14553 31331 14611 31337
rect 14553 31297 14565 31331
rect 14599 31297 14611 31331
rect 14553 31291 14611 31297
rect 14645 31331 14703 31337
rect 14645 31297 14657 31331
rect 14691 31297 14703 31331
rect 14645 31291 14703 31297
rect 14366 31220 14372 31272
rect 14424 31260 14430 31272
rect 14660 31260 14688 31291
rect 14734 31288 14740 31340
rect 14792 31328 14798 31340
rect 14921 31331 14979 31337
rect 14792 31300 14837 31328
rect 14792 31288 14798 31300
rect 14921 31297 14933 31331
rect 14967 31297 14979 31331
rect 14921 31291 14979 31297
rect 15749 31331 15807 31337
rect 15749 31297 15761 31331
rect 15795 31328 15807 31331
rect 15838 31328 15844 31340
rect 15795 31300 15844 31328
rect 15795 31297 15807 31300
rect 15749 31291 15807 31297
rect 14424 31232 14688 31260
rect 14936 31260 14964 31291
rect 15838 31288 15844 31300
rect 15896 31328 15902 31340
rect 16669 31331 16727 31337
rect 16669 31328 16681 31331
rect 15896 31300 16681 31328
rect 15896 31288 15902 31300
rect 16669 31297 16681 31300
rect 16715 31297 16727 31331
rect 16942 31328 16948 31340
rect 16903 31300 16948 31328
rect 16669 31291 16727 31297
rect 16942 31288 16948 31300
rect 17000 31288 17006 31340
rect 20346 31288 20352 31340
rect 20404 31328 20410 31340
rect 20625 31331 20683 31337
rect 20625 31328 20637 31331
rect 20404 31300 20637 31328
rect 20404 31288 20410 31300
rect 20625 31297 20637 31300
rect 20671 31297 20683 31331
rect 20806 31328 20812 31340
rect 20767 31300 20812 31328
rect 20625 31291 20683 31297
rect 20806 31288 20812 31300
rect 20864 31288 20870 31340
rect 21008 31337 21036 31368
rect 21913 31365 21925 31368
rect 21959 31365 21971 31399
rect 24305 31399 24363 31405
rect 24305 31396 24317 31399
rect 21913 31359 21971 31365
rect 23308 31368 24317 31396
rect 20901 31331 20959 31337
rect 20901 31297 20913 31331
rect 20947 31297 20959 31331
rect 20901 31291 20959 31297
rect 20993 31331 21051 31337
rect 20993 31297 21005 31331
rect 21039 31297 21051 31331
rect 22002 31328 22008 31340
rect 21963 31300 22008 31328
rect 20993 31291 21051 31297
rect 16482 31260 16488 31272
rect 14936 31232 16488 31260
rect 14424 31220 14430 31232
rect 16482 31220 16488 31232
rect 16540 31220 16546 31272
rect 20916 31260 20944 31291
rect 22002 31288 22008 31300
rect 22060 31288 22066 31340
rect 21358 31260 21364 31272
rect 20916 31232 21364 31260
rect 21358 31220 21364 31232
rect 21416 31220 21422 31272
rect 21542 31220 21548 31272
rect 21600 31260 21606 31272
rect 23308 31260 23336 31368
rect 24305 31365 24317 31368
rect 24351 31396 24363 31399
rect 25682 31396 25688 31408
rect 24351 31368 25688 31396
rect 24351 31365 24363 31368
rect 24305 31359 24363 31365
rect 25682 31356 25688 31368
rect 25740 31356 25746 31408
rect 26252 31396 26280 31424
rect 26252 31368 27292 31396
rect 23382 31288 23388 31340
rect 23440 31328 23446 31340
rect 23440 31300 23485 31328
rect 23440 31288 23446 31300
rect 23566 31288 23572 31340
rect 23624 31328 23630 31340
rect 23624 31300 23669 31328
rect 23624 31288 23630 31300
rect 24210 31288 24216 31340
rect 24268 31328 24274 31340
rect 24489 31331 24547 31337
rect 24489 31328 24501 31331
rect 24268 31300 24501 31328
rect 24268 31288 24274 31300
rect 24489 31297 24501 31300
rect 24535 31328 24547 31331
rect 24762 31328 24768 31340
rect 24535 31300 24768 31328
rect 24535 31297 24547 31300
rect 24489 31291 24547 31297
rect 24762 31288 24768 31300
rect 24820 31288 24826 31340
rect 25866 31288 25872 31340
rect 25924 31328 25930 31340
rect 27264 31337 27292 31368
rect 27338 31356 27344 31408
rect 27396 31396 27402 31408
rect 28442 31396 28448 31408
rect 27396 31368 27476 31396
rect 28403 31368 28448 31396
rect 27396 31356 27402 31368
rect 27448 31337 27476 31368
rect 28442 31356 28448 31368
rect 28500 31356 28506 31408
rect 30374 31396 30380 31408
rect 29748 31368 30380 31396
rect 25961 31331 26019 31337
rect 25961 31328 25973 31331
rect 25924 31300 25973 31328
rect 25924 31288 25930 31300
rect 25961 31297 25973 31300
rect 26007 31297 26019 31331
rect 25961 31291 26019 31297
rect 26237 31331 26295 31337
rect 26237 31297 26249 31331
rect 26283 31297 26295 31331
rect 26237 31291 26295 31297
rect 27249 31331 27307 31337
rect 27249 31297 27261 31331
rect 27295 31297 27307 31331
rect 27249 31291 27307 31297
rect 27433 31331 27491 31337
rect 27433 31297 27445 31331
rect 27479 31297 27491 31331
rect 27433 31291 27491 31297
rect 28629 31331 28687 31337
rect 28629 31297 28641 31331
rect 28675 31328 28687 31331
rect 28994 31328 29000 31340
rect 28675 31300 29000 31328
rect 28675 31297 28687 31300
rect 28629 31291 28687 31297
rect 26252 31260 26280 31291
rect 28994 31288 29000 31300
rect 29052 31288 29058 31340
rect 29748 31337 29776 31368
rect 30374 31356 30380 31368
rect 30432 31356 30438 31408
rect 29733 31331 29791 31337
rect 29733 31297 29745 31331
rect 29779 31297 29791 31331
rect 29733 31291 29791 31297
rect 29917 31331 29975 31337
rect 29917 31297 29929 31331
rect 29963 31328 29975 31331
rect 30484 31328 30512 31436
rect 30834 31424 30840 31436
rect 30892 31424 30898 31476
rect 32306 31424 32312 31476
rect 32364 31473 32370 31476
rect 32364 31467 32383 31473
rect 32371 31433 32383 31467
rect 34054 31464 34060 31476
rect 34015 31436 34060 31464
rect 32364 31427 32383 31433
rect 32364 31424 32370 31427
rect 34054 31424 34060 31436
rect 34112 31424 34118 31476
rect 34422 31424 34428 31476
rect 34480 31464 34486 31476
rect 35621 31467 35679 31473
rect 35621 31464 35633 31467
rect 34480 31436 35633 31464
rect 34480 31424 34486 31436
rect 35621 31433 35633 31436
rect 35667 31433 35679 31467
rect 38286 31464 38292 31476
rect 38247 31436 38292 31464
rect 35621 31427 35679 31433
rect 38286 31424 38292 31436
rect 38344 31424 38350 31476
rect 38470 31464 38476 31476
rect 38431 31436 38476 31464
rect 38470 31424 38476 31436
rect 38528 31424 38534 31476
rect 39022 31424 39028 31476
rect 39080 31464 39086 31476
rect 39117 31467 39175 31473
rect 39117 31464 39129 31467
rect 39080 31436 39129 31464
rect 39080 31424 39086 31436
rect 39117 31433 39129 31436
rect 39163 31433 39175 31467
rect 39482 31464 39488 31476
rect 39443 31436 39488 31464
rect 39117 31427 39175 31433
rect 39482 31424 39488 31436
rect 39540 31424 39546 31476
rect 40218 31464 40224 31476
rect 40179 31436 40224 31464
rect 40218 31424 40224 31436
rect 40276 31424 40282 31476
rect 41506 31464 41512 31476
rect 41467 31436 41512 31464
rect 41506 31424 41512 31436
rect 41564 31424 41570 31476
rect 32125 31399 32183 31405
rect 30576 31368 32076 31396
rect 30576 31337 30604 31368
rect 29963 31300 30512 31328
rect 30561 31331 30619 31337
rect 29963 31297 29975 31300
rect 29917 31291 29975 31297
rect 30561 31297 30573 31331
rect 30607 31297 30619 31331
rect 30561 31291 30619 31297
rect 30745 31331 30803 31337
rect 30745 31297 30757 31331
rect 30791 31297 30803 31331
rect 30745 31291 30803 31297
rect 26326 31260 26332 31272
rect 21600 31232 23336 31260
rect 26239 31232 26332 31260
rect 21600 31220 21606 31232
rect 26326 31220 26332 31232
rect 26384 31260 26390 31272
rect 27154 31260 27160 31272
rect 26384 31232 27160 31260
rect 26384 31220 26390 31232
rect 27154 31220 27160 31232
rect 27212 31220 27218 31272
rect 27341 31263 27399 31269
rect 27341 31229 27353 31263
rect 27387 31229 27399 31263
rect 27341 31223 27399 31229
rect 10318 31152 10324 31204
rect 10376 31192 10382 31204
rect 26878 31192 26884 31204
rect 10376 31164 26884 31192
rect 10376 31152 10382 31164
rect 26878 31152 26884 31164
rect 26936 31152 26942 31204
rect 20346 31084 20352 31136
rect 20404 31124 20410 31136
rect 23290 31124 23296 31136
rect 20404 31096 23296 31124
rect 20404 31084 20410 31096
rect 23290 31084 23296 31096
rect 23348 31084 23354 31136
rect 23477 31127 23535 31133
rect 23477 31093 23489 31127
rect 23523 31124 23535 31127
rect 24854 31124 24860 31136
rect 23523 31096 24860 31124
rect 23523 31093 23535 31096
rect 23477 31087 23535 31093
rect 24854 31084 24860 31096
rect 24912 31084 24918 31136
rect 25777 31127 25835 31133
rect 25777 31093 25789 31127
rect 25823 31124 25835 31127
rect 25866 31124 25872 31136
rect 25823 31096 25872 31124
rect 25823 31093 25835 31096
rect 25777 31087 25835 31093
rect 25866 31084 25872 31096
rect 25924 31084 25930 31136
rect 25958 31084 25964 31136
rect 26016 31124 26022 31136
rect 27356 31124 27384 31223
rect 30760 31192 30788 31291
rect 30834 31288 30840 31340
rect 30892 31328 30898 31340
rect 31389 31331 31447 31337
rect 31389 31328 31401 31331
rect 30892 31300 31401 31328
rect 30892 31288 30898 31300
rect 31389 31297 31401 31300
rect 31435 31297 31447 31331
rect 31389 31291 31447 31297
rect 31481 31331 31539 31337
rect 31481 31297 31493 31331
rect 31527 31328 31539 31331
rect 31527 31300 31754 31328
rect 31527 31297 31539 31300
rect 31481 31291 31539 31297
rect 31205 31263 31263 31269
rect 31205 31229 31217 31263
rect 31251 31260 31263 31263
rect 31570 31260 31576 31272
rect 31251 31232 31576 31260
rect 31251 31229 31263 31232
rect 31205 31223 31263 31229
rect 31570 31220 31576 31232
rect 31628 31220 31634 31272
rect 31297 31195 31355 31201
rect 31297 31192 31309 31195
rect 30760 31164 31309 31192
rect 31297 31161 31309 31164
rect 31343 31161 31355 31195
rect 31297 31155 31355 31161
rect 26016 31096 27384 31124
rect 30745 31127 30803 31133
rect 26016 31084 26022 31096
rect 30745 31093 30757 31127
rect 30791 31124 30803 31127
rect 30834 31124 30840 31136
rect 30791 31096 30840 31124
rect 30791 31093 30803 31096
rect 30745 31087 30803 31093
rect 30834 31084 30840 31096
rect 30892 31084 30898 31136
rect 31726 31124 31754 31300
rect 32048 31192 32076 31368
rect 32125 31365 32137 31399
rect 32171 31396 32183 31399
rect 32214 31396 32220 31408
rect 32171 31368 32220 31396
rect 32171 31365 32183 31368
rect 32125 31359 32183 31365
rect 32214 31356 32220 31368
rect 32272 31356 32278 31408
rect 33134 31356 33140 31408
rect 33192 31396 33198 31408
rect 33413 31399 33471 31405
rect 33413 31396 33425 31399
rect 33192 31368 33425 31396
rect 33192 31356 33198 31368
rect 33413 31365 33425 31368
rect 33459 31365 33471 31399
rect 33413 31359 33471 31365
rect 33597 31399 33655 31405
rect 33597 31365 33609 31399
rect 33643 31396 33655 31399
rect 34514 31396 34520 31408
rect 33643 31368 34520 31396
rect 33643 31365 33655 31368
rect 33597 31359 33655 31365
rect 34514 31356 34520 31368
rect 34572 31356 34578 31408
rect 35526 31396 35532 31408
rect 34716 31368 35532 31396
rect 34241 31331 34299 31337
rect 34241 31297 34253 31331
rect 34287 31297 34299 31331
rect 34241 31291 34299 31297
rect 32493 31195 32551 31201
rect 32493 31192 32505 31195
rect 32048 31164 32505 31192
rect 32493 31161 32505 31164
rect 32539 31192 32551 31195
rect 32766 31192 32772 31204
rect 32539 31164 32772 31192
rect 32539 31161 32551 31164
rect 32493 31155 32551 31161
rect 32766 31152 32772 31164
rect 32824 31152 32830 31204
rect 34256 31192 34284 31291
rect 34422 31288 34428 31340
rect 34480 31328 34486 31340
rect 34716 31337 34744 31368
rect 35526 31356 35532 31368
rect 35584 31356 35590 31408
rect 35805 31399 35863 31405
rect 35805 31365 35817 31399
rect 35851 31396 35863 31399
rect 37274 31396 37280 31408
rect 35851 31368 37280 31396
rect 35851 31365 35863 31368
rect 35805 31359 35863 31365
rect 37274 31356 37280 31368
rect 37332 31396 37338 31408
rect 38197 31399 38255 31405
rect 38197 31396 38209 31399
rect 37332 31368 38209 31396
rect 37332 31356 37338 31368
rect 38197 31365 38209 31368
rect 38243 31365 38255 31399
rect 39666 31396 39672 31408
rect 38197 31359 38255 31365
rect 39316 31368 39672 31396
rect 34609 31331 34667 31337
rect 34609 31328 34621 31331
rect 34480 31300 34621 31328
rect 34480 31288 34486 31300
rect 34609 31297 34621 31300
rect 34655 31297 34667 31331
rect 34609 31291 34667 31297
rect 34701 31331 34759 31337
rect 34701 31297 34713 31331
rect 34747 31297 34759 31331
rect 35434 31328 35440 31340
rect 35395 31300 35440 31328
rect 34701 31291 34759 31297
rect 35434 31288 35440 31300
rect 35492 31288 35498 31340
rect 37918 31328 37924 31340
rect 37879 31300 37924 31328
rect 37918 31288 37924 31300
rect 37976 31288 37982 31340
rect 38105 31331 38163 31337
rect 38105 31297 38117 31331
rect 38151 31328 38163 31331
rect 38286 31328 38292 31340
rect 38151 31300 38292 31328
rect 38151 31297 38163 31300
rect 38105 31291 38163 31297
rect 38286 31288 38292 31300
rect 38344 31288 38350 31340
rect 39316 31337 39344 31368
rect 39666 31356 39672 31368
rect 39724 31356 39730 31408
rect 39301 31331 39359 31337
rect 39301 31297 39313 31331
rect 39347 31297 39359 31331
rect 39301 31291 39359 31297
rect 39574 31288 39580 31340
rect 39632 31328 39638 31340
rect 39632 31300 39677 31328
rect 39632 31288 39638 31300
rect 39942 31288 39948 31340
rect 40000 31328 40006 31340
rect 40037 31331 40095 31337
rect 40037 31328 40049 31331
rect 40000 31300 40049 31328
rect 40000 31288 40006 31300
rect 40037 31297 40049 31300
rect 40083 31297 40095 31331
rect 40037 31291 40095 31297
rect 40310 31288 40316 31340
rect 40368 31328 40374 31340
rect 40773 31331 40831 31337
rect 40773 31328 40785 31331
rect 40368 31300 40785 31328
rect 40368 31288 40374 31300
rect 40773 31297 40785 31300
rect 40819 31297 40831 31331
rect 41414 31328 41420 31340
rect 41375 31300 41420 31328
rect 40773 31291 40831 31297
rect 41414 31288 41420 31300
rect 41472 31288 41478 31340
rect 34790 31192 34796 31204
rect 34256 31164 34796 31192
rect 34790 31152 34796 31164
rect 34848 31152 34854 31204
rect 34974 31152 34980 31204
rect 35032 31152 35038 31204
rect 35253 31195 35311 31201
rect 35253 31161 35265 31195
rect 35299 31161 35311 31195
rect 35253 31155 35311 31161
rect 32309 31127 32367 31133
rect 32309 31124 32321 31127
rect 31726 31096 32321 31124
rect 32309 31093 32321 31096
rect 32355 31124 32367 31127
rect 32398 31124 32404 31136
rect 32355 31096 32404 31124
rect 32355 31093 32367 31096
rect 32309 31087 32367 31093
rect 32398 31084 32404 31096
rect 32456 31084 32462 31136
rect 34330 31124 34336 31136
rect 34291 31096 34336 31124
rect 34330 31084 34336 31096
rect 34388 31084 34394 31136
rect 34698 31084 34704 31136
rect 34756 31124 34762 31136
rect 34992 31124 35020 31152
rect 35268 31124 35296 31155
rect 34756 31096 35296 31124
rect 34756 31084 34762 31096
rect 1104 31034 42872 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 42872 31034
rect 1104 30960 42872 30982
rect 14734 30880 14740 30932
rect 14792 30920 14798 30932
rect 15013 30923 15071 30929
rect 15013 30920 15025 30923
rect 14792 30892 15025 30920
rect 14792 30880 14798 30892
rect 15013 30889 15025 30892
rect 15059 30889 15071 30923
rect 15194 30920 15200 30932
rect 15013 30883 15071 30889
rect 15120 30892 15200 30920
rect 15120 30852 15148 30892
rect 15194 30880 15200 30892
rect 15252 30920 15258 30932
rect 16206 30920 16212 30932
rect 15252 30892 16212 30920
rect 15252 30880 15258 30892
rect 16206 30880 16212 30892
rect 16264 30880 16270 30932
rect 17586 30920 17592 30932
rect 17547 30892 17592 30920
rect 17586 30880 17592 30892
rect 17644 30880 17650 30932
rect 21358 30920 21364 30932
rect 21319 30892 21364 30920
rect 21358 30880 21364 30892
rect 21416 30880 21422 30932
rect 22554 30920 22560 30932
rect 22515 30892 22560 30920
rect 22554 30880 22560 30892
rect 22612 30880 22618 30932
rect 23290 30880 23296 30932
rect 23348 30920 23354 30932
rect 25038 30920 25044 30932
rect 23348 30892 25044 30920
rect 23348 30880 23354 30892
rect 25038 30880 25044 30892
rect 25096 30880 25102 30932
rect 25774 30920 25780 30932
rect 25735 30892 25780 30920
rect 25774 30880 25780 30892
rect 25832 30880 25838 30932
rect 26878 30880 26884 30932
rect 26936 30920 26942 30932
rect 32125 30923 32183 30929
rect 26936 30892 31754 30920
rect 26936 30880 26942 30892
rect 16574 30852 16580 30864
rect 14936 30824 15148 30852
rect 15580 30824 16580 30852
rect 14277 30719 14335 30725
rect 14277 30685 14289 30719
rect 14323 30685 14335 30719
rect 14277 30679 14335 30685
rect 13722 30608 13728 30660
rect 13780 30648 13786 30660
rect 14292 30648 14320 30679
rect 14366 30676 14372 30728
rect 14424 30716 14430 30728
rect 14936 30725 14964 30824
rect 14921 30719 14979 30725
rect 14424 30688 14469 30716
rect 14424 30676 14430 30688
rect 14921 30685 14933 30719
rect 14967 30685 14979 30719
rect 14921 30679 14979 30685
rect 15105 30719 15163 30725
rect 15105 30685 15117 30719
rect 15151 30716 15163 30719
rect 15580 30716 15608 30824
rect 16574 30812 16580 30824
rect 16632 30812 16638 30864
rect 20990 30812 20996 30864
rect 21048 30852 21054 30864
rect 25130 30852 25136 30864
rect 21048 30824 23428 30852
rect 21048 30812 21054 30824
rect 19242 30784 19248 30796
rect 16546 30756 19248 30784
rect 16546 30728 16574 30756
rect 19242 30744 19248 30756
rect 19300 30744 19306 30796
rect 20441 30787 20499 30793
rect 20441 30753 20453 30787
rect 20487 30784 20499 30787
rect 20806 30784 20812 30796
rect 20487 30756 20812 30784
rect 20487 30753 20499 30756
rect 20441 30747 20499 30753
rect 20806 30744 20812 30756
rect 20864 30744 20870 30796
rect 23293 30787 23351 30793
rect 23293 30784 23305 30787
rect 21836 30756 23305 30784
rect 15151 30688 15608 30716
rect 15749 30719 15807 30725
rect 15151 30685 15163 30688
rect 15105 30679 15163 30685
rect 15749 30685 15761 30719
rect 15795 30685 15807 30719
rect 15749 30679 15807 30685
rect 15841 30719 15899 30725
rect 15841 30685 15853 30719
rect 15887 30716 15899 30719
rect 16206 30716 16212 30728
rect 15887 30688 16212 30716
rect 15887 30685 15899 30688
rect 15841 30679 15899 30685
rect 15654 30648 15660 30660
rect 13780 30620 15660 30648
rect 13780 30608 13786 30620
rect 15654 30608 15660 30620
rect 15712 30608 15718 30660
rect 14093 30583 14151 30589
rect 14093 30549 14105 30583
rect 14139 30580 14151 30583
rect 14182 30580 14188 30592
rect 14139 30552 14188 30580
rect 14139 30549 14151 30552
rect 14093 30543 14151 30549
rect 14182 30540 14188 30552
rect 14240 30540 14246 30592
rect 15764 30580 15792 30679
rect 16206 30676 16212 30688
rect 16264 30676 16270 30728
rect 16482 30676 16488 30728
rect 16540 30716 16574 30728
rect 16666 30716 16672 30728
rect 16540 30688 16585 30716
rect 16627 30688 16672 30716
rect 16540 30679 16549 30688
rect 16540 30676 16546 30679
rect 16666 30676 16672 30688
rect 16724 30676 16730 30728
rect 16761 30719 16819 30725
rect 16761 30685 16773 30719
rect 16807 30685 16819 30719
rect 16761 30679 16819 30685
rect 16853 30719 16911 30725
rect 16853 30685 16865 30719
rect 16899 30716 16911 30719
rect 17218 30716 17224 30728
rect 16899 30688 17224 30716
rect 16899 30685 16911 30688
rect 16853 30679 16911 30685
rect 16025 30651 16083 30657
rect 16025 30617 16037 30651
rect 16071 30648 16083 30651
rect 16776 30648 16804 30679
rect 17218 30676 17224 30688
rect 17276 30676 17282 30728
rect 17589 30719 17647 30725
rect 17589 30685 17601 30719
rect 17635 30685 17647 30719
rect 17770 30716 17776 30728
rect 17731 30688 17776 30716
rect 17589 30679 17647 30685
rect 17604 30648 17632 30679
rect 17770 30676 17776 30688
rect 17828 30676 17834 30728
rect 20622 30716 20628 30728
rect 20583 30688 20628 30716
rect 20622 30676 20628 30688
rect 20680 30676 20686 30728
rect 20901 30719 20959 30725
rect 20901 30685 20913 30719
rect 20947 30716 20959 30719
rect 20990 30716 20996 30728
rect 20947 30688 20996 30716
rect 20947 30685 20959 30688
rect 20901 30679 20959 30685
rect 20990 30676 20996 30688
rect 21048 30676 21054 30728
rect 21542 30716 21548 30728
rect 21503 30688 21548 30716
rect 21542 30676 21548 30688
rect 21600 30676 21606 30728
rect 21836 30725 21864 30756
rect 23293 30753 23305 30756
rect 23339 30753 23351 30787
rect 23293 30747 23351 30753
rect 23400 30725 23428 30824
rect 24688 30824 25136 30852
rect 21821 30719 21879 30725
rect 21821 30685 21833 30719
rect 21867 30685 21879 30719
rect 23201 30719 23259 30725
rect 23201 30716 23213 30719
rect 21821 30679 21879 30685
rect 21928 30688 23213 30716
rect 16071 30620 17632 30648
rect 20640 30648 20668 30676
rect 21928 30648 21956 30688
rect 23201 30685 23213 30688
rect 23247 30685 23259 30719
rect 23201 30679 23259 30685
rect 23385 30719 23443 30725
rect 23385 30685 23397 30719
rect 23431 30685 23443 30719
rect 23385 30679 23443 30685
rect 23566 30676 23572 30728
rect 23624 30716 23630 30728
rect 24688 30725 24716 30824
rect 25130 30812 25136 30824
rect 25188 30812 25194 30864
rect 28813 30855 28871 30861
rect 28813 30821 28825 30855
rect 28859 30852 28871 30855
rect 28994 30852 29000 30864
rect 28859 30824 29000 30852
rect 28859 30821 28871 30824
rect 28813 30815 28871 30821
rect 28994 30812 29000 30824
rect 29052 30812 29058 30864
rect 31726 30852 31754 30892
rect 32125 30889 32137 30923
rect 32171 30920 32183 30923
rect 32398 30920 32404 30932
rect 32171 30892 32404 30920
rect 32171 30889 32183 30892
rect 32125 30883 32183 30889
rect 32398 30880 32404 30892
rect 32456 30880 32462 30932
rect 32766 30920 32772 30932
rect 32727 30892 32772 30920
rect 32766 30880 32772 30892
rect 32824 30880 32830 30932
rect 34330 30880 34336 30932
rect 34388 30920 34394 30932
rect 34885 30923 34943 30929
rect 34885 30920 34897 30923
rect 34388 30892 34897 30920
rect 34388 30880 34394 30892
rect 34885 30889 34897 30892
rect 34931 30920 34943 30923
rect 35069 30923 35127 30929
rect 34931 30892 35020 30920
rect 34931 30889 34943 30892
rect 34885 30883 34943 30889
rect 34790 30852 34796 30864
rect 31726 30824 34796 30852
rect 34790 30812 34796 30824
rect 34848 30812 34854 30864
rect 34992 30852 35020 30892
rect 35069 30889 35081 30923
rect 35115 30920 35127 30923
rect 35342 30920 35348 30932
rect 35115 30892 35348 30920
rect 35115 30889 35127 30892
rect 35069 30883 35127 30889
rect 35342 30880 35348 30892
rect 35400 30920 35406 30932
rect 35621 30923 35679 30929
rect 35621 30920 35633 30923
rect 35400 30892 35633 30920
rect 35400 30880 35406 30892
rect 35621 30889 35633 30892
rect 35667 30889 35679 30923
rect 38562 30920 38568 30932
rect 38523 30892 38568 30920
rect 35621 30883 35679 30889
rect 38562 30880 38568 30892
rect 38620 30880 38626 30932
rect 38749 30923 38807 30929
rect 38749 30889 38761 30923
rect 38795 30920 38807 30923
rect 39114 30920 39120 30932
rect 38795 30892 39120 30920
rect 38795 30889 38807 30892
rect 38749 30883 38807 30889
rect 39114 30880 39120 30892
rect 39172 30920 39178 30932
rect 39574 30920 39580 30932
rect 39172 30892 39580 30920
rect 39172 30880 39178 30892
rect 39574 30880 39580 30892
rect 39632 30880 39638 30932
rect 41509 30923 41567 30929
rect 41509 30889 41521 30923
rect 41555 30920 41567 30923
rect 41966 30920 41972 30932
rect 41555 30892 41972 30920
rect 41555 30889 41567 30892
rect 41509 30883 41567 30889
rect 41966 30880 41972 30892
rect 42024 30880 42030 30932
rect 34992 30824 35112 30852
rect 27157 30787 27215 30793
rect 27157 30753 27169 30787
rect 27203 30784 27215 30787
rect 28534 30784 28540 30796
rect 27203 30756 28540 30784
rect 27203 30753 27215 30756
rect 27157 30747 27215 30753
rect 28534 30744 28540 30756
rect 28592 30744 28598 30796
rect 32585 30787 32643 30793
rect 32585 30753 32597 30787
rect 32631 30784 32643 30787
rect 35084 30784 35112 30824
rect 35158 30812 35164 30864
rect 35216 30852 35222 30864
rect 35216 30824 41460 30852
rect 35216 30812 35222 30824
rect 35434 30784 35440 30796
rect 32631 30756 34836 30784
rect 35084 30756 35440 30784
rect 32631 30753 32643 30756
rect 32585 30747 32643 30753
rect 24880 30725 24886 30728
rect 24673 30719 24731 30725
rect 24673 30716 24685 30719
rect 23624 30688 24685 30716
rect 23624 30676 23630 30688
rect 24673 30685 24685 30688
rect 24719 30685 24731 30719
rect 24673 30679 24731 30685
rect 24765 30719 24823 30725
rect 24765 30685 24777 30719
rect 24811 30685 24823 30719
rect 24765 30679 24823 30685
rect 24862 30719 24886 30725
rect 24862 30685 24874 30719
rect 24862 30679 24886 30685
rect 22646 30648 22652 30660
rect 20640 30620 21956 30648
rect 22607 30620 22652 30648
rect 16071 30617 16083 30620
rect 16025 30611 16083 30617
rect 22646 30608 22652 30620
rect 22704 30608 22710 30660
rect 24780 30648 24808 30679
rect 24880 30676 24886 30679
rect 24938 30676 24944 30728
rect 25038 30716 25044 30728
rect 24999 30688 25044 30716
rect 25038 30676 25044 30688
rect 25096 30676 25102 30728
rect 27062 30676 27068 30728
rect 27120 30716 27126 30728
rect 27801 30719 27859 30725
rect 27801 30716 27813 30719
rect 27120 30688 27813 30716
rect 27120 30676 27126 30688
rect 27801 30685 27813 30688
rect 27847 30685 27859 30719
rect 27801 30679 27859 30685
rect 30374 30676 30380 30728
rect 30432 30716 30438 30728
rect 30745 30719 30803 30725
rect 30745 30716 30757 30719
rect 30432 30688 30757 30716
rect 30432 30676 30438 30688
rect 30745 30685 30757 30688
rect 30791 30685 30803 30719
rect 30745 30679 30803 30685
rect 30834 30676 30840 30728
rect 30892 30716 30898 30728
rect 31001 30719 31059 30725
rect 31001 30716 31013 30719
rect 30892 30688 31013 30716
rect 30892 30676 30898 30688
rect 31001 30685 31013 30688
rect 31047 30685 31059 30719
rect 31001 30679 31059 30685
rect 31570 30676 31576 30728
rect 31628 30716 31634 30728
rect 32600 30716 32628 30747
rect 31628 30688 32628 30716
rect 32861 30719 32919 30725
rect 31628 30676 31634 30688
rect 32861 30685 32873 30719
rect 32907 30716 32919 30719
rect 33226 30716 33232 30728
rect 32907 30688 33232 30716
rect 32907 30685 32919 30688
rect 32861 30679 32919 30685
rect 33226 30676 33232 30688
rect 33284 30716 33290 30728
rect 33962 30716 33968 30728
rect 33284 30688 33968 30716
rect 33284 30676 33290 30688
rect 33962 30676 33968 30688
rect 34020 30716 34026 30728
rect 34422 30716 34428 30728
rect 34020 30688 34428 30716
rect 34020 30676 34026 30688
rect 34422 30676 34428 30688
rect 34480 30676 34486 30728
rect 26234 30648 26240 30660
rect 24780 30620 26240 30648
rect 26234 30608 26240 30620
rect 26292 30608 26298 30660
rect 26912 30651 26970 30657
rect 26912 30617 26924 30651
rect 26958 30648 26970 30651
rect 26958 30620 27660 30648
rect 26958 30617 26970 30620
rect 26912 30611 26970 30617
rect 15838 30580 15844 30592
rect 15751 30552 15844 30580
rect 15838 30540 15844 30552
rect 15896 30580 15902 30592
rect 16942 30580 16948 30592
rect 15896 30552 16948 30580
rect 15896 30540 15902 30552
rect 16942 30540 16948 30552
rect 17000 30540 17006 30592
rect 17129 30583 17187 30589
rect 17129 30549 17141 30583
rect 17175 30580 17187 30583
rect 18230 30580 18236 30592
rect 17175 30552 18236 30580
rect 17175 30549 17187 30552
rect 17129 30543 17187 30549
rect 18230 30540 18236 30552
rect 18288 30540 18294 30592
rect 20530 30540 20536 30592
rect 20588 30580 20594 30592
rect 20809 30583 20867 30589
rect 20809 30580 20821 30583
rect 20588 30552 20821 30580
rect 20588 30540 20594 30552
rect 20809 30549 20821 30552
rect 20855 30580 20867 30583
rect 21729 30583 21787 30589
rect 21729 30580 21741 30583
rect 20855 30552 21741 30580
rect 20855 30549 20867 30552
rect 20809 30543 20867 30549
rect 21729 30549 21741 30552
rect 21775 30549 21787 30583
rect 24394 30580 24400 30592
rect 24355 30552 24400 30580
rect 21729 30543 21787 30549
rect 24394 30540 24400 30552
rect 24452 30540 24458 30592
rect 27632 30589 27660 30620
rect 28442 30608 28448 30660
rect 28500 30648 28506 30660
rect 28626 30648 28632 30660
rect 28500 30620 28632 30648
rect 28500 30608 28506 30620
rect 28626 30608 28632 30620
rect 28684 30608 28690 30660
rect 33410 30608 33416 30660
rect 33468 30648 33474 30660
rect 34698 30648 34704 30660
rect 33468 30620 34704 30648
rect 33468 30608 33474 30620
rect 34698 30608 34704 30620
rect 34756 30608 34762 30660
rect 34808 30648 34836 30756
rect 35434 30744 35440 30756
rect 35492 30744 35498 30796
rect 35618 30744 35624 30796
rect 35676 30784 35682 30796
rect 35805 30787 35863 30793
rect 35805 30784 35817 30787
rect 35676 30756 35817 30784
rect 35676 30744 35682 30756
rect 35805 30753 35817 30756
rect 35851 30753 35863 30787
rect 37918 30784 37924 30796
rect 35805 30747 35863 30753
rect 37568 30756 37924 30784
rect 35526 30716 35532 30728
rect 35487 30688 35532 30716
rect 35526 30676 35532 30688
rect 35584 30676 35590 30728
rect 35636 30648 35664 30744
rect 36265 30719 36323 30725
rect 36265 30716 36277 30719
rect 35820 30688 36277 30716
rect 35820 30657 35848 30688
rect 36265 30685 36277 30688
rect 36311 30685 36323 30719
rect 36265 30679 36323 30685
rect 36449 30719 36507 30725
rect 36449 30685 36461 30719
rect 36495 30716 36507 30719
rect 36998 30716 37004 30728
rect 36495 30688 37004 30716
rect 36495 30685 36507 30688
rect 36449 30679 36507 30685
rect 36998 30676 37004 30688
rect 37056 30716 37062 30728
rect 37568 30725 37596 30756
rect 37918 30744 37924 30756
rect 37976 30784 37982 30796
rect 37976 30756 38424 30784
rect 37976 30744 37982 30756
rect 37461 30719 37519 30725
rect 37461 30716 37473 30719
rect 37056 30688 37473 30716
rect 37056 30676 37062 30688
rect 37461 30685 37473 30688
rect 37507 30685 37519 30719
rect 37461 30679 37519 30685
rect 37553 30719 37611 30725
rect 37553 30685 37565 30719
rect 37599 30685 37611 30719
rect 37553 30679 37611 30685
rect 37737 30719 37795 30725
rect 37737 30685 37749 30719
rect 37783 30716 37795 30719
rect 38286 30716 38292 30728
rect 37783 30688 38292 30716
rect 37783 30685 37795 30688
rect 37737 30679 37795 30685
rect 34808 30620 35664 30648
rect 35805 30651 35863 30657
rect 35805 30617 35817 30651
rect 35851 30617 35863 30651
rect 37476 30648 37504 30679
rect 38286 30676 38292 30688
rect 38344 30676 38350 30728
rect 38396 30657 38424 30756
rect 41432 30725 41460 30824
rect 41417 30719 41475 30725
rect 41417 30685 41429 30719
rect 41463 30716 41475 30719
rect 41874 30716 41880 30728
rect 41463 30688 41880 30716
rect 41463 30685 41475 30688
rect 41417 30679 41475 30685
rect 41874 30676 41880 30688
rect 41932 30676 41938 30728
rect 38381 30651 38439 30657
rect 37476 30620 38056 30648
rect 35805 30611 35863 30617
rect 27617 30583 27675 30589
rect 27617 30549 27629 30583
rect 27663 30549 27675 30583
rect 27617 30543 27675 30549
rect 32585 30583 32643 30589
rect 32585 30549 32597 30583
rect 32631 30580 32643 30583
rect 32674 30580 32680 30592
rect 32631 30552 32680 30580
rect 32631 30549 32643 30552
rect 32585 30543 32643 30549
rect 32674 30540 32680 30552
rect 32732 30540 32738 30592
rect 34146 30540 34152 30592
rect 34204 30580 34210 30592
rect 34901 30583 34959 30589
rect 34901 30580 34913 30583
rect 34204 30552 34913 30580
rect 34204 30540 34210 30552
rect 34901 30549 34913 30552
rect 34947 30549 34959 30583
rect 34901 30543 34959 30549
rect 36357 30583 36415 30589
rect 36357 30549 36369 30583
rect 36403 30580 36415 30583
rect 36446 30580 36452 30592
rect 36403 30552 36452 30580
rect 36403 30549 36415 30552
rect 36357 30543 36415 30549
rect 36446 30540 36452 30552
rect 36504 30540 36510 30592
rect 37918 30580 37924 30592
rect 37879 30552 37924 30580
rect 37918 30540 37924 30552
rect 37976 30540 37982 30592
rect 38028 30580 38056 30620
rect 38381 30617 38393 30651
rect 38427 30617 38439 30651
rect 38381 30611 38439 30617
rect 38581 30583 38639 30589
rect 38581 30580 38593 30583
rect 38028 30552 38593 30580
rect 38581 30549 38593 30552
rect 38627 30549 38639 30583
rect 38581 30543 38639 30549
rect 1104 30490 42872 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 42872 30490
rect 1104 30416 42872 30438
rect 13173 30379 13231 30385
rect 13173 30345 13185 30379
rect 13219 30376 13231 30379
rect 13998 30376 14004 30388
rect 13219 30348 14004 30376
rect 13219 30345 13231 30348
rect 13173 30339 13231 30345
rect 13998 30336 14004 30348
rect 14056 30336 14062 30388
rect 14366 30336 14372 30388
rect 14424 30376 14430 30388
rect 15105 30379 15163 30385
rect 15105 30376 15117 30379
rect 14424 30348 15117 30376
rect 14424 30336 14430 30348
rect 15105 30345 15117 30348
rect 15151 30345 15163 30379
rect 16666 30376 16672 30388
rect 16627 30348 16672 30376
rect 15105 30339 15163 30345
rect 16666 30336 16672 30348
rect 16724 30336 16730 30388
rect 20743 30379 20801 30385
rect 20456 30348 20668 30376
rect 14918 30308 14924 30320
rect 14292 30280 14924 30308
rect 13081 30243 13139 30249
rect 13081 30209 13093 30243
rect 13127 30209 13139 30243
rect 13081 30203 13139 30209
rect 13357 30243 13415 30249
rect 13357 30209 13369 30243
rect 13403 30240 13415 30243
rect 13403 30212 13952 30240
rect 13403 30209 13415 30212
rect 13357 30203 13415 30209
rect 13096 30172 13124 30203
rect 13722 30172 13728 30184
rect 13096 30144 13728 30172
rect 13722 30132 13728 30144
rect 13780 30132 13786 30184
rect 13924 30172 13952 30212
rect 13998 30200 14004 30252
rect 14056 30240 14062 30252
rect 14182 30240 14188 30252
rect 14056 30212 14101 30240
rect 14143 30212 14188 30240
rect 14056 30200 14062 30212
rect 14182 30200 14188 30212
rect 14240 30200 14246 30252
rect 14292 30249 14320 30280
rect 14918 30268 14924 30280
rect 14976 30308 14982 30320
rect 20456 30308 20484 30348
rect 14976 30280 20484 30308
rect 20533 30311 20591 30317
rect 14976 30268 14982 30280
rect 14277 30243 14335 30249
rect 14277 30209 14289 30243
rect 14323 30209 14335 30243
rect 14277 30203 14335 30209
rect 14369 30243 14427 30249
rect 14369 30209 14381 30243
rect 14415 30240 14427 30243
rect 14458 30240 14464 30252
rect 14415 30212 14464 30240
rect 14415 30209 14427 30212
rect 14369 30203 14427 30209
rect 14458 30200 14464 30212
rect 14516 30200 14522 30252
rect 14550 30200 14556 30252
rect 14608 30240 14614 30252
rect 14826 30240 14832 30252
rect 14608 30212 14832 30240
rect 14608 30200 14614 30212
rect 14826 30200 14832 30212
rect 14884 30200 14890 30252
rect 17328 30249 17356 30280
rect 20533 30277 20545 30311
rect 20579 30277 20591 30311
rect 20640 30308 20668 30348
rect 20743 30345 20755 30379
rect 20789 30376 20801 30379
rect 21358 30376 21364 30388
rect 20789 30348 21364 30376
rect 20789 30345 20801 30348
rect 20743 30339 20801 30345
rect 21358 30336 21364 30348
rect 21416 30336 21422 30388
rect 23293 30379 23351 30385
rect 23293 30345 23305 30379
rect 23339 30376 23351 30379
rect 23566 30376 23572 30388
rect 23339 30348 23572 30376
rect 23339 30345 23351 30348
rect 23293 30339 23351 30345
rect 23566 30336 23572 30348
rect 23624 30336 23630 30388
rect 25498 30376 25504 30388
rect 25459 30348 25504 30376
rect 25498 30336 25504 30348
rect 25556 30336 25562 30388
rect 25869 30379 25927 30385
rect 25869 30345 25881 30379
rect 25915 30376 25927 30379
rect 26234 30376 26240 30388
rect 25915 30348 26240 30376
rect 25915 30345 25927 30348
rect 25869 30339 25927 30345
rect 26234 30336 26240 30348
rect 26292 30336 26298 30388
rect 27985 30379 28043 30385
rect 27985 30345 27997 30379
rect 28031 30345 28043 30379
rect 34146 30376 34152 30388
rect 27985 30339 28043 30345
rect 33336 30348 34152 30376
rect 21542 30308 21548 30320
rect 20640 30280 21548 30308
rect 20533 30271 20591 30277
rect 15197 30243 15255 30249
rect 15197 30209 15209 30243
rect 15243 30240 15255 30243
rect 16945 30243 17003 30249
rect 16945 30240 16957 30243
rect 15243 30212 16957 30240
rect 15243 30209 15255 30212
rect 15197 30203 15255 30209
rect 16945 30209 16957 30212
rect 16991 30209 17003 30243
rect 16945 30203 17003 30209
rect 17313 30243 17371 30249
rect 17313 30209 17325 30243
rect 17359 30209 17371 30243
rect 17313 30203 17371 30209
rect 17865 30243 17923 30249
rect 17865 30209 17877 30243
rect 17911 30241 17923 30243
rect 18049 30243 18107 30249
rect 17911 30213 18000 30241
rect 17911 30209 17923 30213
rect 17865 30203 17923 30209
rect 15212 30172 15240 30203
rect 13924 30144 15240 30172
rect 15746 30132 15752 30184
rect 15804 30172 15810 30184
rect 16853 30175 16911 30181
rect 16853 30172 16865 30175
rect 15804 30144 16865 30172
rect 15804 30132 15810 30144
rect 16853 30141 16865 30144
rect 16899 30141 16911 30175
rect 16853 30135 16911 30141
rect 11974 30064 11980 30116
rect 12032 30104 12038 30116
rect 13817 30107 13875 30113
rect 13817 30104 13829 30107
rect 12032 30076 13829 30104
rect 12032 30064 12038 30076
rect 13817 30073 13829 30076
rect 13863 30073 13875 30107
rect 16960 30104 16988 30203
rect 17218 30172 17224 30184
rect 17179 30144 17224 30172
rect 17218 30132 17224 30144
rect 17276 30132 17282 30184
rect 17972 30172 18000 30213
rect 18049 30209 18061 30243
rect 18095 30240 18107 30243
rect 18506 30240 18512 30252
rect 18095 30212 18512 30240
rect 18095 30209 18107 30212
rect 18049 30203 18107 30209
rect 18506 30200 18512 30212
rect 18564 30200 18570 30252
rect 19633 30243 19691 30249
rect 19633 30209 19645 30243
rect 19679 30240 19691 30243
rect 19794 30240 19800 30252
rect 19679 30212 19800 30240
rect 19679 30209 19691 30212
rect 19633 30203 19691 30209
rect 19794 30200 19800 30212
rect 19852 30200 19858 30252
rect 20548 30240 20576 30271
rect 21542 30268 21548 30280
rect 21600 30268 21606 30320
rect 24394 30268 24400 30320
rect 24452 30317 24458 30320
rect 24452 30308 24464 30317
rect 24452 30280 24497 30308
rect 24452 30271 24464 30280
rect 24452 30268 24458 30271
rect 25774 30268 25780 30320
rect 25832 30308 25838 30320
rect 28000 30308 28028 30339
rect 28690 30311 28748 30317
rect 28690 30308 28702 30311
rect 25832 30280 27016 30308
rect 28000 30280 28702 30308
rect 25832 30268 25838 30280
rect 22186 30240 22192 30252
rect 20548 30212 22192 30240
rect 22186 30200 22192 30212
rect 22244 30200 22250 30252
rect 22281 30243 22339 30249
rect 22281 30209 22293 30243
rect 22327 30240 22339 30243
rect 22462 30240 22468 30252
rect 22327 30212 22468 30240
rect 22327 30209 22339 30212
rect 22281 30203 22339 30209
rect 22462 30200 22468 30212
rect 22520 30200 22526 30252
rect 24670 30240 24676 30252
rect 24631 30212 24676 30240
rect 24670 30200 24676 30212
rect 24728 30200 24734 30252
rect 25682 30240 25688 30252
rect 25643 30212 25688 30240
rect 25682 30200 25688 30212
rect 25740 30200 25746 30252
rect 26988 30249 27016 30280
rect 28690 30277 28702 30280
rect 28736 30277 28748 30311
rect 28690 30271 28748 30277
rect 25961 30243 26019 30249
rect 25961 30209 25973 30243
rect 26007 30209 26019 30243
rect 25961 30203 26019 30209
rect 26973 30243 27031 30249
rect 26973 30209 26985 30243
rect 27019 30209 27031 30243
rect 27154 30240 27160 30252
rect 27115 30212 27160 30240
rect 26973 30203 27031 30209
rect 19889 30175 19947 30181
rect 17880 30144 18644 30172
rect 17770 30104 17776 30116
rect 16960 30076 17776 30104
rect 13817 30067 13875 30073
rect 17770 30064 17776 30076
rect 17828 30064 17834 30116
rect 13357 30039 13415 30045
rect 13357 30005 13369 30039
rect 13403 30036 13415 30039
rect 14458 30036 14464 30048
rect 13403 30008 14464 30036
rect 13403 30005 13415 30008
rect 13357 29999 13415 30005
rect 14458 29996 14464 30008
rect 14516 29996 14522 30048
rect 16574 29996 16580 30048
rect 16632 30036 16638 30048
rect 17880 30036 17908 30144
rect 17957 30107 18015 30113
rect 17957 30073 17969 30107
rect 18003 30104 18015 30107
rect 18414 30104 18420 30116
rect 18003 30076 18420 30104
rect 18003 30073 18015 30076
rect 17957 30067 18015 30073
rect 18414 30064 18420 30076
rect 18472 30064 18478 30116
rect 18506 30036 18512 30048
rect 16632 30008 17908 30036
rect 18467 30008 18512 30036
rect 16632 29996 16638 30008
rect 18506 29996 18512 30008
rect 18564 29996 18570 30048
rect 18616 30036 18644 30144
rect 19889 30141 19901 30175
rect 19935 30172 19947 30175
rect 20714 30172 20720 30184
rect 19935 30144 20720 30172
rect 19935 30141 19947 30144
rect 19889 30135 19947 30141
rect 20714 30132 20720 30144
rect 20772 30132 20778 30184
rect 23382 30172 23388 30184
rect 22066 30144 23388 30172
rect 22066 30104 22094 30144
rect 23382 30132 23388 30144
rect 23440 30132 23446 30184
rect 25976 30172 26004 30203
rect 27154 30200 27160 30212
rect 27212 30200 27218 30252
rect 27798 30240 27804 30252
rect 27759 30212 27804 30240
rect 27798 30200 27804 30212
rect 27856 30200 27862 30252
rect 28445 30243 28503 30249
rect 28445 30209 28457 30243
rect 28491 30240 28503 30243
rect 28534 30240 28540 30252
rect 28491 30212 28540 30240
rect 28491 30209 28503 30212
rect 28445 30203 28503 30209
rect 28534 30200 28540 30212
rect 28592 30200 28598 30252
rect 32674 30240 32680 30252
rect 32635 30212 32680 30240
rect 32674 30200 32680 30212
rect 32732 30200 32738 30252
rect 33336 30249 33364 30348
rect 34146 30336 34152 30348
rect 34204 30336 34210 30388
rect 35345 30379 35403 30385
rect 35345 30345 35357 30379
rect 35391 30376 35403 30379
rect 35526 30376 35532 30388
rect 35391 30348 35532 30376
rect 35391 30345 35403 30348
rect 35345 30339 35403 30345
rect 35526 30336 35532 30348
rect 35584 30336 35590 30388
rect 33410 30268 33416 30320
rect 33468 30308 33474 30320
rect 33781 30311 33839 30317
rect 33468 30280 33513 30308
rect 33468 30268 33474 30280
rect 33781 30277 33793 30311
rect 33827 30308 33839 30311
rect 34425 30311 34483 30317
rect 34425 30308 34437 30311
rect 33827 30280 34437 30308
rect 33827 30277 33839 30280
rect 33781 30271 33839 30277
rect 34425 30277 34437 30280
rect 34471 30277 34483 30311
rect 34425 30271 34483 30277
rect 34514 30268 34520 30320
rect 34572 30308 34578 30320
rect 34572 30280 36768 30308
rect 34572 30268 34578 30280
rect 32861 30243 32919 30249
rect 32861 30209 32873 30243
rect 32907 30240 32919 30243
rect 33321 30243 33379 30249
rect 33321 30240 33333 30243
rect 32907 30212 33333 30240
rect 32907 30209 32919 30212
rect 32861 30203 32919 30209
rect 33321 30209 33333 30212
rect 33367 30209 33379 30243
rect 33321 30203 33379 30209
rect 33597 30243 33655 30249
rect 33597 30209 33609 30243
rect 33643 30209 33655 30243
rect 33597 30203 33655 30209
rect 34793 30243 34851 30249
rect 34793 30209 34805 30243
rect 34839 30240 34851 30243
rect 35342 30240 35348 30252
rect 34839 30212 35348 30240
rect 34839 30209 34851 30212
rect 34793 30203 34851 30209
rect 27065 30175 27123 30181
rect 27065 30172 27077 30175
rect 25976 30144 27077 30172
rect 27065 30141 27077 30144
rect 27111 30141 27123 30175
rect 33612 30172 33640 30203
rect 35342 30200 35348 30212
rect 35400 30200 35406 30252
rect 36446 30200 36452 30252
rect 36504 30249 36510 30252
rect 36740 30249 36768 30280
rect 37568 30280 39436 30308
rect 37568 30249 37596 30280
rect 37826 30249 37832 30252
rect 36504 30240 36516 30249
rect 36725 30243 36783 30249
rect 36504 30212 36549 30240
rect 36504 30203 36516 30212
rect 36725 30209 36737 30243
rect 36771 30240 36783 30243
rect 37553 30243 37611 30249
rect 37553 30240 37565 30243
rect 36771 30212 37565 30240
rect 36771 30209 36783 30212
rect 36725 30203 36783 30209
rect 37553 30209 37565 30212
rect 37599 30209 37611 30243
rect 37553 30203 37611 30209
rect 37820 30203 37832 30249
rect 37884 30240 37890 30252
rect 39408 30249 39436 30280
rect 39666 30249 39672 30252
rect 39393 30243 39451 30249
rect 37884 30212 37920 30240
rect 36504 30200 36510 30203
rect 37826 30200 37832 30203
rect 37884 30200 37890 30212
rect 39393 30209 39405 30243
rect 39439 30209 39451 30243
rect 39393 30203 39451 30209
rect 39660 30203 39672 30249
rect 39724 30240 39730 30252
rect 41785 30243 41843 30249
rect 39724 30212 39760 30240
rect 39666 30200 39672 30203
rect 39724 30200 39730 30212
rect 41785 30209 41797 30243
rect 41831 30240 41843 30243
rect 42150 30240 42156 30252
rect 41831 30212 42156 30240
rect 41831 30209 41843 30212
rect 41785 30203 41843 30209
rect 42150 30200 42156 30212
rect 42208 30200 42214 30252
rect 34330 30172 34336 30184
rect 33612 30144 34336 30172
rect 27065 30135 27123 30141
rect 34330 30132 34336 30144
rect 34388 30132 34394 30184
rect 19904 30076 22094 30104
rect 19904 30036 19932 30076
rect 34146 30064 34152 30116
rect 34204 30104 34210 30116
rect 34204 30076 34468 30104
rect 34204 30064 34210 30076
rect 18616 30008 19932 30036
rect 20717 30039 20775 30045
rect 20717 30005 20729 30039
rect 20763 30036 20775 30039
rect 20806 30036 20812 30048
rect 20763 30008 20812 30036
rect 20763 30005 20775 30008
rect 20717 29999 20775 30005
rect 20806 29996 20812 30008
rect 20864 29996 20870 30048
rect 20901 30039 20959 30045
rect 20901 30005 20913 30039
rect 20947 30036 20959 30039
rect 20990 30036 20996 30048
rect 20947 30008 20996 30036
rect 20947 30005 20959 30008
rect 20901 29999 20959 30005
rect 20990 29996 20996 30008
rect 21048 29996 21054 30048
rect 22278 29996 22284 30048
rect 22336 30036 22342 30048
rect 22373 30039 22431 30045
rect 22373 30036 22385 30039
rect 22336 30008 22385 30036
rect 22336 29996 22342 30008
rect 22373 30005 22385 30008
rect 22419 30005 22431 30039
rect 22373 29999 22431 30005
rect 28626 29996 28632 30048
rect 28684 30036 28690 30048
rect 29825 30039 29883 30045
rect 29825 30036 29837 30039
rect 28684 30008 29837 30036
rect 28684 29996 28690 30008
rect 29825 30005 29837 30008
rect 29871 30005 29883 30039
rect 32674 30036 32680 30048
rect 32635 30008 32680 30036
rect 29825 29999 29883 30005
rect 32674 29996 32680 30008
rect 32732 29996 32738 30048
rect 34238 30036 34244 30048
rect 34199 30008 34244 30036
rect 34238 29996 34244 30008
rect 34296 29996 34302 30048
rect 34440 30045 34468 30076
rect 38562 30064 38568 30116
rect 38620 30104 38626 30116
rect 38933 30107 38991 30113
rect 38933 30104 38945 30107
rect 38620 30076 38945 30104
rect 38620 30064 38626 30076
rect 38933 30073 38945 30076
rect 38979 30073 38991 30107
rect 38933 30067 38991 30073
rect 34425 30039 34483 30045
rect 34425 30005 34437 30039
rect 34471 30036 34483 30039
rect 37734 30036 37740 30048
rect 34471 30008 37740 30036
rect 34471 30005 34483 30008
rect 34425 29999 34483 30005
rect 37734 29996 37740 30008
rect 37792 29996 37798 30048
rect 39574 29996 39580 30048
rect 39632 30036 39638 30048
rect 40773 30039 40831 30045
rect 40773 30036 40785 30039
rect 39632 30008 40785 30036
rect 39632 29996 39638 30008
rect 40773 30005 40785 30008
rect 40819 30005 40831 30039
rect 40773 29999 40831 30005
rect 1104 29946 42872 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 42872 29946
rect 1104 29872 42872 29894
rect 8018 29792 8024 29844
rect 8076 29832 8082 29844
rect 22462 29832 22468 29844
rect 8076 29804 22468 29832
rect 8076 29792 8082 29804
rect 22462 29792 22468 29804
rect 22520 29792 22526 29844
rect 22833 29835 22891 29841
rect 22833 29801 22845 29835
rect 22879 29832 22891 29835
rect 22922 29832 22928 29844
rect 22879 29804 22928 29832
rect 22879 29801 22891 29804
rect 22833 29795 22891 29801
rect 14369 29767 14427 29773
rect 14369 29733 14381 29767
rect 14415 29764 14427 29767
rect 14918 29764 14924 29776
rect 14415 29736 14924 29764
rect 14415 29733 14427 29736
rect 14369 29727 14427 29733
rect 14918 29724 14924 29736
rect 14976 29724 14982 29776
rect 16758 29764 16764 29776
rect 15764 29736 16764 29764
rect 14458 29696 14464 29708
rect 14419 29668 14464 29696
rect 14458 29656 14464 29668
rect 14516 29656 14522 29708
rect 11701 29631 11759 29637
rect 11701 29597 11713 29631
rect 11747 29628 11759 29631
rect 14274 29628 14280 29640
rect 11747 29600 12112 29628
rect 14235 29600 14280 29628
rect 11747 29597 11759 29600
rect 11701 29591 11759 29597
rect 12084 29572 12112 29600
rect 14274 29588 14280 29600
rect 14332 29588 14338 29640
rect 14550 29588 14556 29640
rect 14608 29628 14614 29640
rect 14608 29600 14653 29628
rect 14608 29588 14614 29600
rect 14734 29588 14740 29640
rect 14792 29628 14798 29640
rect 14792 29600 14837 29628
rect 14792 29588 14798 29600
rect 14918 29588 14924 29640
rect 14976 29628 14982 29640
rect 15197 29631 15255 29637
rect 15197 29628 15209 29631
rect 14976 29600 15209 29628
rect 14976 29588 14982 29600
rect 15197 29597 15209 29600
rect 15243 29597 15255 29631
rect 15470 29628 15476 29640
rect 15431 29600 15476 29628
rect 15197 29591 15255 29597
rect 15470 29588 15476 29600
rect 15528 29588 15534 29640
rect 15764 29637 15792 29736
rect 16758 29724 16764 29736
rect 16816 29764 16822 29776
rect 17129 29767 17187 29773
rect 17129 29764 17141 29767
rect 16816 29736 17141 29764
rect 16816 29724 16822 29736
rect 17129 29733 17141 29736
rect 17175 29733 17187 29767
rect 17129 29727 17187 29733
rect 18506 29724 18512 29776
rect 18564 29764 18570 29776
rect 18564 29736 19564 29764
rect 18564 29724 18570 29736
rect 19536 29696 19564 29736
rect 19794 29724 19800 29776
rect 19852 29764 19858 29776
rect 19889 29767 19947 29773
rect 19889 29764 19901 29767
rect 19852 29736 19901 29764
rect 19852 29724 19858 29736
rect 19889 29733 19901 29736
rect 19935 29733 19947 29767
rect 19889 29727 19947 29733
rect 22370 29724 22376 29776
rect 22428 29764 22434 29776
rect 22848 29764 22876 29795
rect 22922 29792 22928 29804
rect 22980 29792 22986 29844
rect 25866 29832 25872 29844
rect 25827 29804 25872 29832
rect 25866 29792 25872 29804
rect 25924 29792 25930 29844
rect 26053 29835 26111 29841
rect 26053 29801 26065 29835
rect 26099 29832 26111 29835
rect 27062 29832 27068 29844
rect 26099 29804 27068 29832
rect 26099 29801 26111 29804
rect 26053 29795 26111 29801
rect 27062 29792 27068 29804
rect 27120 29792 27126 29844
rect 27798 29792 27804 29844
rect 27856 29832 27862 29844
rect 29549 29835 29607 29841
rect 29549 29832 29561 29835
rect 27856 29804 29561 29832
rect 27856 29792 27862 29804
rect 29549 29801 29561 29804
rect 29595 29801 29607 29835
rect 29730 29832 29736 29844
rect 29691 29804 29736 29832
rect 29549 29795 29607 29801
rect 29730 29792 29736 29804
rect 29788 29792 29794 29844
rect 30650 29832 30656 29844
rect 30392 29804 30656 29832
rect 22428 29736 22876 29764
rect 22428 29724 22434 29736
rect 23382 29724 23388 29776
rect 23440 29764 23446 29776
rect 23477 29767 23535 29773
rect 23477 29764 23489 29767
rect 23440 29736 23489 29764
rect 23440 29724 23446 29736
rect 23477 29733 23489 29736
rect 23523 29733 23535 29767
rect 30392 29764 30420 29804
rect 30650 29792 30656 29804
rect 30708 29792 30714 29844
rect 33962 29832 33968 29844
rect 33923 29804 33968 29832
rect 33962 29792 33968 29804
rect 34020 29792 34026 29844
rect 35434 29792 35440 29844
rect 35492 29832 35498 29844
rect 36081 29835 36139 29841
rect 36081 29832 36093 29835
rect 35492 29804 36093 29832
rect 35492 29792 35498 29804
rect 36081 29801 36093 29804
rect 36127 29801 36139 29835
rect 37734 29832 37740 29844
rect 37695 29804 37740 29832
rect 36081 29795 36139 29801
rect 37734 29792 37740 29804
rect 37792 29792 37798 29844
rect 39666 29792 39672 29844
rect 39724 29832 39730 29844
rect 39853 29835 39911 29841
rect 39853 29832 39865 29835
rect 39724 29804 39865 29832
rect 39724 29792 39730 29804
rect 39853 29801 39865 29804
rect 39899 29801 39911 29835
rect 39853 29795 39911 29801
rect 23477 29727 23535 29733
rect 29012 29736 30420 29764
rect 29012 29708 29040 29736
rect 19536 29668 19656 29696
rect 15749 29631 15807 29637
rect 15749 29597 15761 29631
rect 15795 29597 15807 29631
rect 15930 29628 15936 29640
rect 15891 29600 15936 29628
rect 15749 29591 15807 29597
rect 15930 29588 15936 29600
rect 15988 29588 15994 29640
rect 16206 29588 16212 29640
rect 16264 29628 16270 29640
rect 16485 29631 16543 29637
rect 16485 29628 16497 29631
rect 16264 29600 16497 29628
rect 16264 29588 16270 29600
rect 16485 29597 16497 29600
rect 16531 29597 16543 29631
rect 18506 29628 18512 29640
rect 16485 29591 16543 29597
rect 18156 29600 18512 29628
rect 11974 29569 11980 29572
rect 11968 29560 11980 29569
rect 11935 29532 11980 29560
rect 11968 29523 11980 29532
rect 11974 29520 11980 29523
rect 12032 29520 12038 29572
rect 12066 29520 12072 29572
rect 12124 29560 12130 29572
rect 18156 29560 18184 29600
rect 18506 29588 18512 29600
rect 18564 29588 18570 29640
rect 18966 29588 18972 29640
rect 19024 29628 19030 29640
rect 19242 29628 19248 29640
rect 19024 29600 19248 29628
rect 19024 29588 19030 29600
rect 19242 29588 19248 29600
rect 19300 29588 19306 29640
rect 19628 29637 19656 29668
rect 25130 29656 25136 29708
rect 25188 29696 25194 29708
rect 28442 29696 28448 29708
rect 25188 29668 28448 29696
rect 25188 29656 25194 29668
rect 28442 29656 28448 29668
rect 28500 29656 28506 29708
rect 28994 29696 29000 29708
rect 28955 29668 29000 29696
rect 28994 29656 29000 29668
rect 29052 29656 29058 29708
rect 37752 29696 37780 29792
rect 38105 29767 38163 29773
rect 38105 29733 38117 29767
rect 38151 29764 38163 29767
rect 39114 29764 39120 29776
rect 38151 29736 39120 29764
rect 38151 29733 38163 29736
rect 38105 29727 38163 29733
rect 39114 29724 39120 29736
rect 39172 29764 39178 29776
rect 40221 29767 40279 29773
rect 40221 29764 40233 29767
rect 39172 29736 40233 29764
rect 39172 29724 39178 29736
rect 40221 29733 40233 29736
rect 40267 29733 40279 29767
rect 40221 29727 40279 29733
rect 38657 29699 38715 29705
rect 38657 29696 38669 29699
rect 37752 29668 38669 29696
rect 38657 29665 38669 29668
rect 38703 29665 38715 29699
rect 38657 29659 38715 29665
rect 38841 29699 38899 29705
rect 38841 29665 38853 29699
rect 38887 29696 38899 29699
rect 38887 29668 40080 29696
rect 38887 29665 38899 29668
rect 38841 29659 38899 29665
rect 19429 29631 19487 29637
rect 19429 29628 19441 29631
rect 19352 29600 19441 29628
rect 12124 29532 18184 29560
rect 12124 29520 12130 29532
rect 18230 29520 18236 29572
rect 18288 29569 18294 29572
rect 18288 29560 18300 29569
rect 18288 29532 18333 29560
rect 18288 29523 18300 29532
rect 18288 29520 18294 29523
rect 18414 29520 18420 29572
rect 18472 29560 18478 29572
rect 19352 29560 19380 29600
rect 19429 29597 19441 29600
rect 19475 29597 19487 29631
rect 19429 29591 19487 29597
rect 19521 29631 19579 29637
rect 19521 29597 19533 29631
rect 19567 29597 19579 29631
rect 19521 29591 19579 29597
rect 19613 29631 19671 29637
rect 19613 29597 19625 29631
rect 19659 29597 19671 29631
rect 20438 29628 20444 29640
rect 20399 29600 20444 29628
rect 19613 29591 19671 29597
rect 18472 29532 19380 29560
rect 19536 29560 19564 29591
rect 20438 29588 20444 29600
rect 20496 29588 20502 29640
rect 22925 29631 22983 29637
rect 22925 29597 22937 29631
rect 22971 29628 22983 29631
rect 28721 29631 28779 29637
rect 22971 29600 25728 29628
rect 22971 29597 22983 29600
rect 22925 29591 22983 29597
rect 20530 29560 20536 29572
rect 19536 29532 20536 29560
rect 18472 29520 18478 29532
rect 20530 29520 20536 29532
rect 20588 29520 20594 29572
rect 20708 29563 20766 29569
rect 20708 29529 20720 29563
rect 20754 29560 20766 29563
rect 20806 29560 20812 29572
rect 20754 29532 20812 29560
rect 20754 29529 20766 29532
rect 20708 29523 20766 29529
rect 20806 29520 20812 29532
rect 20864 29520 20870 29572
rect 23661 29563 23719 29569
rect 23661 29529 23673 29563
rect 23707 29560 23719 29563
rect 23842 29560 23848 29572
rect 23707 29532 23848 29560
rect 23707 29529 23719 29532
rect 23661 29523 23719 29529
rect 23842 29520 23848 29532
rect 23900 29520 23906 29572
rect 25130 29560 25136 29572
rect 25091 29532 25136 29560
rect 25130 29520 25136 29532
rect 25188 29520 25194 29572
rect 25700 29569 25728 29600
rect 28721 29597 28733 29631
rect 28767 29597 28779 29631
rect 30374 29628 30380 29640
rect 30335 29600 30380 29628
rect 28721 29591 28779 29597
rect 25685 29563 25743 29569
rect 25685 29529 25697 29563
rect 25731 29560 25743 29563
rect 25774 29560 25780 29572
rect 25731 29532 25780 29560
rect 25731 29529 25743 29532
rect 25685 29523 25743 29529
rect 25774 29520 25780 29532
rect 25832 29560 25838 29572
rect 28736 29560 28764 29591
rect 30374 29588 30380 29600
rect 30432 29628 30438 29640
rect 32585 29631 32643 29637
rect 32585 29628 32597 29631
rect 30432 29600 32597 29628
rect 30432 29588 30438 29600
rect 32585 29597 32597 29600
rect 32631 29597 32643 29631
rect 32585 29591 32643 29597
rect 32674 29588 32680 29640
rect 32732 29628 32738 29640
rect 32841 29631 32899 29637
rect 32841 29628 32853 29631
rect 32732 29600 32853 29628
rect 32732 29588 32738 29600
rect 32841 29597 32853 29600
rect 32887 29597 32899 29631
rect 34698 29628 34704 29640
rect 34659 29600 34704 29628
rect 32841 29591 32899 29597
rect 34698 29588 34704 29600
rect 34756 29588 34762 29640
rect 39114 29628 39120 29640
rect 39075 29600 39120 29628
rect 39114 29588 39120 29600
rect 39172 29588 39178 29640
rect 40052 29637 40080 29668
rect 40037 29631 40095 29637
rect 40037 29597 40049 29631
rect 40083 29597 40095 29631
rect 40037 29591 40095 29597
rect 40313 29631 40371 29637
rect 40313 29597 40325 29631
rect 40359 29597 40371 29631
rect 40313 29591 40371 29597
rect 29917 29563 29975 29569
rect 29917 29560 29929 29563
rect 25832 29532 29929 29560
rect 25832 29520 25838 29532
rect 29917 29529 29929 29532
rect 29963 29529 29975 29563
rect 29917 29523 29975 29529
rect 30006 29520 30012 29572
rect 30064 29560 30070 29572
rect 30622 29563 30680 29569
rect 30622 29560 30634 29563
rect 30064 29532 30634 29560
rect 30064 29520 30070 29532
rect 30622 29529 30634 29532
rect 30668 29529 30680 29563
rect 30622 29523 30680 29529
rect 34790 29520 34796 29572
rect 34848 29560 34854 29572
rect 34946 29563 35004 29569
rect 34946 29560 34958 29563
rect 34848 29532 34958 29560
rect 34848 29520 34854 29532
rect 34946 29529 34958 29532
rect 34992 29529 35004 29563
rect 34946 29523 35004 29529
rect 37737 29563 37795 29569
rect 37737 29529 37749 29563
rect 37783 29560 37795 29563
rect 37918 29560 37924 29572
rect 37783 29532 37924 29560
rect 37783 29529 37795 29532
rect 37737 29523 37795 29529
rect 37918 29520 37924 29532
rect 37976 29520 37982 29572
rect 39025 29563 39083 29569
rect 39025 29529 39037 29563
rect 39071 29560 39083 29563
rect 39482 29560 39488 29572
rect 39071 29532 39488 29560
rect 39071 29529 39083 29532
rect 39025 29523 39083 29529
rect 39482 29520 39488 29532
rect 39540 29560 39546 29572
rect 40328 29560 40356 29591
rect 42058 29560 42064 29572
rect 39540 29532 40356 29560
rect 42019 29532 42064 29560
rect 39540 29520 39546 29532
rect 42058 29520 42064 29532
rect 42116 29520 42122 29572
rect 13078 29492 13084 29504
rect 13039 29464 13084 29492
rect 13078 29452 13084 29464
rect 13136 29452 13142 29504
rect 14090 29492 14096 29504
rect 14051 29464 14096 29492
rect 14090 29452 14096 29464
rect 14148 29452 14154 29504
rect 15286 29492 15292 29504
rect 15247 29464 15292 29492
rect 15286 29452 15292 29464
rect 15344 29452 15350 29504
rect 16577 29495 16635 29501
rect 16577 29461 16589 29495
rect 16623 29492 16635 29495
rect 17126 29492 17132 29504
rect 16623 29464 17132 29492
rect 16623 29461 16635 29464
rect 16577 29455 16635 29461
rect 17126 29452 17132 29464
rect 17184 29452 17190 29504
rect 20622 29452 20628 29504
rect 20680 29492 20686 29504
rect 21821 29495 21879 29501
rect 21821 29492 21833 29495
rect 20680 29464 21833 29492
rect 20680 29452 20686 29464
rect 21821 29461 21833 29464
rect 21867 29461 21879 29495
rect 21821 29455 21879 29461
rect 24857 29495 24915 29501
rect 24857 29461 24869 29495
rect 24903 29492 24915 29495
rect 24946 29492 24952 29504
rect 24903 29464 24952 29492
rect 24903 29461 24915 29464
rect 24857 29455 24915 29461
rect 24946 29452 24952 29464
rect 25004 29492 25010 29504
rect 25222 29492 25228 29504
rect 25004 29464 25228 29492
rect 25004 29452 25010 29464
rect 25222 29452 25228 29464
rect 25280 29452 25286 29504
rect 25498 29452 25504 29504
rect 25556 29492 25562 29504
rect 25885 29495 25943 29501
rect 25885 29492 25897 29495
rect 25556 29464 25897 29492
rect 25556 29452 25562 29464
rect 25885 29461 25897 29464
rect 25931 29461 25943 29495
rect 25885 29455 25943 29461
rect 28994 29452 29000 29504
rect 29052 29492 29058 29504
rect 29707 29495 29765 29501
rect 29707 29492 29719 29495
rect 29052 29464 29719 29492
rect 29052 29452 29058 29464
rect 29707 29461 29719 29464
rect 29753 29461 29765 29495
rect 29707 29455 29765 29461
rect 30742 29452 30748 29504
rect 30800 29492 30806 29504
rect 31757 29495 31815 29501
rect 31757 29492 31769 29495
rect 30800 29464 31769 29492
rect 30800 29452 30806 29464
rect 31757 29461 31769 29464
rect 31803 29461 31815 29495
rect 37550 29492 37556 29504
rect 37511 29464 37556 29492
rect 31757 29455 31815 29461
rect 37550 29452 37556 29464
rect 37608 29452 37614 29504
rect 41966 29492 41972 29504
rect 41927 29464 41972 29492
rect 41966 29452 41972 29464
rect 42024 29452 42030 29504
rect 1104 29402 42872 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 42872 29402
rect 1104 29328 42872 29350
rect 15746 29288 15752 29300
rect 15707 29260 15752 29288
rect 15746 29248 15752 29260
rect 15804 29248 15810 29300
rect 15917 29291 15975 29297
rect 15917 29257 15929 29291
rect 15963 29288 15975 29291
rect 16206 29288 16212 29300
rect 15963 29260 16212 29288
rect 15963 29257 15975 29260
rect 15917 29251 15975 29257
rect 16206 29248 16212 29260
rect 16264 29248 16270 29300
rect 20806 29288 20812 29300
rect 20767 29260 20812 29288
rect 20806 29248 20812 29260
rect 20864 29248 20870 29300
rect 23569 29291 23627 29297
rect 23569 29288 23581 29291
rect 22572 29260 23581 29288
rect 12336 29223 12394 29229
rect 12336 29189 12348 29223
rect 12382 29220 12394 29223
rect 14090 29220 14096 29232
rect 12382 29192 14096 29220
rect 12382 29189 12394 29192
rect 12336 29183 12394 29189
rect 14090 29180 14096 29192
rect 14148 29180 14154 29232
rect 16117 29223 16175 29229
rect 16117 29189 16129 29223
rect 16163 29220 16175 29223
rect 16482 29220 16488 29232
rect 16163 29192 16488 29220
rect 16163 29189 16175 29192
rect 16117 29183 16175 29189
rect 16482 29180 16488 29192
rect 16540 29220 16546 29232
rect 17218 29220 17224 29232
rect 16540 29192 17224 29220
rect 16540 29180 16546 29192
rect 12066 29152 12072 29164
rect 12027 29124 12072 29152
rect 12066 29112 12072 29124
rect 12124 29112 12130 29164
rect 13078 29112 13084 29164
rect 13136 29152 13142 29164
rect 14829 29155 14887 29161
rect 14829 29152 14841 29155
rect 13136 29124 14841 29152
rect 13136 29112 13142 29124
rect 14829 29121 14841 29124
rect 14875 29152 14887 29155
rect 15470 29152 15476 29164
rect 14875 29124 15476 29152
rect 14875 29121 14887 29124
rect 14829 29115 14887 29121
rect 15470 29112 15476 29124
rect 15528 29112 15534 29164
rect 16758 29152 16764 29164
rect 16719 29124 16764 29152
rect 16758 29112 16764 29124
rect 16816 29112 16822 29164
rect 17052 29161 17080 29192
rect 17218 29180 17224 29192
rect 17276 29180 17282 29232
rect 18506 29180 18512 29232
rect 18564 29220 18570 29232
rect 18690 29220 18696 29232
rect 18564 29192 18696 29220
rect 18564 29180 18570 29192
rect 18690 29180 18696 29192
rect 18748 29220 18754 29232
rect 19426 29220 19432 29232
rect 18748 29192 19432 29220
rect 18748 29180 18754 29192
rect 19426 29180 19432 29192
rect 19484 29220 19490 29232
rect 20438 29220 20444 29232
rect 19484 29192 20444 29220
rect 19484 29180 19490 29192
rect 20438 29180 20444 29192
rect 20496 29180 20502 29232
rect 17037 29155 17095 29161
rect 17037 29121 17049 29155
rect 17083 29121 17095 29155
rect 17037 29115 17095 29121
rect 19613 29155 19671 29161
rect 19613 29121 19625 29155
rect 19659 29152 19671 29155
rect 20898 29152 20904 29164
rect 19659 29124 20904 29152
rect 19659 29121 19671 29124
rect 19613 29115 19671 29121
rect 20898 29112 20904 29124
rect 20956 29112 20962 29164
rect 20990 29112 20996 29164
rect 21048 29152 21054 29164
rect 22572 29161 22600 29260
rect 23569 29257 23581 29260
rect 23615 29257 23627 29291
rect 26602 29288 26608 29300
rect 23569 29251 23627 29257
rect 23676 29260 26608 29288
rect 23382 29220 23388 29232
rect 22756 29192 23388 29220
rect 22756 29161 22784 29192
rect 23382 29180 23388 29192
rect 23440 29180 23446 29232
rect 23676 29161 23704 29260
rect 26602 29248 26608 29260
rect 26660 29248 26666 29300
rect 28721 29291 28779 29297
rect 28721 29257 28733 29291
rect 28767 29288 28779 29291
rect 29730 29288 29736 29300
rect 28767 29260 29736 29288
rect 28767 29257 28779 29260
rect 28721 29251 28779 29257
rect 29730 29248 29736 29260
rect 29788 29248 29794 29300
rect 29825 29291 29883 29297
rect 29825 29257 29837 29291
rect 29871 29288 29883 29291
rect 30006 29288 30012 29300
rect 29871 29260 30012 29288
rect 29871 29257 29883 29260
rect 29825 29251 29883 29257
rect 30006 29248 30012 29260
rect 30064 29248 30070 29300
rect 34701 29291 34759 29297
rect 34701 29257 34713 29291
rect 34747 29288 34759 29291
rect 34790 29288 34796 29300
rect 34747 29260 34796 29288
rect 34747 29257 34759 29260
rect 34701 29251 34759 29257
rect 34790 29248 34796 29260
rect 34848 29248 34854 29300
rect 37826 29288 37832 29300
rect 37787 29260 37832 29288
rect 37826 29248 37832 29260
rect 37884 29248 37890 29300
rect 24121 29223 24179 29229
rect 24121 29189 24133 29223
rect 24167 29189 24179 29223
rect 24121 29183 24179 29189
rect 24337 29223 24395 29229
rect 24337 29189 24349 29223
rect 24383 29220 24395 29223
rect 24854 29220 24860 29232
rect 24383 29192 24860 29220
rect 24383 29189 24395 29192
rect 24337 29183 24395 29189
rect 22557 29155 22615 29161
rect 21048 29124 21093 29152
rect 21048 29112 21054 29124
rect 22557 29121 22569 29155
rect 22603 29121 22615 29155
rect 22557 29115 22615 29121
rect 22740 29155 22798 29161
rect 22740 29121 22752 29155
rect 22786 29121 22798 29155
rect 22740 29115 22798 29121
rect 23661 29155 23719 29161
rect 23661 29121 23673 29155
rect 23707 29121 23719 29155
rect 24136 29152 24164 29183
rect 24854 29180 24860 29192
rect 24912 29180 24918 29232
rect 25774 29180 25780 29232
rect 25832 29220 25838 29232
rect 25869 29223 25927 29229
rect 25869 29220 25881 29223
rect 25832 29192 25881 29220
rect 25832 29180 25838 29192
rect 25869 29189 25881 29192
rect 25915 29189 25927 29223
rect 25869 29183 25927 29189
rect 25958 29180 25964 29232
rect 26016 29220 26022 29232
rect 26069 29223 26127 29229
rect 26069 29220 26081 29223
rect 26016 29192 26081 29220
rect 26016 29180 26022 29192
rect 26069 29189 26081 29192
rect 26115 29189 26127 29223
rect 26069 29183 26127 29189
rect 28368 29192 29592 29220
rect 25792 29152 25820 29180
rect 28368 29164 28396 29192
rect 26973 29155 27031 29161
rect 26973 29152 26985 29155
rect 24136 29124 25820 29152
rect 26252 29124 26985 29152
rect 23661 29115 23719 29121
rect 13998 29044 14004 29096
rect 14056 29084 14062 29096
rect 14553 29087 14611 29093
rect 14553 29084 14565 29087
rect 14056 29056 14565 29084
rect 14056 29044 14062 29056
rect 14553 29053 14565 29056
rect 14599 29053 14611 29087
rect 14553 29047 14611 29053
rect 22278 29044 22284 29096
rect 22336 29084 22342 29096
rect 22649 29087 22707 29093
rect 22649 29084 22661 29087
rect 22336 29056 22661 29084
rect 22336 29044 22342 29056
rect 22649 29053 22661 29056
rect 22695 29053 22707 29087
rect 22649 29047 22707 29053
rect 22833 29087 22891 29093
rect 22833 29053 22845 29087
rect 22879 29053 22891 29087
rect 22833 29047 22891 29053
rect 14734 28976 14740 29028
rect 14792 29016 14798 29028
rect 17218 29016 17224 29028
rect 14792 28988 17224 29016
rect 14792 28976 14798 28988
rect 17218 28976 17224 28988
rect 17276 29016 17282 29028
rect 22370 29016 22376 29028
rect 17276 28988 22376 29016
rect 17276 28976 17282 28988
rect 22370 28976 22376 28988
rect 22428 28976 22434 29028
rect 22554 28976 22560 29028
rect 22612 29016 22618 29028
rect 22848 29016 22876 29047
rect 22612 28988 22876 29016
rect 23017 29019 23075 29025
rect 22612 28976 22618 28988
rect 23017 28985 23029 29019
rect 23063 29016 23075 29019
rect 24489 29019 24547 29025
rect 23063 28988 24348 29016
rect 23063 28985 23075 28988
rect 23017 28979 23075 28985
rect 24320 28960 24348 28988
rect 24489 28985 24501 29019
rect 24535 29016 24547 29019
rect 24578 29016 24584 29028
rect 24535 28988 24584 29016
rect 24535 28985 24547 28988
rect 24489 28979 24547 28985
rect 24578 28976 24584 28988
rect 24636 28976 24642 29028
rect 26252 29025 26280 29124
rect 26973 29121 26985 29124
rect 27019 29121 27031 29155
rect 26973 29115 27031 29121
rect 28261 29155 28319 29161
rect 28261 29121 28273 29155
rect 28307 29121 28319 29155
rect 28261 29115 28319 29121
rect 28276 29084 28304 29115
rect 28350 29112 28356 29164
rect 28408 29152 28414 29164
rect 28408 29124 28453 29152
rect 28408 29112 28414 29124
rect 28534 29112 28540 29164
rect 28592 29152 28598 29164
rect 29178 29152 29184 29164
rect 28592 29124 28637 29152
rect 29139 29124 29184 29152
rect 28592 29112 28598 29124
rect 29178 29112 29184 29124
rect 29236 29112 29242 29164
rect 29362 29152 29368 29164
rect 29323 29124 29368 29152
rect 29362 29112 29368 29124
rect 29420 29112 29426 29164
rect 29564 29161 29592 29192
rect 29457 29155 29515 29161
rect 29457 29121 29469 29155
rect 29503 29121 29515 29155
rect 29457 29115 29515 29121
rect 29549 29155 29607 29161
rect 29549 29121 29561 29155
rect 29595 29152 29607 29155
rect 30742 29152 30748 29164
rect 29595 29124 29684 29152
rect 30703 29124 30748 29152
rect 29595 29121 29607 29124
rect 29549 29115 29607 29121
rect 29086 29084 29092 29096
rect 28276 29056 29092 29084
rect 29086 29044 29092 29056
rect 29144 29084 29150 29096
rect 29472 29084 29500 29115
rect 29144 29056 29500 29084
rect 29656 29084 29684 29124
rect 30742 29112 30748 29124
rect 30800 29112 30806 29164
rect 34238 29112 34244 29164
rect 34296 29152 34302 29164
rect 34517 29155 34575 29161
rect 34517 29152 34529 29155
rect 34296 29124 34529 29152
rect 34296 29112 34302 29124
rect 34517 29121 34529 29124
rect 34563 29121 34575 29155
rect 34517 29115 34575 29121
rect 37550 29112 37556 29164
rect 37608 29152 37614 29164
rect 38013 29155 38071 29161
rect 38013 29152 38025 29155
rect 37608 29124 38025 29152
rect 37608 29112 37614 29124
rect 38013 29121 38025 29124
rect 38059 29121 38071 29155
rect 38013 29115 38071 29121
rect 31021 29087 31079 29093
rect 31021 29084 31033 29087
rect 29656 29056 31033 29084
rect 29144 29044 29150 29056
rect 31021 29053 31033 29056
rect 31067 29053 31079 29087
rect 31021 29047 31079 29053
rect 26237 29019 26295 29025
rect 26237 28985 26249 29019
rect 26283 28985 26295 29019
rect 26237 28979 26295 28985
rect 1670 28948 1676 28960
rect 1631 28920 1676 28948
rect 1670 28908 1676 28920
rect 1728 28908 1734 28960
rect 13446 28948 13452 28960
rect 13407 28920 13452 28948
rect 13446 28908 13452 28920
rect 13504 28908 13510 28960
rect 15838 28908 15844 28960
rect 15896 28948 15902 28960
rect 15933 28951 15991 28957
rect 15933 28948 15945 28951
rect 15896 28920 15945 28948
rect 15896 28908 15902 28920
rect 15933 28917 15945 28920
rect 15979 28917 15991 28951
rect 24302 28948 24308 28960
rect 24215 28920 24308 28948
rect 15933 28911 15991 28917
rect 24302 28908 24308 28920
rect 24360 28908 24366 28960
rect 26053 28951 26111 28957
rect 26053 28917 26065 28951
rect 26099 28948 26111 28951
rect 26326 28948 26332 28960
rect 26099 28920 26332 28948
rect 26099 28917 26111 28920
rect 26053 28911 26111 28917
rect 26326 28908 26332 28920
rect 26384 28908 26390 28960
rect 27154 28948 27160 28960
rect 27115 28920 27160 28948
rect 27154 28908 27160 28920
rect 27212 28908 27218 28960
rect 41782 28948 41788 28960
rect 41743 28920 41788 28948
rect 41782 28908 41788 28920
rect 41840 28908 41846 28960
rect 1104 28858 42872 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 42872 28858
rect 1104 28784 42872 28806
rect 14550 28704 14556 28756
rect 14608 28744 14614 28756
rect 14645 28747 14703 28753
rect 14645 28744 14657 28747
rect 14608 28716 14657 28744
rect 14608 28704 14614 28716
rect 14645 28713 14657 28716
rect 14691 28713 14703 28747
rect 14645 28707 14703 28713
rect 20898 28704 20904 28756
rect 20956 28744 20962 28756
rect 21726 28744 21732 28756
rect 20956 28716 21732 28744
rect 20956 28704 20962 28716
rect 21726 28704 21732 28716
rect 21784 28704 21790 28756
rect 22646 28744 22652 28756
rect 22066 28716 22652 28744
rect 14918 28676 14924 28688
rect 14200 28648 14924 28676
rect 1397 28611 1455 28617
rect 1397 28577 1409 28611
rect 1443 28608 1455 28611
rect 1670 28608 1676 28620
rect 1443 28580 1676 28608
rect 1443 28577 1455 28580
rect 1397 28571 1455 28577
rect 1670 28568 1676 28580
rect 1728 28568 1734 28620
rect 2774 28608 2780 28620
rect 2735 28580 2780 28608
rect 2774 28568 2780 28580
rect 2832 28568 2838 28620
rect 13446 28568 13452 28620
rect 13504 28608 13510 28620
rect 14200 28617 14228 28648
rect 14918 28636 14924 28648
rect 14976 28636 14982 28688
rect 14185 28611 14243 28617
rect 14185 28608 14197 28611
rect 13504 28580 14197 28608
rect 13504 28568 13510 28580
rect 13556 28549 13584 28580
rect 14185 28577 14197 28580
rect 14231 28577 14243 28611
rect 14366 28608 14372 28620
rect 14327 28580 14372 28608
rect 14185 28571 14243 28577
rect 14366 28568 14372 28580
rect 14424 28568 14430 28620
rect 14461 28611 14519 28617
rect 14461 28577 14473 28611
rect 14507 28608 14519 28611
rect 15746 28608 15752 28620
rect 14507 28580 15752 28608
rect 14507 28577 14519 28580
rect 14461 28571 14519 28577
rect 15746 28568 15752 28580
rect 15804 28568 15810 28620
rect 16390 28568 16396 28620
rect 16448 28608 16454 28620
rect 16448 28580 16620 28608
rect 16448 28568 16454 28580
rect 13541 28543 13599 28549
rect 13541 28509 13553 28543
rect 13587 28509 13599 28543
rect 13541 28503 13599 28509
rect 13998 28500 14004 28552
rect 14056 28540 14062 28552
rect 14277 28543 14335 28549
rect 14277 28540 14289 28543
rect 14056 28512 14289 28540
rect 14056 28500 14062 28512
rect 14277 28509 14289 28512
rect 14323 28509 14335 28543
rect 14277 28503 14335 28509
rect 15838 28500 15844 28552
rect 15896 28540 15902 28552
rect 16592 28549 16620 28580
rect 17236 28580 17632 28608
rect 16209 28543 16267 28549
rect 16209 28540 16221 28543
rect 15896 28512 16221 28540
rect 15896 28500 15902 28512
rect 16209 28509 16221 28512
rect 16255 28509 16267 28543
rect 16209 28503 16267 28509
rect 16577 28543 16635 28549
rect 16577 28509 16589 28543
rect 16623 28509 16635 28543
rect 16577 28503 16635 28509
rect 16942 28500 16948 28552
rect 17000 28540 17006 28552
rect 17236 28549 17264 28580
rect 17221 28543 17279 28549
rect 17221 28540 17233 28543
rect 17000 28512 17233 28540
rect 17000 28500 17006 28512
rect 17221 28509 17233 28512
rect 17267 28509 17279 28543
rect 17402 28540 17408 28552
rect 17363 28512 17408 28540
rect 17221 28503 17279 28509
rect 17402 28500 17408 28512
rect 17460 28500 17466 28552
rect 17604 28540 17632 28580
rect 19426 28568 19432 28620
rect 19484 28608 19490 28620
rect 19613 28611 19671 28617
rect 19613 28608 19625 28611
rect 19484 28580 19625 28608
rect 19484 28568 19490 28580
rect 19613 28577 19625 28580
rect 19659 28577 19671 28611
rect 19613 28571 19671 28577
rect 21637 28543 21695 28549
rect 17604 28512 20392 28540
rect 1581 28475 1639 28481
rect 1581 28441 1593 28475
rect 1627 28472 1639 28475
rect 2130 28472 2136 28484
rect 1627 28444 2136 28472
rect 1627 28441 1639 28444
rect 1581 28435 1639 28441
rect 2130 28432 2136 28444
rect 2188 28432 2194 28484
rect 15930 28432 15936 28484
rect 15988 28472 15994 28484
rect 16393 28475 16451 28481
rect 16393 28472 16405 28475
rect 15988 28444 16405 28472
rect 15988 28432 15994 28444
rect 16393 28441 16405 28444
rect 16439 28441 16451 28475
rect 16393 28435 16451 28441
rect 16482 28432 16488 28484
rect 16540 28472 16546 28484
rect 19880 28475 19938 28481
rect 16540 28444 16585 28472
rect 16540 28432 16546 28444
rect 19880 28441 19892 28475
rect 19926 28472 19938 28475
rect 20254 28472 20260 28484
rect 19926 28444 20260 28472
rect 19926 28441 19938 28444
rect 19880 28435 19938 28441
rect 20254 28432 20260 28444
rect 20312 28432 20318 28484
rect 20364 28472 20392 28512
rect 21637 28509 21649 28543
rect 21683 28540 21695 28543
rect 22066 28540 22094 28716
rect 22646 28704 22652 28716
rect 22704 28744 22710 28756
rect 26878 28744 26884 28756
rect 22704 28716 26884 28744
rect 22704 28704 22710 28716
rect 26878 28704 26884 28716
rect 26936 28744 26942 28756
rect 31662 28744 31668 28756
rect 26936 28716 31668 28744
rect 26936 28704 26942 28716
rect 31662 28704 31668 28716
rect 31720 28704 31726 28756
rect 22554 28636 22560 28688
rect 22612 28676 22618 28688
rect 23477 28679 23535 28685
rect 22612 28648 22692 28676
rect 22612 28636 22618 28648
rect 22462 28608 22468 28620
rect 22423 28580 22468 28608
rect 22462 28568 22468 28580
rect 22520 28568 22526 28620
rect 22664 28617 22692 28648
rect 23477 28645 23489 28679
rect 23523 28676 23535 28679
rect 23658 28676 23664 28688
rect 23523 28648 23664 28676
rect 23523 28645 23535 28648
rect 23477 28639 23535 28645
rect 23658 28636 23664 28648
rect 23716 28636 23722 28688
rect 24854 28676 24860 28688
rect 24815 28648 24860 28676
rect 24854 28636 24860 28648
rect 24912 28636 24918 28688
rect 28810 28676 28816 28688
rect 27816 28648 28816 28676
rect 22649 28611 22707 28617
rect 22649 28577 22661 28611
rect 22695 28577 22707 28611
rect 22649 28571 22707 28577
rect 25317 28611 25375 28617
rect 25317 28577 25329 28611
rect 25363 28608 25375 28611
rect 25958 28608 25964 28620
rect 25363 28580 25964 28608
rect 25363 28577 25375 28580
rect 25317 28571 25375 28577
rect 25958 28568 25964 28580
rect 26016 28568 26022 28620
rect 22370 28540 22376 28552
rect 21683 28512 22094 28540
rect 22331 28512 22376 28540
rect 21683 28509 21695 28512
rect 21637 28503 21695 28509
rect 22370 28500 22376 28512
rect 22428 28500 22434 28552
rect 22557 28543 22615 28549
rect 22557 28509 22569 28543
rect 22603 28540 22615 28543
rect 23293 28543 23351 28549
rect 23293 28540 23305 28543
rect 22603 28512 23305 28540
rect 22603 28509 22615 28512
rect 22557 28503 22615 28509
rect 23293 28509 23305 28512
rect 23339 28540 23351 28543
rect 23842 28540 23848 28552
rect 23339 28512 23848 28540
rect 23339 28509 23351 28512
rect 23293 28503 23351 28509
rect 23842 28500 23848 28512
rect 23900 28500 23906 28552
rect 25225 28543 25283 28549
rect 25225 28509 25237 28543
rect 25271 28540 25283 28543
rect 26234 28540 26240 28552
rect 25271 28512 26240 28540
rect 25271 28509 25283 28512
rect 25225 28503 25283 28509
rect 26234 28500 26240 28512
rect 26292 28500 26298 28552
rect 26993 28543 27051 28549
rect 26993 28509 27005 28543
rect 27039 28540 27051 28543
rect 27154 28540 27160 28552
rect 27039 28512 27160 28540
rect 27039 28509 27051 28512
rect 26993 28503 27051 28509
rect 27154 28500 27160 28512
rect 27212 28500 27218 28552
rect 27816 28549 27844 28648
rect 28810 28636 28816 28648
rect 28868 28636 28874 28688
rect 28905 28679 28963 28685
rect 28905 28645 28917 28679
rect 28951 28676 28963 28679
rect 29362 28676 29368 28688
rect 28951 28648 29368 28676
rect 28951 28645 28963 28648
rect 28905 28639 28963 28645
rect 29362 28636 29368 28648
rect 29420 28636 29426 28688
rect 28077 28611 28135 28617
rect 28077 28577 28089 28611
rect 28123 28608 28135 28611
rect 41322 28608 41328 28620
rect 28123 28597 28856 28608
rect 28123 28580 28948 28597
rect 41283 28580 41328 28608
rect 28123 28577 28135 28580
rect 28077 28571 28135 28577
rect 28828 28569 28948 28580
rect 27249 28543 27307 28549
rect 27249 28509 27261 28543
rect 27295 28509 27307 28543
rect 27249 28503 27307 28509
rect 27801 28543 27859 28549
rect 27801 28509 27813 28543
rect 27847 28509 27859 28543
rect 27801 28503 27859 28509
rect 23658 28472 23664 28484
rect 20364 28444 23664 28472
rect 23658 28432 23664 28444
rect 23716 28432 23722 28484
rect 27264 28472 27292 28503
rect 27890 28500 27896 28552
rect 27948 28540 27954 28552
rect 27948 28512 27993 28540
rect 27948 28500 27954 28512
rect 28350 28500 28356 28552
rect 28408 28540 28414 28552
rect 28537 28543 28595 28549
rect 28537 28540 28549 28543
rect 28408 28512 28549 28540
rect 28408 28500 28414 28512
rect 28537 28509 28549 28512
rect 28583 28509 28595 28543
rect 28537 28503 28595 28509
rect 28626 28500 28632 28552
rect 28684 28549 28690 28552
rect 28684 28543 28733 28549
rect 28684 28509 28687 28543
rect 28721 28509 28733 28543
rect 28920 28540 28948 28569
rect 41322 28568 41328 28580
rect 41380 28568 41386 28620
rect 41782 28568 41788 28620
rect 41840 28608 41846 28620
rect 42153 28611 42211 28617
rect 42153 28608 42165 28611
rect 41840 28580 42165 28608
rect 41840 28568 41846 28580
rect 42153 28577 42165 28580
rect 42199 28577 42211 28611
rect 42153 28571 42211 28577
rect 28997 28543 29055 28549
rect 28997 28540 29009 28543
rect 28920 28512 29009 28540
rect 28684 28503 28733 28509
rect 28997 28509 29009 28512
rect 29043 28540 29055 28543
rect 29178 28540 29184 28552
rect 29043 28512 29184 28540
rect 29043 28509 29055 28512
rect 28997 28503 29055 28509
rect 28684 28500 28690 28503
rect 29178 28500 29184 28512
rect 29236 28540 29242 28552
rect 29549 28543 29607 28549
rect 29549 28540 29561 28543
rect 29236 28512 29561 28540
rect 29236 28500 29242 28512
rect 29549 28509 29561 28512
rect 29595 28509 29607 28543
rect 29549 28503 29607 28509
rect 29638 28500 29644 28552
rect 29696 28540 29702 28552
rect 29733 28543 29791 28549
rect 29733 28540 29745 28543
rect 29696 28512 29745 28540
rect 29696 28500 29702 28512
rect 29733 28509 29745 28512
rect 29779 28509 29791 28543
rect 29733 28503 29791 28509
rect 30374 28500 30380 28552
rect 30432 28540 30438 28552
rect 30561 28543 30619 28549
rect 30561 28540 30573 28543
rect 30432 28512 30573 28540
rect 30432 28500 30438 28512
rect 30561 28509 30573 28512
rect 30607 28509 30619 28543
rect 30561 28503 30619 28509
rect 30392 28472 30420 28500
rect 27264 28444 30420 28472
rect 30466 28432 30472 28484
rect 30524 28472 30530 28484
rect 30806 28475 30864 28481
rect 30806 28472 30818 28475
rect 30524 28444 30818 28472
rect 30524 28432 30530 28444
rect 30806 28441 30818 28444
rect 30852 28441 30864 28475
rect 30806 28435 30864 28441
rect 41414 28432 41420 28484
rect 41472 28472 41478 28484
rect 41969 28475 42027 28481
rect 41969 28472 41981 28475
rect 41472 28444 41981 28472
rect 41472 28432 41478 28444
rect 41969 28441 41981 28444
rect 42015 28441 42027 28475
rect 41969 28435 42027 28441
rect 13449 28407 13507 28413
rect 13449 28373 13461 28407
rect 13495 28404 13507 28407
rect 14274 28404 14280 28416
rect 13495 28376 14280 28404
rect 13495 28373 13507 28376
rect 13449 28367 13507 28373
rect 14274 28364 14280 28376
rect 14332 28404 14338 28416
rect 14550 28404 14556 28416
rect 14332 28376 14556 28404
rect 14332 28364 14338 28376
rect 14550 28364 14556 28376
rect 14608 28364 14614 28416
rect 16761 28407 16819 28413
rect 16761 28373 16773 28407
rect 16807 28404 16819 28407
rect 17310 28404 17316 28416
rect 16807 28376 17316 28404
rect 16807 28373 16819 28376
rect 16761 28367 16819 28373
rect 17310 28364 17316 28376
rect 17368 28364 17374 28416
rect 17405 28407 17463 28413
rect 17405 28373 17417 28407
rect 17451 28404 17463 28407
rect 18230 28404 18236 28416
rect 17451 28376 18236 28404
rect 17451 28373 17463 28376
rect 17405 28367 17463 28373
rect 18230 28364 18236 28376
rect 18288 28364 18294 28416
rect 20993 28407 21051 28413
rect 20993 28373 21005 28407
rect 21039 28404 21051 28407
rect 21174 28404 21180 28416
rect 21039 28376 21180 28404
rect 21039 28373 21051 28376
rect 20993 28367 21051 28373
rect 21174 28364 21180 28376
rect 21232 28364 21238 28416
rect 22833 28407 22891 28413
rect 22833 28373 22845 28407
rect 22879 28404 22891 28407
rect 25682 28404 25688 28416
rect 22879 28376 25688 28404
rect 22879 28373 22891 28376
rect 22833 28367 22891 28373
rect 25682 28364 25688 28376
rect 25740 28364 25746 28416
rect 25866 28404 25872 28416
rect 25827 28376 25872 28404
rect 25866 28364 25872 28376
rect 25924 28364 25930 28416
rect 28077 28407 28135 28413
rect 28077 28373 28089 28407
rect 28123 28404 28135 28407
rect 28994 28404 29000 28416
rect 28123 28376 29000 28404
rect 28123 28373 28135 28376
rect 28077 28367 28135 28373
rect 28994 28364 29000 28376
rect 29052 28364 29058 28416
rect 29270 28364 29276 28416
rect 29328 28404 29334 28416
rect 29549 28407 29607 28413
rect 29549 28404 29561 28407
rect 29328 28376 29561 28404
rect 29328 28364 29334 28376
rect 29549 28373 29561 28376
rect 29595 28373 29607 28407
rect 29549 28367 29607 28373
rect 31386 28364 31392 28416
rect 31444 28404 31450 28416
rect 31941 28407 31999 28413
rect 31941 28404 31953 28407
rect 31444 28376 31953 28404
rect 31444 28364 31450 28376
rect 31941 28373 31953 28376
rect 31987 28373 31999 28407
rect 31941 28367 31999 28373
rect 1104 28314 42872 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 42872 28314
rect 1104 28240 42872 28262
rect 2130 28200 2136 28212
rect 2091 28172 2136 28200
rect 2130 28160 2136 28172
rect 2188 28160 2194 28212
rect 17770 28200 17776 28212
rect 16132 28172 17540 28200
rect 17731 28172 17776 28200
rect 13998 28092 14004 28144
rect 14056 28132 14062 28144
rect 14642 28132 14648 28144
rect 14056 28104 14648 28132
rect 14056 28092 14062 28104
rect 14642 28092 14648 28104
rect 14700 28092 14706 28144
rect 16132 28141 16160 28172
rect 16117 28135 16175 28141
rect 16117 28101 16129 28135
rect 16163 28101 16175 28135
rect 16117 28095 16175 28101
rect 17034 28092 17040 28144
rect 17092 28132 17098 28144
rect 17092 28104 17137 28132
rect 17092 28092 17098 28104
rect 2225 28067 2283 28073
rect 2225 28033 2237 28067
rect 2271 28064 2283 28067
rect 2590 28064 2596 28076
rect 2271 28036 2596 28064
rect 2271 28033 2283 28036
rect 2225 28027 2283 28033
rect 2590 28024 2596 28036
rect 2648 28024 2654 28076
rect 12710 28064 12716 28076
rect 12671 28036 12716 28064
rect 12710 28024 12716 28036
rect 12768 28024 12774 28076
rect 14458 28064 14464 28076
rect 14419 28036 14464 28064
rect 14458 28024 14464 28036
rect 14516 28024 14522 28076
rect 14550 28024 14556 28076
rect 14608 28064 14614 28076
rect 15565 28067 15623 28073
rect 15565 28064 15577 28067
rect 14608 28036 15577 28064
rect 14608 28024 14614 28036
rect 15488 27928 15516 28036
rect 15565 28033 15577 28036
rect 15611 28033 15623 28067
rect 15838 28064 15844 28076
rect 15799 28036 15844 28064
rect 15565 28027 15623 28033
rect 15838 28024 15844 28036
rect 15896 28024 15902 28076
rect 15930 28024 15936 28076
rect 15988 28064 15994 28076
rect 16807 28067 16865 28073
rect 16807 28064 16819 28067
rect 15988 28036 16033 28064
rect 16132 28036 16819 28064
rect 15988 28024 15994 28036
rect 15654 27996 15660 28008
rect 15567 27968 15660 27996
rect 15654 27956 15660 27968
rect 15712 27996 15718 28008
rect 16132 27996 16160 28036
rect 16807 28033 16819 28036
rect 16853 28033 16865 28067
rect 16807 28027 16865 28033
rect 16945 28067 17003 28073
rect 16945 28033 16957 28067
rect 16991 28033 17003 28067
rect 16945 28027 17003 28033
rect 15712 27968 16160 27996
rect 15712 27956 15718 27968
rect 16960 27928 16988 28027
rect 17126 28024 17132 28076
rect 17184 28064 17190 28076
rect 17220 28067 17278 28073
rect 17220 28064 17232 28067
rect 17184 28036 17232 28064
rect 17184 28024 17190 28036
rect 17220 28033 17232 28036
rect 17266 28033 17278 28067
rect 17220 28027 17278 28033
rect 17310 28024 17316 28076
rect 17368 28064 17374 28076
rect 17512 28064 17540 28172
rect 17770 28160 17776 28172
rect 17828 28160 17834 28212
rect 20254 28200 20260 28212
rect 20215 28172 20260 28200
rect 20254 28160 20260 28172
rect 20312 28160 20318 28212
rect 26326 28200 26332 28212
rect 26287 28172 26332 28200
rect 26326 28160 26332 28172
rect 26384 28160 26390 28212
rect 27890 28160 27896 28212
rect 27948 28200 27954 28212
rect 28442 28200 28448 28212
rect 27948 28172 28448 28200
rect 27948 28160 27954 28172
rect 28442 28160 28448 28172
rect 28500 28160 28506 28212
rect 28629 28203 28687 28209
rect 28629 28169 28641 28203
rect 28675 28200 28687 28203
rect 29638 28200 29644 28212
rect 28675 28172 29644 28200
rect 28675 28169 28687 28172
rect 28629 28163 28687 28169
rect 29638 28160 29644 28172
rect 29696 28160 29702 28212
rect 29733 28203 29791 28209
rect 29733 28169 29745 28203
rect 29779 28200 29791 28203
rect 30466 28200 30472 28212
rect 29779 28172 30472 28200
rect 29779 28169 29791 28172
rect 29733 28163 29791 28169
rect 30466 28160 30472 28172
rect 30524 28160 30530 28212
rect 41414 28200 41420 28212
rect 41375 28172 41420 28200
rect 41414 28160 41420 28172
rect 41472 28160 41478 28212
rect 19797 28135 19855 28141
rect 19797 28101 19809 28135
rect 19843 28132 19855 28135
rect 20346 28132 20352 28144
rect 19843 28104 20352 28132
rect 19843 28101 19855 28104
rect 19797 28095 19855 28101
rect 20346 28092 20352 28104
rect 20404 28092 20410 28144
rect 21726 28092 21732 28144
rect 21784 28132 21790 28144
rect 22833 28135 22891 28141
rect 22833 28132 22845 28135
rect 21784 28104 22845 28132
rect 21784 28092 21790 28104
rect 22833 28101 22845 28104
rect 22879 28101 22891 28135
rect 22833 28095 22891 28101
rect 25866 28092 25872 28144
rect 25924 28132 25930 28144
rect 26050 28132 26056 28144
rect 25924 28104 26056 28132
rect 25924 28092 25930 28104
rect 26050 28092 26056 28104
rect 26108 28132 26114 28144
rect 26145 28135 26203 28141
rect 26145 28132 26157 28135
rect 26108 28104 26157 28132
rect 26108 28092 26114 28104
rect 26145 28101 26157 28104
rect 26191 28101 26203 28135
rect 30377 28135 30435 28141
rect 26145 28095 26203 28101
rect 28276 28104 29684 28132
rect 18141 28067 18199 28073
rect 18141 28064 18153 28067
rect 17368 28036 17413 28064
rect 17512 28036 18153 28064
rect 17368 28024 17374 28036
rect 18141 28033 18153 28036
rect 18187 28033 18199 28067
rect 18141 28027 18199 28033
rect 18230 28024 18236 28076
rect 18288 28064 18294 28076
rect 18782 28064 18788 28076
rect 18288 28036 18333 28064
rect 18743 28036 18788 28064
rect 18288 28024 18294 28036
rect 18782 28024 18788 28036
rect 18840 28064 18846 28076
rect 19613 28067 19671 28073
rect 19613 28064 19625 28067
rect 18840 28036 19625 28064
rect 18840 28024 18846 28036
rect 19613 28033 19625 28036
rect 19659 28033 19671 28067
rect 20438 28064 20444 28076
rect 20399 28036 20444 28064
rect 19613 28027 19671 28033
rect 20438 28024 20444 28036
rect 20496 28024 20502 28076
rect 24112 28067 24170 28073
rect 24112 28033 24124 28067
rect 24158 28064 24170 28067
rect 24394 28064 24400 28076
rect 24158 28036 24400 28064
rect 24158 28033 24170 28036
rect 24112 28027 24170 28033
rect 24394 28024 24400 28036
rect 24452 28024 24458 28076
rect 25774 28024 25780 28076
rect 25832 28064 25838 28076
rect 28276 28073 28304 28104
rect 25961 28067 26019 28073
rect 25961 28064 25973 28067
rect 25832 28036 25973 28064
rect 25832 28024 25838 28036
rect 25961 28033 25973 28036
rect 26007 28033 26019 28067
rect 25961 28027 26019 28033
rect 28261 28067 28319 28073
rect 28261 28033 28273 28067
rect 28307 28033 28319 28067
rect 28442 28064 28448 28076
rect 28403 28036 28448 28064
rect 28261 28027 28319 28033
rect 28442 28024 28448 28036
rect 28500 28024 28506 28076
rect 29086 28064 29092 28076
rect 29047 28036 29092 28064
rect 29086 28024 29092 28036
rect 29144 28024 29150 28076
rect 29518 28073 29546 28104
rect 29252 28067 29310 28073
rect 29252 28033 29264 28067
rect 29298 28064 29310 28067
rect 29352 28067 29410 28073
rect 29298 28033 29316 28064
rect 29252 28027 29316 28033
rect 29352 28033 29364 28067
rect 29398 28033 29410 28067
rect 29352 28027 29410 28033
rect 29477 28067 29546 28073
rect 29477 28033 29489 28067
rect 29523 28036 29546 28067
rect 29656 28064 29684 28104
rect 30377 28101 30389 28135
rect 30423 28132 30435 28135
rect 31573 28135 31631 28141
rect 31573 28132 31585 28135
rect 30423 28104 31585 28132
rect 30423 28101 30435 28104
rect 30377 28095 30435 28101
rect 31573 28101 31585 28104
rect 31619 28132 31631 28135
rect 32766 28132 32772 28144
rect 31619 28104 31754 28132
rect 32727 28104 32772 28132
rect 31619 28101 31631 28104
rect 31573 28095 31631 28101
rect 31294 28064 31300 28076
rect 29656 28036 31300 28064
rect 29523 28033 29535 28036
rect 29477 28027 29535 28033
rect 17862 27956 17868 28008
rect 17920 27996 17926 28008
rect 17957 27999 18015 28005
rect 17957 27996 17969 27999
rect 17920 27968 17969 27996
rect 17920 27956 17926 27968
rect 17957 27965 17969 27968
rect 18003 27965 18015 27999
rect 17957 27959 18015 27965
rect 18046 27956 18052 28008
rect 18104 27996 18110 28008
rect 23017 27999 23075 28005
rect 18104 27968 18149 27996
rect 18104 27956 18110 27968
rect 23017 27965 23029 27999
rect 23063 27996 23075 27999
rect 23658 27996 23664 28008
rect 23063 27968 23664 27996
rect 23063 27965 23075 27968
rect 23017 27959 23075 27965
rect 23658 27956 23664 27968
rect 23716 27996 23722 28008
rect 23845 27999 23903 28005
rect 23845 27996 23857 27999
rect 23716 27968 23857 27996
rect 23716 27956 23722 27968
rect 23845 27965 23857 27968
rect 23891 27965 23903 27999
rect 23845 27959 23903 27965
rect 28169 27999 28227 28005
rect 28169 27965 28181 27999
rect 28215 27965 28227 27999
rect 28169 27959 28227 27965
rect 28353 27999 28411 28005
rect 28353 27965 28365 27999
rect 28399 27996 28411 27999
rect 28994 27996 29000 28008
rect 28399 27968 29000 27996
rect 28399 27965 28411 27968
rect 28353 27959 28411 27965
rect 15488 27900 16988 27928
rect 28184 27928 28212 27959
rect 28994 27956 29000 27968
rect 29052 27956 29058 28008
rect 29288 27940 29316 28027
rect 29380 27940 29408 28027
rect 31294 28024 31300 28036
rect 31352 28024 31358 28076
rect 31389 28067 31447 28073
rect 31389 28033 31401 28067
rect 31435 28064 31447 28067
rect 31478 28064 31484 28076
rect 31435 28036 31484 28064
rect 31435 28033 31447 28036
rect 31389 28027 31447 28033
rect 31478 28024 31484 28036
rect 31536 28024 31542 28076
rect 28810 27928 28816 27940
rect 28184 27900 28816 27928
rect 28810 27888 28816 27900
rect 28868 27928 28874 27940
rect 29086 27928 29092 27940
rect 28868 27900 29092 27928
rect 28868 27888 28874 27900
rect 29086 27888 29092 27900
rect 29144 27888 29150 27940
rect 29270 27888 29276 27940
rect 29328 27888 29334 27940
rect 29362 27888 29368 27940
rect 29420 27888 29426 27940
rect 31726 27928 31754 28104
rect 32766 28092 32772 28104
rect 32824 28092 32830 28144
rect 33226 28092 33232 28144
rect 33284 28132 33290 28144
rect 33565 28135 33623 28141
rect 33565 28132 33577 28135
rect 33284 28104 33577 28132
rect 33284 28092 33290 28104
rect 33565 28101 33577 28104
rect 33611 28101 33623 28135
rect 33565 28095 33623 28101
rect 33781 28135 33839 28141
rect 33781 28101 33793 28135
rect 33827 28101 33839 28135
rect 33781 28095 33839 28101
rect 32582 28064 32588 28076
rect 32543 28036 32588 28064
rect 32582 28024 32588 28036
rect 32640 28024 32646 28076
rect 32858 28024 32864 28076
rect 32916 28064 32922 28076
rect 33796 28064 33824 28095
rect 32916 28036 33824 28064
rect 34885 28067 34943 28073
rect 32916 28024 32922 28036
rect 34885 28033 34897 28067
rect 34931 28064 34943 28067
rect 41230 28064 41236 28076
rect 34931 28036 41236 28064
rect 34931 28033 34943 28036
rect 34885 28027 34943 28033
rect 41230 28024 41236 28036
rect 41288 28064 41294 28076
rect 41325 28067 41383 28073
rect 41325 28064 41337 28067
rect 41288 28036 41337 28064
rect 41288 28024 41294 28036
rect 41325 28033 41337 28036
rect 41371 28033 41383 28067
rect 41325 28027 41383 28033
rect 32490 27928 32496 27940
rect 31726 27900 32496 27928
rect 32490 27888 32496 27900
rect 32548 27888 32554 27940
rect 32953 27931 33011 27937
rect 32953 27897 32965 27931
rect 32999 27928 33011 27931
rect 32999 27900 33640 27928
rect 32999 27897 33011 27900
rect 32953 27891 33011 27897
rect 12526 27860 12532 27872
rect 12487 27832 12532 27860
rect 12526 27820 12532 27832
rect 12584 27820 12590 27872
rect 14829 27863 14887 27869
rect 14829 27829 14841 27863
rect 14875 27860 14887 27863
rect 15102 27860 15108 27872
rect 14875 27832 15108 27860
rect 14875 27829 14887 27832
rect 14829 27823 14887 27829
rect 15102 27820 15108 27832
rect 15160 27820 15166 27872
rect 16669 27863 16727 27869
rect 16669 27829 16681 27863
rect 16715 27860 16727 27863
rect 16758 27860 16764 27872
rect 16715 27832 16764 27860
rect 16715 27829 16727 27832
rect 16669 27823 16727 27829
rect 16758 27820 16764 27832
rect 16816 27820 16822 27872
rect 18966 27860 18972 27872
rect 18927 27832 18972 27860
rect 18966 27820 18972 27832
rect 19024 27820 19030 27872
rect 25225 27863 25283 27869
rect 25225 27829 25237 27863
rect 25271 27860 25283 27863
rect 26234 27860 26240 27872
rect 25271 27832 26240 27860
rect 25271 27829 25283 27832
rect 25225 27823 25283 27829
rect 26234 27820 26240 27832
rect 26292 27860 26298 27872
rect 27430 27860 27436 27872
rect 26292 27832 27436 27860
rect 26292 27820 26298 27832
rect 27430 27820 27436 27832
rect 27488 27820 27494 27872
rect 28166 27820 28172 27872
rect 28224 27860 28230 27872
rect 28626 27860 28632 27872
rect 28224 27832 28632 27860
rect 28224 27820 28230 27832
rect 28626 27820 28632 27832
rect 28684 27820 28690 27872
rect 30285 27863 30343 27869
rect 30285 27829 30297 27863
rect 30331 27860 30343 27863
rect 30374 27860 30380 27872
rect 30331 27832 30380 27860
rect 30331 27829 30343 27832
rect 30285 27823 30343 27829
rect 30374 27820 30380 27832
rect 30432 27860 30438 27872
rect 31662 27860 31668 27872
rect 30432 27832 31668 27860
rect 30432 27820 30438 27832
rect 31662 27820 31668 27832
rect 31720 27820 31726 27872
rect 33410 27860 33416 27872
rect 33371 27832 33416 27860
rect 33410 27820 33416 27832
rect 33468 27820 33474 27872
rect 33612 27869 33640 27900
rect 33597 27863 33655 27869
rect 33597 27829 33609 27863
rect 33643 27829 33655 27863
rect 33597 27823 33655 27829
rect 34885 27863 34943 27869
rect 34885 27829 34897 27863
rect 34931 27860 34943 27863
rect 35618 27860 35624 27872
rect 34931 27832 35624 27860
rect 34931 27829 34943 27832
rect 34885 27823 34943 27829
rect 35618 27820 35624 27832
rect 35676 27820 35682 27872
rect 1104 27770 42872 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 42872 27770
rect 1104 27696 42872 27718
rect 17862 27656 17868 27668
rect 16776 27628 17868 27656
rect 15381 27591 15439 27597
rect 15381 27557 15393 27591
rect 15427 27588 15439 27591
rect 16776 27588 16804 27628
rect 17862 27616 17868 27628
rect 17920 27616 17926 27668
rect 20349 27659 20407 27665
rect 20349 27625 20361 27659
rect 20395 27625 20407 27659
rect 20349 27619 20407 27625
rect 15427 27560 16804 27588
rect 16853 27591 16911 27597
rect 15427 27557 15439 27560
rect 15381 27551 15439 27557
rect 16853 27557 16865 27591
rect 16899 27588 16911 27591
rect 18046 27588 18052 27600
rect 16899 27560 18052 27588
rect 16899 27557 16911 27560
rect 16853 27551 16911 27557
rect 18046 27548 18052 27560
rect 18104 27548 18110 27600
rect 18598 27588 18604 27600
rect 18511 27560 18604 27588
rect 18598 27548 18604 27560
rect 18656 27588 18662 27600
rect 20162 27588 20168 27600
rect 18656 27560 20168 27588
rect 18656 27548 18662 27560
rect 20162 27548 20168 27560
rect 20220 27548 20226 27600
rect 20364 27588 20392 27619
rect 20438 27616 20444 27668
rect 20496 27656 20502 27668
rect 20533 27659 20591 27665
rect 20533 27656 20545 27659
rect 20496 27628 20545 27656
rect 20496 27616 20502 27628
rect 20533 27625 20545 27628
rect 20579 27625 20591 27659
rect 20533 27619 20591 27625
rect 21174 27616 21180 27668
rect 21232 27656 21238 27668
rect 22557 27659 22615 27665
rect 22557 27656 22569 27659
rect 21232 27628 22569 27656
rect 21232 27616 21238 27628
rect 22557 27625 22569 27628
rect 22603 27625 22615 27659
rect 24394 27656 24400 27668
rect 24355 27628 24400 27656
rect 22557 27619 22615 27625
rect 24394 27616 24400 27628
rect 24452 27616 24458 27668
rect 25958 27656 25964 27668
rect 25919 27628 25964 27656
rect 25958 27616 25964 27628
rect 26016 27616 26022 27668
rect 28166 27656 28172 27668
rect 28127 27628 28172 27656
rect 28166 27616 28172 27628
rect 28224 27616 28230 27668
rect 28810 27656 28816 27668
rect 28771 27628 28816 27656
rect 28810 27616 28816 27628
rect 28868 27616 28874 27668
rect 29086 27616 29092 27668
rect 29144 27656 29150 27668
rect 29549 27659 29607 27665
rect 29549 27656 29561 27659
rect 29144 27628 29561 27656
rect 29144 27616 29150 27628
rect 29549 27625 29561 27628
rect 29595 27625 29607 27659
rect 31573 27659 31631 27665
rect 31573 27656 31585 27659
rect 29549 27619 29607 27625
rect 30116 27628 31585 27656
rect 30116 27600 30144 27628
rect 31573 27625 31585 27628
rect 31619 27656 31631 27659
rect 32582 27656 32588 27668
rect 31619 27628 32588 27656
rect 31619 27625 31631 27628
rect 31573 27619 31631 27625
rect 32582 27616 32588 27628
rect 32640 27616 32646 27668
rect 20993 27591 21051 27597
rect 20993 27588 21005 27591
rect 20364 27560 21005 27588
rect 20993 27557 21005 27560
rect 21039 27557 21051 27591
rect 22370 27588 22376 27600
rect 22331 27560 22376 27588
rect 20993 27551 21051 27557
rect 22370 27548 22376 27560
rect 22428 27588 22434 27600
rect 23753 27591 23811 27597
rect 22428 27560 23428 27588
rect 22428 27548 22434 27560
rect 11882 27520 11888 27532
rect 11843 27492 11888 27520
rect 11882 27480 11888 27492
rect 11940 27480 11946 27532
rect 16390 27520 16396 27532
rect 16351 27492 16396 27520
rect 16390 27480 16396 27492
rect 16448 27480 16454 27532
rect 17126 27520 17132 27532
rect 16592 27492 17132 27520
rect 12152 27455 12210 27461
rect 12152 27421 12164 27455
rect 12198 27452 12210 27455
rect 12526 27452 12532 27464
rect 12198 27424 12532 27452
rect 12198 27421 12210 27424
rect 12152 27415 12210 27421
rect 12526 27412 12532 27424
rect 12584 27412 12590 27464
rect 14458 27452 14464 27464
rect 14419 27424 14464 27452
rect 14458 27412 14464 27424
rect 14516 27412 14522 27464
rect 14642 27452 14648 27464
rect 14603 27424 14648 27452
rect 14642 27412 14648 27424
rect 14700 27412 14706 27464
rect 15102 27452 15108 27464
rect 15063 27424 15108 27452
rect 15102 27412 15108 27424
rect 15160 27412 15166 27464
rect 16301 27455 16359 27461
rect 16301 27421 16313 27455
rect 16347 27452 16359 27455
rect 16482 27452 16488 27464
rect 16347 27424 16488 27452
rect 16347 27421 16359 27424
rect 16301 27415 16359 27421
rect 16482 27412 16488 27424
rect 16540 27412 16546 27464
rect 16592 27461 16620 27492
rect 17126 27480 17132 27492
rect 17184 27480 17190 27532
rect 17402 27480 17408 27532
rect 17460 27520 17466 27532
rect 23290 27520 23296 27532
rect 17460 27492 23296 27520
rect 17460 27480 17466 27492
rect 23290 27480 23296 27492
rect 23348 27480 23354 27532
rect 23400 27529 23428 27560
rect 23753 27557 23765 27591
rect 23799 27588 23811 27591
rect 24486 27588 24492 27600
rect 23799 27560 24492 27588
rect 23799 27557 23811 27560
rect 23753 27551 23811 27557
rect 24486 27548 24492 27560
rect 24544 27588 24550 27600
rect 25130 27588 25136 27600
rect 24544 27560 25136 27588
rect 24544 27548 24550 27560
rect 25130 27548 25136 27560
rect 25188 27548 25194 27600
rect 29733 27591 29791 27597
rect 29733 27557 29745 27591
rect 29779 27588 29791 27591
rect 30098 27588 30104 27600
rect 29779 27560 30104 27588
rect 29779 27557 29791 27560
rect 29733 27551 29791 27557
rect 30098 27548 30104 27560
rect 30156 27548 30162 27600
rect 30837 27591 30895 27597
rect 30837 27588 30849 27591
rect 30208 27560 30849 27588
rect 30208 27532 30236 27560
rect 30837 27557 30849 27560
rect 30883 27557 30895 27591
rect 30837 27551 30895 27557
rect 23385 27523 23443 27529
rect 23385 27489 23397 27523
rect 23431 27489 23443 27523
rect 28902 27520 28908 27532
rect 23385 27483 23443 27489
rect 28000 27492 28908 27520
rect 16577 27455 16635 27461
rect 16577 27421 16589 27455
rect 16623 27421 16635 27455
rect 16577 27415 16635 27421
rect 16669 27455 16727 27461
rect 16669 27421 16681 27455
rect 16715 27452 16727 27455
rect 17034 27452 17040 27464
rect 16715 27424 17040 27452
rect 16715 27421 16727 27424
rect 16669 27415 16727 27421
rect 17034 27412 17040 27424
rect 17092 27452 17098 27464
rect 17586 27452 17592 27464
rect 17092 27424 17592 27452
rect 17092 27412 17098 27424
rect 17586 27412 17592 27424
rect 17644 27412 17650 27464
rect 19981 27455 20039 27461
rect 19981 27421 19993 27455
rect 20027 27452 20039 27455
rect 20806 27452 20812 27464
rect 20027 27424 20812 27452
rect 20027 27421 20039 27424
rect 19981 27415 20039 27421
rect 20806 27412 20812 27424
rect 20864 27412 20870 27464
rect 21174 27452 21180 27464
rect 21135 27424 21180 27452
rect 21174 27412 21180 27424
rect 21232 27412 21238 27464
rect 21450 27452 21456 27464
rect 21411 27424 21456 27452
rect 21450 27412 21456 27424
rect 21508 27412 21514 27464
rect 22925 27455 22983 27461
rect 22925 27421 22937 27455
rect 22971 27452 22983 27455
rect 23198 27452 23204 27464
rect 22971 27424 23204 27452
rect 22971 27421 22983 27424
rect 22925 27415 22983 27421
rect 23198 27412 23204 27424
rect 23256 27412 23262 27464
rect 24578 27452 24584 27464
rect 24539 27424 24584 27452
rect 24578 27412 24584 27424
rect 24636 27412 24642 27464
rect 25038 27412 25044 27464
rect 25096 27452 25102 27464
rect 25774 27452 25780 27464
rect 25096 27424 25780 27452
rect 25096 27412 25102 27424
rect 25774 27412 25780 27424
rect 25832 27452 25838 27464
rect 25869 27455 25927 27461
rect 25869 27452 25881 27455
rect 25832 27424 25881 27452
rect 25832 27412 25838 27424
rect 25869 27421 25881 27424
rect 25915 27421 25927 27455
rect 26050 27452 26056 27464
rect 26011 27424 26056 27452
rect 25869 27415 25927 27421
rect 26050 27412 26056 27424
rect 26108 27452 26114 27464
rect 26605 27455 26663 27461
rect 26605 27452 26617 27455
rect 26108 27424 26617 27452
rect 26108 27412 26114 27424
rect 26605 27421 26617 27424
rect 26651 27421 26663 27455
rect 26605 27415 26663 27421
rect 27798 27412 27804 27464
rect 27856 27452 27862 27464
rect 28000 27461 28028 27492
rect 28902 27480 28908 27492
rect 28960 27480 28966 27532
rect 28994 27480 29000 27532
rect 29052 27520 29058 27532
rect 30190 27520 30196 27532
rect 29052 27492 30196 27520
rect 29052 27480 29058 27492
rect 30190 27480 30196 27492
rect 30248 27480 30254 27532
rect 31662 27480 31668 27532
rect 31720 27520 31726 27532
rect 32769 27523 32827 27529
rect 32769 27520 32781 27523
rect 31720 27492 32781 27520
rect 31720 27480 31726 27492
rect 32769 27489 32781 27492
rect 32815 27489 32827 27523
rect 32769 27483 32827 27489
rect 27985 27455 28043 27461
rect 27985 27452 27997 27455
rect 27856 27424 27997 27452
rect 27856 27412 27862 27424
rect 27985 27421 27997 27424
rect 28031 27421 28043 27455
rect 27985 27415 28043 27421
rect 28169 27455 28227 27461
rect 28169 27421 28181 27455
rect 28215 27452 28227 27455
rect 28534 27452 28540 27464
rect 28215 27424 28540 27452
rect 28215 27421 28227 27424
rect 28169 27415 28227 27421
rect 28534 27412 28540 27424
rect 28592 27412 28598 27464
rect 28626 27412 28632 27464
rect 28684 27452 28690 27464
rect 29086 27452 29092 27464
rect 28684 27424 29092 27452
rect 28684 27412 28690 27424
rect 29086 27412 29092 27424
rect 29144 27452 29150 27464
rect 29362 27452 29368 27464
rect 29144 27424 29368 27452
rect 29144 27412 29150 27424
rect 29362 27412 29368 27424
rect 29420 27412 29426 27464
rect 32125 27455 32183 27461
rect 32125 27421 32137 27455
rect 32171 27452 32183 27455
rect 33410 27452 33416 27464
rect 32171 27424 33416 27452
rect 32171 27421 32183 27424
rect 32125 27415 32183 27421
rect 33410 27412 33416 27424
rect 33468 27412 33474 27464
rect 41417 27455 41475 27461
rect 41417 27421 41429 27455
rect 41463 27452 41475 27455
rect 41506 27452 41512 27464
rect 41463 27424 41512 27452
rect 41463 27421 41475 27424
rect 41417 27415 41475 27421
rect 41506 27412 41512 27424
rect 41564 27412 41570 27464
rect 15381 27387 15439 27393
rect 15381 27353 15393 27387
rect 15427 27384 15439 27387
rect 16758 27384 16764 27396
rect 15427 27356 16764 27384
rect 15427 27353 15439 27356
rect 15381 27347 15439 27353
rect 16758 27344 16764 27356
rect 16816 27344 16822 27396
rect 18138 27344 18144 27396
rect 18196 27384 18202 27396
rect 18325 27387 18383 27393
rect 18325 27384 18337 27387
rect 18196 27356 18337 27384
rect 18196 27344 18202 27356
rect 18325 27353 18337 27356
rect 18371 27384 18383 27387
rect 18782 27384 18788 27396
rect 18371 27356 18788 27384
rect 18371 27353 18383 27356
rect 18325 27347 18383 27353
rect 18782 27344 18788 27356
rect 18840 27344 18846 27396
rect 20349 27387 20407 27393
rect 20349 27353 20361 27387
rect 20395 27384 20407 27387
rect 20990 27384 20996 27396
rect 20395 27356 20996 27384
rect 20395 27353 20407 27356
rect 20349 27347 20407 27353
rect 20990 27344 20996 27356
rect 21048 27384 21054 27396
rect 21048 27356 22968 27384
rect 21048 27344 21054 27356
rect 13262 27316 13268 27328
rect 13223 27288 13268 27316
rect 13262 27276 13268 27288
rect 13320 27276 13326 27328
rect 14645 27319 14703 27325
rect 14645 27285 14657 27319
rect 14691 27316 14703 27319
rect 15197 27319 15255 27325
rect 15197 27316 15209 27319
rect 14691 27288 15209 27316
rect 14691 27285 14703 27288
rect 14645 27279 14703 27285
rect 15197 27285 15209 27288
rect 15243 27285 15255 27319
rect 15197 27279 15255 27285
rect 21361 27319 21419 27325
rect 21361 27285 21373 27319
rect 21407 27316 21419 27319
rect 21726 27316 21732 27328
rect 21407 27288 21732 27316
rect 21407 27285 21419 27288
rect 21361 27279 21419 27285
rect 21726 27276 21732 27288
rect 21784 27276 21790 27328
rect 22554 27316 22560 27328
rect 22515 27288 22560 27316
rect 22554 27276 22560 27288
rect 22612 27276 22618 27328
rect 22940 27316 22968 27356
rect 27890 27344 27896 27396
rect 27948 27384 27954 27396
rect 28781 27387 28839 27393
rect 28781 27384 28793 27387
rect 27948 27356 28793 27384
rect 27948 27344 27954 27356
rect 28781 27353 28793 27356
rect 28827 27353 28839 27387
rect 28994 27384 29000 27396
rect 28955 27356 29000 27384
rect 28781 27347 28839 27353
rect 28994 27344 29000 27356
rect 29052 27344 29058 27396
rect 30009 27387 30067 27393
rect 30009 27353 30021 27387
rect 30055 27353 30067 27387
rect 30009 27347 30067 27353
rect 23845 27319 23903 27325
rect 23845 27316 23857 27319
rect 22940 27288 23857 27316
rect 23845 27285 23857 27288
rect 23891 27285 23903 27319
rect 26694 27316 26700 27328
rect 26655 27288 26700 27316
rect 23845 27279 23903 27285
rect 26694 27276 26700 27288
rect 26752 27276 26758 27328
rect 28626 27276 28632 27328
rect 28684 27316 28690 27328
rect 28684 27288 28729 27316
rect 28684 27276 28690 27288
rect 28902 27276 28908 27328
rect 28960 27316 28966 27328
rect 29822 27316 29828 27328
rect 28960 27288 29828 27316
rect 28960 27276 28966 27288
rect 29822 27276 29828 27288
rect 29880 27316 29886 27328
rect 30024 27316 30052 27347
rect 30742 27344 30748 27396
rect 30800 27384 30806 27396
rect 30837 27387 30895 27393
rect 30837 27384 30849 27387
rect 30800 27356 30849 27384
rect 30800 27344 30806 27356
rect 30837 27353 30849 27356
rect 30883 27353 30895 27387
rect 33014 27387 33072 27393
rect 33014 27384 33026 27387
rect 30837 27347 30895 27353
rect 32324 27356 33026 27384
rect 29880 27288 30052 27316
rect 29880 27276 29886 27288
rect 30282 27276 30288 27328
rect 30340 27316 30346 27328
rect 31297 27319 31355 27325
rect 31297 27316 31309 27319
rect 30340 27288 31309 27316
rect 30340 27276 30346 27288
rect 31297 27285 31309 27288
rect 31343 27285 31355 27319
rect 31297 27279 31355 27285
rect 31386 27276 31392 27328
rect 31444 27316 31450 27328
rect 32324 27325 32352 27356
rect 33014 27353 33026 27356
rect 33060 27353 33072 27387
rect 33014 27347 33072 27353
rect 32309 27319 32367 27325
rect 31444 27288 31489 27316
rect 31444 27276 31450 27288
rect 32309 27285 32321 27319
rect 32355 27285 32367 27319
rect 32309 27279 32367 27285
rect 32766 27276 32772 27328
rect 32824 27316 32830 27328
rect 34146 27316 34152 27328
rect 32824 27288 34152 27316
rect 32824 27276 32830 27288
rect 34146 27276 34152 27288
rect 34204 27276 34210 27328
rect 41509 27319 41567 27325
rect 41509 27285 41521 27319
rect 41555 27316 41567 27319
rect 41690 27316 41696 27328
rect 41555 27288 41696 27316
rect 41555 27285 41567 27288
rect 41509 27279 41567 27285
rect 41690 27276 41696 27288
rect 41748 27276 41754 27328
rect 1104 27226 42872 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 42872 27226
rect 1104 27152 42872 27174
rect 12710 27072 12716 27124
rect 12768 27112 12774 27124
rect 12989 27115 13047 27121
rect 12989 27112 13001 27115
rect 12768 27084 13001 27112
rect 12768 27072 12774 27084
rect 12989 27081 13001 27084
rect 13035 27081 13047 27115
rect 12989 27075 13047 27081
rect 19426 27072 19432 27124
rect 19484 27112 19490 27124
rect 20625 27115 20683 27121
rect 20625 27112 20637 27115
rect 19484 27084 20637 27112
rect 19484 27072 19490 27084
rect 20625 27081 20637 27084
rect 20671 27081 20683 27115
rect 23198 27112 23204 27124
rect 23159 27084 23204 27112
rect 20625 27075 20683 27081
rect 23198 27072 23204 27084
rect 23256 27072 23262 27124
rect 23290 27072 23296 27124
rect 23348 27112 23354 27124
rect 24029 27115 24087 27121
rect 23348 27084 23704 27112
rect 23348 27072 23354 27084
rect 20806 27044 20812 27056
rect 15488 27016 20024 27044
rect 13173 26979 13231 26985
rect 13173 26945 13185 26979
rect 13219 26976 13231 26979
rect 14734 26976 14740 26988
rect 13219 26948 14740 26976
rect 13219 26945 13231 26948
rect 13173 26939 13231 26945
rect 14734 26936 14740 26948
rect 14792 26936 14798 26988
rect 15286 26976 15292 26988
rect 15199 26948 15292 26976
rect 15286 26936 15292 26948
rect 15344 26976 15350 26988
rect 15488 26976 15516 27016
rect 15344 26948 15516 26976
rect 15565 26979 15623 26985
rect 15344 26936 15350 26948
rect 15565 26945 15577 26979
rect 15611 26976 15623 26979
rect 15654 26976 15660 26988
rect 15611 26948 15660 26976
rect 15611 26945 15623 26948
rect 15565 26939 15623 26945
rect 13262 26868 13268 26920
rect 13320 26908 13326 26920
rect 13357 26911 13415 26917
rect 13357 26908 13369 26911
rect 13320 26880 13369 26908
rect 13320 26868 13326 26880
rect 13357 26877 13369 26880
rect 13403 26877 13415 26911
rect 13357 26871 13415 26877
rect 13372 26772 13400 26871
rect 14458 26868 14464 26920
rect 14516 26908 14522 26920
rect 15473 26911 15531 26917
rect 15473 26908 15485 26911
rect 14516 26880 15485 26908
rect 14516 26868 14522 26880
rect 15473 26877 15485 26880
rect 15519 26877 15531 26911
rect 15473 26871 15531 26877
rect 15378 26840 15384 26852
rect 15339 26812 15384 26840
rect 15378 26800 15384 26812
rect 15436 26800 15442 26852
rect 15580 26772 15608 26939
rect 15654 26936 15660 26948
rect 15712 26936 15718 26988
rect 16666 26976 16672 26988
rect 16627 26948 16672 26976
rect 16666 26936 16672 26948
rect 16724 26936 16730 26988
rect 19518 26936 19524 26988
rect 19576 26976 19582 26988
rect 19806 26979 19864 26985
rect 19806 26976 19818 26979
rect 19576 26948 19818 26976
rect 19576 26936 19582 26948
rect 19806 26945 19818 26948
rect 19852 26945 19864 26979
rect 19806 26939 19864 26945
rect 16942 26908 16948 26920
rect 16903 26880 16948 26908
rect 16942 26868 16948 26880
rect 17000 26868 17006 26920
rect 19996 26908 20024 27016
rect 20548 27016 20812 27044
rect 20548 26985 20576 27016
rect 20806 27004 20812 27016
rect 20864 27004 20870 27056
rect 23566 27044 23572 27056
rect 21836 27016 23572 27044
rect 21836 26985 21864 27016
rect 23566 27004 23572 27016
rect 23624 27004 23630 27056
rect 23676 27053 23704 27084
rect 24029 27081 24041 27115
rect 24075 27112 24087 27115
rect 27798 27112 27804 27124
rect 24075 27084 27804 27112
rect 24075 27081 24087 27084
rect 24029 27075 24087 27081
rect 27798 27072 27804 27084
rect 27856 27072 27862 27124
rect 27890 27072 27896 27124
rect 27948 27112 27954 27124
rect 28077 27115 28135 27121
rect 28077 27112 28089 27115
rect 27948 27084 28089 27112
rect 27948 27072 27954 27084
rect 28077 27081 28089 27084
rect 28123 27081 28135 27115
rect 41966 27112 41972 27124
rect 28077 27075 28135 27081
rect 31726 27084 41972 27112
rect 23661 27047 23719 27053
rect 23661 27013 23673 27047
rect 23707 27013 23719 27047
rect 23661 27007 23719 27013
rect 20073 26979 20131 26985
rect 20073 26945 20085 26979
rect 20119 26976 20131 26979
rect 20533 26979 20591 26985
rect 20119 26948 20484 26976
rect 20119 26945 20131 26948
rect 20073 26939 20131 26945
rect 20456 26908 20484 26948
rect 20533 26945 20545 26979
rect 20579 26945 20591 26979
rect 21821 26979 21879 26985
rect 21821 26976 21833 26979
rect 20533 26939 20591 26945
rect 20916 26948 21833 26976
rect 20916 26908 20944 26948
rect 21821 26945 21833 26948
rect 21867 26945 21879 26979
rect 21821 26939 21879 26945
rect 21910 26936 21916 26988
rect 21968 26976 21974 26988
rect 22077 26979 22135 26985
rect 22077 26976 22089 26979
rect 21968 26948 22089 26976
rect 21968 26936 21974 26948
rect 22077 26945 22089 26948
rect 22123 26945 22135 26979
rect 23676 26976 23704 27007
rect 23842 27004 23848 27056
rect 23900 27053 23906 27056
rect 23900 27047 23919 27053
rect 23907 27013 23919 27047
rect 31726 27044 31754 27084
rect 41966 27072 41972 27084
rect 42024 27072 42030 27124
rect 33226 27044 33232 27056
rect 23900 27007 23919 27013
rect 23952 27016 31754 27044
rect 33060 27016 33232 27044
rect 23900 27004 23906 27007
rect 23952 26976 23980 27016
rect 23676 26948 23980 26976
rect 22077 26939 22135 26945
rect 25590 26936 25596 26988
rect 25648 26976 25654 26988
rect 26053 26979 26111 26985
rect 26053 26976 26065 26979
rect 25648 26948 26065 26976
rect 25648 26936 25654 26948
rect 26053 26945 26065 26948
rect 26099 26945 26111 26979
rect 26053 26939 26111 26945
rect 28261 26979 28319 26985
rect 28261 26945 28273 26979
rect 28307 26976 28319 26979
rect 28350 26976 28356 26988
rect 28307 26948 28356 26976
rect 28307 26945 28319 26948
rect 28261 26939 28319 26945
rect 28350 26936 28356 26948
rect 28408 26936 28414 26988
rect 28810 26936 28816 26988
rect 28868 26976 28874 26988
rect 28905 26979 28963 26985
rect 28905 26976 28917 26979
rect 28868 26948 28917 26976
rect 28868 26936 28874 26948
rect 28905 26945 28917 26948
rect 28951 26945 28963 26979
rect 29178 26976 29184 26988
rect 29139 26948 29184 26976
rect 28905 26939 28963 26945
rect 29178 26936 29184 26948
rect 29236 26936 29242 26988
rect 30742 26936 30748 26988
rect 30800 26976 30806 26988
rect 30929 26979 30987 26985
rect 30929 26976 30941 26979
rect 30800 26948 30941 26976
rect 30800 26936 30806 26948
rect 30929 26945 30941 26948
rect 30975 26945 30987 26979
rect 31386 26976 31392 26988
rect 31347 26948 31392 26976
rect 30929 26939 30987 26945
rect 31386 26936 31392 26948
rect 31444 26936 31450 26988
rect 32769 26979 32827 26985
rect 32769 26945 32781 26979
rect 32815 26976 32827 26979
rect 32858 26976 32864 26988
rect 32815 26948 32864 26976
rect 32815 26945 32827 26948
rect 32769 26939 32827 26945
rect 32858 26936 32864 26948
rect 32916 26936 32922 26988
rect 33060 26985 33088 27016
rect 33226 27004 33232 27016
rect 33284 27004 33290 27056
rect 34698 27044 34704 27056
rect 33888 27016 34704 27044
rect 32953 26979 33011 26985
rect 32953 26945 32965 26979
rect 32999 26945 33011 26979
rect 32953 26939 33011 26945
rect 33045 26979 33103 26985
rect 33045 26945 33057 26979
rect 33091 26945 33103 26979
rect 33045 26939 33103 26945
rect 33137 26979 33195 26985
rect 33137 26945 33149 26979
rect 33183 26976 33195 26979
rect 33778 26976 33784 26988
rect 33183 26948 33784 26976
rect 33183 26945 33195 26948
rect 33137 26939 33195 26945
rect 19996 26880 20116 26908
rect 20456 26880 20944 26908
rect 20088 26840 20116 26880
rect 20990 26868 20996 26920
rect 21048 26908 21054 26920
rect 28442 26908 28448 26920
rect 21048 26880 21093 26908
rect 28355 26880 28448 26908
rect 21048 26868 21054 26880
rect 28442 26868 28448 26880
rect 28500 26908 28506 26920
rect 28500 26880 30052 26908
rect 28500 26868 28506 26880
rect 20088 26812 20944 26840
rect 13372 26744 15608 26772
rect 15749 26775 15807 26781
rect 15749 26741 15761 26775
rect 15795 26772 15807 26775
rect 16761 26775 16819 26781
rect 16761 26772 16773 26775
rect 15795 26744 16773 26772
rect 15795 26741 15807 26744
rect 15749 26735 15807 26741
rect 16761 26741 16773 26744
rect 16807 26741 16819 26775
rect 16761 26735 16819 26741
rect 16850 26732 16856 26784
rect 16908 26772 16914 26784
rect 18693 26775 18751 26781
rect 16908 26744 16953 26772
rect 16908 26732 16914 26744
rect 18693 26741 18705 26775
rect 18739 26772 18751 26775
rect 19426 26772 19432 26784
rect 18739 26744 19432 26772
rect 18739 26741 18751 26744
rect 18693 26735 18751 26741
rect 19426 26732 19432 26744
rect 19484 26732 19490 26784
rect 19702 26732 19708 26784
rect 19760 26772 19766 26784
rect 20809 26775 20867 26781
rect 20809 26772 20821 26775
rect 19760 26744 20821 26772
rect 19760 26732 19766 26744
rect 20809 26741 20821 26744
rect 20855 26741 20867 26775
rect 20916 26772 20944 26812
rect 22940 26812 23888 26840
rect 22940 26772 22968 26812
rect 23860 26781 23888 26812
rect 30024 26784 30052 26880
rect 30834 26868 30840 26920
rect 30892 26908 30898 26920
rect 31205 26911 31263 26917
rect 31205 26908 31217 26911
rect 30892 26880 31217 26908
rect 30892 26868 30898 26880
rect 31205 26877 31217 26880
rect 31251 26877 31263 26911
rect 32968 26908 32996 26939
rect 33778 26936 33784 26948
rect 33836 26936 33842 26988
rect 33888 26985 33916 27016
rect 34698 27004 34704 27016
rect 34756 27004 34762 27056
rect 41690 27044 41696 27056
rect 41651 27016 41696 27044
rect 41690 27004 41696 27016
rect 41748 27004 41754 27056
rect 33873 26979 33931 26985
rect 33873 26945 33885 26979
rect 33919 26945 33931 26979
rect 34129 26979 34187 26985
rect 34129 26976 34141 26979
rect 33873 26939 33931 26945
rect 33980 26948 34141 26976
rect 33318 26908 33324 26920
rect 32968 26880 33324 26908
rect 31205 26871 31263 26877
rect 33318 26868 33324 26880
rect 33376 26868 33382 26920
rect 33413 26911 33471 26917
rect 33413 26877 33425 26911
rect 33459 26908 33471 26911
rect 33980 26908 34008 26948
rect 34129 26945 34141 26948
rect 34175 26945 34187 26979
rect 34129 26939 34187 26945
rect 41322 26908 41328 26920
rect 33459 26880 34008 26908
rect 41283 26880 41328 26908
rect 33459 26877 33471 26880
rect 33413 26871 33471 26877
rect 41322 26868 41328 26880
rect 41380 26868 41386 26920
rect 41874 26908 41880 26920
rect 41835 26880 41880 26908
rect 41874 26868 41880 26880
rect 41932 26868 41938 26920
rect 20916 26744 22968 26772
rect 23845 26775 23903 26781
rect 20809 26735 20867 26741
rect 23845 26741 23857 26775
rect 23891 26741 23903 26775
rect 23845 26735 23903 26741
rect 26237 26775 26295 26781
rect 26237 26741 26249 26775
rect 26283 26772 26295 26775
rect 26326 26772 26332 26784
rect 26283 26744 26332 26772
rect 26283 26741 26295 26744
rect 26237 26735 26295 26741
rect 26326 26732 26332 26744
rect 26384 26732 26390 26784
rect 30006 26732 30012 26784
rect 30064 26772 30070 26784
rect 30282 26772 30288 26784
rect 30064 26744 30288 26772
rect 30064 26732 30070 26744
rect 30282 26732 30288 26744
rect 30340 26772 30346 26784
rect 31021 26775 31079 26781
rect 31021 26772 31033 26775
rect 30340 26744 31033 26772
rect 30340 26732 30346 26744
rect 31021 26741 31033 26744
rect 31067 26741 31079 26775
rect 31021 26735 31079 26741
rect 31573 26775 31631 26781
rect 31573 26741 31585 26775
rect 31619 26772 31631 26775
rect 32030 26772 32036 26784
rect 31619 26744 32036 26772
rect 31619 26741 31631 26744
rect 31573 26735 31631 26741
rect 32030 26732 32036 26744
rect 32088 26732 32094 26784
rect 35253 26775 35311 26781
rect 35253 26741 35265 26775
rect 35299 26772 35311 26775
rect 35342 26772 35348 26784
rect 35299 26744 35348 26772
rect 35299 26741 35311 26744
rect 35253 26735 35311 26741
rect 35342 26732 35348 26744
rect 35400 26732 35406 26784
rect 1104 26682 42872 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 42872 26682
rect 1104 26608 42872 26630
rect 15470 26528 15476 26580
rect 15528 26568 15534 26580
rect 16393 26571 16451 26577
rect 16393 26568 16405 26571
rect 15528 26540 16405 26568
rect 15528 26528 15534 26540
rect 16393 26537 16405 26540
rect 16439 26537 16451 26571
rect 19518 26568 19524 26580
rect 19479 26540 19524 26568
rect 16393 26531 16451 26537
rect 19518 26528 19524 26540
rect 19576 26528 19582 26580
rect 19889 26571 19947 26577
rect 19889 26537 19901 26571
rect 19935 26568 19947 26571
rect 20806 26568 20812 26580
rect 19935 26540 20812 26568
rect 19935 26537 19947 26540
rect 19889 26531 19947 26537
rect 20806 26528 20812 26540
rect 20864 26528 20870 26580
rect 21821 26571 21879 26577
rect 21821 26537 21833 26571
rect 21867 26568 21879 26571
rect 21910 26568 21916 26580
rect 21867 26540 21916 26568
rect 21867 26537 21879 26540
rect 21821 26531 21879 26537
rect 21910 26528 21916 26540
rect 21968 26528 21974 26580
rect 25409 26571 25467 26577
rect 25409 26537 25421 26571
rect 25455 26537 25467 26571
rect 25590 26568 25596 26580
rect 25551 26540 25596 26568
rect 25409 26531 25467 26537
rect 13541 26503 13599 26509
rect 13541 26469 13553 26503
rect 13587 26500 13599 26503
rect 14458 26500 14464 26512
rect 13587 26472 14464 26500
rect 13587 26469 13599 26472
rect 13541 26463 13599 26469
rect 12066 26392 12072 26444
rect 12124 26432 12130 26444
rect 14384 26441 14412 26472
rect 14458 26460 14464 26472
rect 14516 26500 14522 26512
rect 14516 26472 14872 26500
rect 14516 26460 14522 26472
rect 12161 26435 12219 26441
rect 12161 26432 12173 26435
rect 12124 26404 12173 26432
rect 12124 26392 12130 26404
rect 12161 26401 12173 26404
rect 12207 26401 12219 26435
rect 12161 26395 12219 26401
rect 14369 26435 14427 26441
rect 14369 26401 14381 26435
rect 14415 26401 14427 26435
rect 14734 26432 14740 26444
rect 14695 26404 14740 26432
rect 14369 26395 14427 26401
rect 12176 26364 12204 26395
rect 14734 26392 14740 26404
rect 14792 26392 14798 26444
rect 14844 26432 14872 26472
rect 15378 26460 15384 26512
rect 15436 26500 15442 26512
rect 15565 26503 15623 26509
rect 15565 26500 15577 26503
rect 15436 26472 15577 26500
rect 15436 26460 15442 26472
rect 15565 26469 15577 26472
rect 15611 26469 15623 26503
rect 22554 26500 22560 26512
rect 15565 26463 15623 26469
rect 16224 26472 17264 26500
rect 15657 26435 15715 26441
rect 15657 26432 15669 26435
rect 14844 26404 15669 26432
rect 15657 26401 15669 26404
rect 15703 26401 15715 26435
rect 15657 26395 15715 26401
rect 12894 26364 12900 26376
rect 12176 26336 12900 26364
rect 12894 26324 12900 26336
rect 12952 26324 12958 26376
rect 14277 26367 14335 26373
rect 14277 26333 14289 26367
rect 14323 26333 14335 26367
rect 14277 26327 14335 26333
rect 15381 26367 15439 26373
rect 15381 26333 15393 26367
rect 15427 26364 15439 26367
rect 15562 26364 15568 26376
rect 15427 26336 15568 26364
rect 15427 26333 15439 26336
rect 15381 26327 15439 26333
rect 12428 26299 12486 26305
rect 12428 26265 12440 26299
rect 12474 26296 12486 26299
rect 14093 26299 14151 26305
rect 14093 26296 14105 26299
rect 12474 26268 14105 26296
rect 12474 26265 12486 26268
rect 12428 26259 12486 26265
rect 14093 26265 14105 26268
rect 14139 26265 14151 26299
rect 14292 26296 14320 26327
rect 15562 26324 15568 26336
rect 15620 26364 15626 26376
rect 16224 26364 16252 26472
rect 16301 26435 16359 26441
rect 16301 26401 16313 26435
rect 16347 26432 16359 26435
rect 16390 26432 16396 26444
rect 16347 26404 16396 26432
rect 16347 26401 16359 26404
rect 16301 26395 16359 26401
rect 16390 26392 16396 26404
rect 16448 26392 16454 26444
rect 15620 26336 16252 26364
rect 16485 26367 16543 26373
rect 15620 26324 15626 26336
rect 16485 26333 16497 26367
rect 16531 26333 16543 26367
rect 16485 26327 16543 26333
rect 16577 26367 16635 26373
rect 16577 26333 16589 26367
rect 16623 26364 16635 26367
rect 16758 26364 16764 26376
rect 16623 26336 16764 26364
rect 16623 26333 16635 26336
rect 16577 26327 16635 26333
rect 15286 26296 15292 26308
rect 14292 26268 15292 26296
rect 14093 26259 14151 26265
rect 15286 26256 15292 26268
rect 15344 26256 15350 26308
rect 16500 26296 16528 26327
rect 16758 26324 16764 26336
rect 16816 26324 16822 26376
rect 17236 26373 17264 26472
rect 19996 26472 22560 26500
rect 19426 26392 19432 26444
rect 19484 26432 19490 26444
rect 19996 26441 20024 26472
rect 22554 26460 22560 26472
rect 22612 26500 22618 26512
rect 23014 26500 23020 26512
rect 22612 26472 23020 26500
rect 22612 26460 22618 26472
rect 23014 26460 23020 26472
rect 23072 26460 23078 26512
rect 25424 26500 25452 26531
rect 25590 26528 25596 26540
rect 25648 26528 25654 26580
rect 26084 26540 28028 26568
rect 26084 26500 26112 26540
rect 25424 26472 26112 26500
rect 19981 26435 20039 26441
rect 19981 26432 19993 26435
rect 19484 26404 19993 26432
rect 19484 26392 19490 26404
rect 19981 26401 19993 26404
rect 20027 26401 20039 26435
rect 19981 26395 20039 26401
rect 20625 26435 20683 26441
rect 20625 26401 20637 26435
rect 20671 26432 20683 26435
rect 20671 26404 21404 26432
rect 20671 26401 20683 26404
rect 20625 26395 20683 26401
rect 17221 26367 17279 26373
rect 17221 26333 17233 26367
rect 17267 26364 17279 26367
rect 17402 26364 17408 26376
rect 17267 26336 17408 26364
rect 17267 26333 17279 26336
rect 17221 26327 17279 26333
rect 17402 26324 17408 26336
rect 17460 26324 17466 26376
rect 19702 26364 19708 26376
rect 19663 26336 19708 26364
rect 19702 26324 19708 26336
rect 19760 26324 19766 26376
rect 20533 26367 20591 26373
rect 20533 26333 20545 26367
rect 20579 26333 20591 26367
rect 20533 26327 20591 26333
rect 20717 26367 20775 26373
rect 20717 26333 20729 26367
rect 20763 26333 20775 26367
rect 20717 26327 20775 26333
rect 16666 26296 16672 26308
rect 16500 26268 16672 26296
rect 16666 26256 16672 26268
rect 16724 26296 16730 26308
rect 16942 26296 16948 26308
rect 16724 26268 16948 26296
rect 16724 26256 16730 26268
rect 16942 26256 16948 26268
rect 17000 26296 17006 26308
rect 17129 26299 17187 26305
rect 17129 26296 17141 26299
rect 17000 26268 17141 26296
rect 17000 26256 17006 26268
rect 17129 26265 17141 26268
rect 17175 26265 17187 26299
rect 17129 26259 17187 26265
rect 15194 26228 15200 26240
rect 15155 26200 15200 26228
rect 15194 26188 15200 26200
rect 15252 26188 15258 26240
rect 20548 26228 20576 26327
rect 20732 26296 20760 26327
rect 20990 26324 20996 26376
rect 21048 26364 21054 26376
rect 21376 26373 21404 26404
rect 23198 26392 23204 26444
rect 23256 26432 23262 26444
rect 23385 26435 23443 26441
rect 23385 26432 23397 26435
rect 23256 26404 23397 26432
rect 23256 26392 23262 26404
rect 23385 26401 23397 26404
rect 23431 26401 23443 26435
rect 23385 26395 23443 26401
rect 23658 26392 23664 26444
rect 23716 26432 23722 26444
rect 26053 26435 26111 26441
rect 26053 26432 26065 26435
rect 23716 26404 26065 26432
rect 23716 26392 23722 26404
rect 26053 26401 26065 26404
rect 26099 26401 26111 26435
rect 26053 26395 26111 26401
rect 21177 26367 21235 26373
rect 21177 26364 21189 26367
rect 21048 26336 21189 26364
rect 21048 26324 21054 26336
rect 21177 26333 21189 26336
rect 21223 26333 21235 26367
rect 21177 26327 21235 26333
rect 21361 26367 21419 26373
rect 21361 26333 21373 26367
rect 21407 26333 21419 26367
rect 21361 26327 21419 26333
rect 21450 26324 21456 26376
rect 21508 26364 21514 26376
rect 21591 26367 21649 26373
rect 21508 26336 21553 26364
rect 21508 26324 21514 26336
rect 21591 26333 21603 26367
rect 21637 26364 21649 26367
rect 21726 26364 21732 26376
rect 21637 26336 21732 26364
rect 21637 26333 21671 26336
rect 21591 26327 21671 26333
rect 21643 26296 21671 26327
rect 21726 26324 21732 26336
rect 21784 26364 21790 26376
rect 23109 26367 23167 26373
rect 23109 26364 23121 26367
rect 21784 26336 23121 26364
rect 21784 26324 21790 26336
rect 23109 26333 23121 26336
rect 23155 26364 23167 26367
rect 23842 26364 23848 26376
rect 23155 26336 23848 26364
rect 23155 26333 23167 26336
rect 23109 26327 23167 26333
rect 23842 26324 23848 26336
rect 23900 26324 23906 26376
rect 24578 26364 24584 26376
rect 24539 26336 24584 26364
rect 24578 26324 24584 26336
rect 24636 26324 24642 26376
rect 25038 26364 25044 26376
rect 24999 26336 25044 26364
rect 25038 26324 25044 26336
rect 25096 26324 25102 26376
rect 26326 26373 26332 26376
rect 26320 26364 26332 26373
rect 26287 26336 26332 26364
rect 26320 26327 26332 26336
rect 26326 26324 26332 26327
rect 26384 26324 26390 26376
rect 28000 26364 28028 26540
rect 28810 26528 28816 26580
rect 28868 26568 28874 26580
rect 29549 26571 29607 26577
rect 29549 26568 29561 26571
rect 28868 26540 29561 26568
rect 28868 26528 28874 26540
rect 29549 26537 29561 26540
rect 29595 26537 29607 26571
rect 29549 26531 29607 26537
rect 30009 26571 30067 26577
rect 30009 26537 30021 26571
rect 30055 26568 30067 26571
rect 30282 26568 30288 26580
rect 30055 26540 30288 26568
rect 30055 26537 30067 26540
rect 30009 26531 30067 26537
rect 30282 26528 30288 26540
rect 30340 26528 30346 26580
rect 31846 26528 31852 26580
rect 31904 26568 31910 26580
rect 32033 26571 32091 26577
rect 32033 26568 32045 26571
rect 31904 26540 32045 26568
rect 31904 26528 31910 26540
rect 32033 26537 32045 26540
rect 32079 26568 32091 26571
rect 32766 26568 32772 26580
rect 32079 26540 32772 26568
rect 32079 26537 32091 26540
rect 32033 26531 32091 26537
rect 32766 26528 32772 26540
rect 32824 26528 32830 26580
rect 33226 26528 33232 26580
rect 33284 26568 33290 26580
rect 34054 26568 34060 26580
rect 33284 26540 34060 26568
rect 33284 26528 33290 26540
rect 34054 26528 34060 26540
rect 34112 26528 34118 26580
rect 41785 26571 41843 26577
rect 41785 26537 41797 26571
rect 41831 26568 41843 26571
rect 41874 26568 41880 26580
rect 41831 26540 41880 26568
rect 41831 26537 41843 26540
rect 41785 26531 41843 26537
rect 41874 26528 41880 26540
rect 41932 26528 41938 26580
rect 28997 26503 29055 26509
rect 28997 26469 29009 26503
rect 29043 26500 29055 26503
rect 29362 26500 29368 26512
rect 29043 26472 29368 26500
rect 29043 26469 29055 26472
rect 28997 26463 29055 26469
rect 29362 26460 29368 26472
rect 29420 26460 29426 26512
rect 32306 26500 32312 26512
rect 30116 26472 32312 26500
rect 28353 26435 28411 26441
rect 28353 26401 28365 26435
rect 28399 26432 28411 26435
rect 29086 26432 29092 26444
rect 28399 26404 29092 26432
rect 28399 26401 28411 26404
rect 28353 26395 28411 26401
rect 29086 26392 29092 26404
rect 29144 26392 29150 26444
rect 29822 26432 29828 26444
rect 29783 26404 29828 26432
rect 29822 26392 29828 26404
rect 29880 26392 29886 26444
rect 28442 26364 28448 26376
rect 28000 26336 28448 26364
rect 28442 26324 28448 26336
rect 28500 26364 28506 26376
rect 28629 26367 28687 26373
rect 28629 26364 28641 26367
rect 28500 26336 28641 26364
rect 28500 26324 28506 26336
rect 28629 26333 28641 26336
rect 28675 26333 28687 26367
rect 28629 26327 28687 26333
rect 28838 26367 28896 26373
rect 28838 26333 28850 26367
rect 28884 26364 28896 26367
rect 28994 26364 29000 26376
rect 28884 26336 29000 26364
rect 28884 26333 28896 26336
rect 28838 26327 28896 26333
rect 28994 26324 29000 26336
rect 29052 26324 29058 26376
rect 30116 26373 30144 26472
rect 32306 26460 32312 26472
rect 32364 26500 32370 26512
rect 32401 26503 32459 26509
rect 32401 26500 32413 26503
rect 32364 26472 32413 26500
rect 32364 26460 32370 26472
rect 32401 26469 32413 26472
rect 32447 26469 32459 26503
rect 32401 26463 32459 26469
rect 33505 26503 33563 26509
rect 33505 26469 33517 26503
rect 33551 26500 33563 26503
rect 34698 26500 34704 26512
rect 33551 26472 34704 26500
rect 33551 26469 33563 26472
rect 33505 26463 33563 26469
rect 34698 26460 34704 26472
rect 34756 26460 34762 26512
rect 30190 26392 30196 26444
rect 30248 26432 30254 26444
rect 31021 26435 31079 26441
rect 31021 26432 31033 26435
rect 30248 26404 31033 26432
rect 30248 26392 30254 26404
rect 31021 26401 31033 26404
rect 31067 26401 31079 26435
rect 31021 26395 31079 26401
rect 32582 26392 32588 26444
rect 32640 26432 32646 26444
rect 32640 26404 34008 26432
rect 32640 26392 32646 26404
rect 30101 26367 30159 26373
rect 30101 26333 30113 26367
rect 30147 26333 30159 26367
rect 30742 26364 30748 26376
rect 30703 26336 30748 26364
rect 30101 26327 30159 26333
rect 20732 26268 21671 26296
rect 28534 26256 28540 26308
rect 28592 26296 28598 26308
rect 30116 26296 30144 26327
rect 30742 26324 30748 26336
rect 30800 26324 30806 26376
rect 32030 26364 32036 26376
rect 31991 26336 32036 26364
rect 32030 26324 32036 26336
rect 32088 26324 32094 26376
rect 32217 26367 32275 26373
rect 32217 26333 32229 26367
rect 32263 26333 32275 26367
rect 32217 26327 32275 26333
rect 28592 26268 30144 26296
rect 32232 26296 32260 26327
rect 32490 26324 32496 26376
rect 32548 26364 32554 26376
rect 33980 26373 34008 26404
rect 33304 26367 33362 26373
rect 33304 26364 33316 26367
rect 32548 26336 33316 26364
rect 32548 26324 32554 26336
rect 33304 26333 33316 26336
rect 33350 26333 33362 26367
rect 33304 26327 33362 26333
rect 33965 26367 34023 26373
rect 33965 26333 33977 26367
rect 34011 26333 34023 26367
rect 34146 26364 34152 26376
rect 34107 26336 34152 26364
rect 33965 26327 34023 26333
rect 34146 26324 34152 26336
rect 34204 26324 34210 26376
rect 34885 26367 34943 26373
rect 34885 26333 34897 26367
rect 34931 26364 34943 26367
rect 35342 26364 35348 26376
rect 34931 26336 35348 26364
rect 34931 26333 34943 26336
rect 34885 26327 34943 26333
rect 35342 26324 35348 26336
rect 35400 26324 35406 26376
rect 33870 26296 33876 26308
rect 32232 26268 33876 26296
rect 28592 26256 28598 26268
rect 33870 26256 33876 26268
rect 33928 26296 33934 26308
rect 34793 26299 34851 26305
rect 34793 26296 34805 26299
rect 33928 26268 34805 26296
rect 33928 26256 33934 26268
rect 34793 26265 34805 26268
rect 34839 26265 34851 26299
rect 34793 26259 34851 26265
rect 21542 26228 21548 26240
rect 20548 26200 21548 26228
rect 21542 26188 21548 26200
rect 21600 26188 21606 26240
rect 24394 26228 24400 26240
rect 24355 26200 24400 26228
rect 24394 26188 24400 26200
rect 24452 26188 24458 26240
rect 25406 26228 25412 26240
rect 25367 26200 25412 26228
rect 25406 26188 25412 26200
rect 25464 26188 25470 26240
rect 27433 26231 27491 26237
rect 27433 26197 27445 26231
rect 27479 26228 27491 26231
rect 27522 26228 27528 26240
rect 27479 26200 27528 26228
rect 27479 26197 27491 26200
rect 27433 26191 27491 26197
rect 27522 26188 27528 26200
rect 27580 26188 27586 26240
rect 28718 26188 28724 26240
rect 28776 26228 28782 26240
rect 28776 26200 28821 26228
rect 28776 26188 28782 26200
rect 1104 26138 42872 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 42872 26138
rect 1104 26064 42872 26086
rect 14369 26027 14427 26033
rect 14369 25993 14381 26027
rect 14415 26024 14427 26027
rect 14734 26024 14740 26036
rect 14415 25996 14740 26024
rect 14415 25993 14427 25996
rect 14369 25987 14427 25993
rect 14734 25984 14740 25996
rect 14792 25984 14798 26036
rect 15473 26027 15531 26033
rect 15473 25993 15485 26027
rect 15519 26024 15531 26027
rect 15562 26024 15568 26036
rect 15519 25996 15568 26024
rect 15519 25993 15531 25996
rect 15473 25987 15531 25993
rect 15562 25984 15568 25996
rect 15620 25984 15626 26036
rect 20806 26024 20812 26036
rect 20767 25996 20812 26024
rect 20806 25984 20812 25996
rect 20864 25984 20870 26036
rect 20972 26027 21030 26033
rect 20972 25993 20984 26027
rect 21018 26024 21030 26027
rect 21542 26024 21548 26036
rect 21018 25996 21548 26024
rect 21018 25993 21030 25996
rect 20972 25987 21030 25993
rect 21542 25984 21548 25996
rect 21600 25984 21606 26036
rect 24946 26024 24952 26036
rect 22066 25996 24952 26024
rect 17862 25956 17868 25968
rect 14568 25928 17868 25956
rect 14568 25897 14596 25928
rect 17862 25916 17868 25928
rect 17920 25956 17926 25968
rect 21174 25956 21180 25968
rect 17920 25928 21036 25956
rect 21087 25928 21180 25956
rect 17920 25916 17926 25928
rect 14553 25891 14611 25897
rect 14553 25857 14565 25891
rect 14599 25857 14611 25891
rect 14553 25851 14611 25857
rect 14737 25891 14795 25897
rect 14737 25857 14749 25891
rect 14783 25888 14795 25891
rect 15194 25888 15200 25900
rect 14783 25860 15200 25888
rect 14783 25857 14795 25860
rect 14737 25851 14795 25857
rect 15194 25848 15200 25860
rect 15252 25848 15258 25900
rect 15381 25891 15439 25897
rect 15381 25857 15393 25891
rect 15427 25857 15439 25891
rect 15381 25851 15439 25857
rect 15657 25891 15715 25897
rect 15657 25857 15669 25891
rect 15703 25888 15715 25891
rect 16850 25888 16856 25900
rect 15703 25860 16856 25888
rect 15703 25857 15715 25860
rect 15657 25851 15715 25857
rect 14829 25823 14887 25829
rect 14829 25789 14841 25823
rect 14875 25820 14887 25823
rect 15396 25820 15424 25851
rect 16850 25848 16856 25860
rect 16908 25848 16914 25900
rect 17954 25848 17960 25900
rect 18012 25888 18018 25900
rect 18426 25891 18484 25897
rect 18426 25888 18438 25891
rect 18012 25860 18438 25888
rect 18012 25848 18018 25860
rect 18426 25857 18438 25860
rect 18472 25857 18484 25891
rect 18690 25888 18696 25900
rect 18651 25860 18696 25888
rect 18426 25851 18484 25857
rect 18690 25848 18696 25860
rect 18748 25848 18754 25900
rect 21008 25888 21036 25928
rect 21174 25916 21180 25928
rect 21232 25956 21238 25968
rect 21450 25956 21456 25968
rect 21232 25928 21456 25956
rect 21232 25916 21238 25928
rect 21450 25916 21456 25928
rect 21508 25916 21514 25968
rect 22066 25888 22094 25996
rect 24946 25984 24952 25996
rect 25004 25984 25010 26036
rect 25406 25984 25412 26036
rect 25464 26024 25470 26036
rect 25501 26027 25559 26033
rect 25501 26024 25513 26027
rect 25464 25996 25513 26024
rect 25464 25984 25470 25996
rect 25501 25993 25513 25996
rect 25547 25993 25559 26027
rect 25501 25987 25559 25993
rect 28629 26027 28687 26033
rect 28629 25993 28641 26027
rect 28675 26024 28687 26027
rect 28810 26024 28816 26036
rect 28675 25996 28816 26024
rect 28675 25993 28687 25996
rect 28629 25987 28687 25993
rect 28810 25984 28816 25996
rect 28868 25984 28874 26036
rect 28994 26024 29000 26036
rect 28955 25996 29000 26024
rect 28994 25984 29000 25996
rect 29052 25984 29058 26036
rect 30742 25984 30748 26036
rect 30800 26024 30806 26036
rect 31021 26027 31079 26033
rect 31021 26024 31033 26027
rect 30800 25996 31033 26024
rect 30800 25984 30806 25996
rect 31021 25993 31033 25996
rect 31067 25993 31079 26027
rect 31021 25987 31079 25993
rect 32493 26027 32551 26033
rect 32493 25993 32505 26027
rect 32539 26024 32551 26027
rect 32858 26024 32864 26036
rect 32539 25996 32864 26024
rect 32539 25993 32551 25996
rect 32493 25987 32551 25993
rect 32858 25984 32864 25996
rect 32916 25984 32922 26036
rect 33318 25984 33324 26036
rect 33376 26024 33382 26036
rect 33873 26027 33931 26033
rect 33873 26024 33885 26027
rect 33376 25996 33885 26024
rect 33376 25984 33382 25996
rect 33873 25993 33885 25996
rect 33919 25993 33931 26027
rect 33873 25987 33931 25993
rect 23928 25959 23986 25965
rect 23928 25925 23940 25959
rect 23974 25956 23986 25959
rect 24394 25956 24400 25968
rect 23974 25928 24400 25956
rect 23974 25925 23986 25928
rect 23928 25919 23986 25925
rect 24394 25916 24400 25928
rect 24452 25916 24458 25968
rect 25869 25959 25927 25965
rect 25869 25925 25881 25959
rect 25915 25956 25927 25959
rect 27522 25956 27528 25968
rect 25915 25928 27528 25956
rect 25915 25925 25927 25928
rect 25869 25919 25927 25925
rect 27522 25916 27528 25928
rect 27580 25916 27586 25968
rect 23014 25888 23020 25900
rect 21008 25860 22094 25888
rect 22975 25860 23020 25888
rect 23014 25848 23020 25860
rect 23072 25848 23078 25900
rect 23658 25888 23664 25900
rect 23619 25860 23664 25888
rect 23658 25848 23664 25860
rect 23716 25848 23722 25900
rect 24302 25848 24308 25900
rect 24360 25888 24366 25900
rect 24360 25860 25452 25888
rect 24360 25848 24366 25860
rect 15562 25820 15568 25832
rect 14875 25792 15240 25820
rect 15396 25792 15568 25820
rect 14875 25789 14887 25792
rect 14829 25783 14887 25789
rect 15212 25764 15240 25792
rect 15562 25780 15568 25792
rect 15620 25780 15626 25832
rect 25424 25820 25452 25860
rect 25498 25848 25504 25900
rect 25556 25888 25562 25900
rect 25685 25891 25743 25897
rect 25685 25888 25697 25891
rect 25556 25860 25697 25888
rect 25556 25848 25562 25860
rect 25685 25857 25697 25860
rect 25731 25857 25743 25891
rect 25685 25851 25743 25857
rect 25961 25891 26019 25897
rect 25961 25857 25973 25891
rect 26007 25857 26019 25891
rect 25961 25851 26019 25857
rect 25976 25820 26004 25851
rect 26326 25848 26332 25900
rect 26384 25888 26390 25900
rect 27341 25891 27399 25897
rect 27341 25888 27353 25891
rect 26384 25860 27353 25888
rect 26384 25848 26390 25860
rect 27341 25857 27353 25860
rect 27387 25857 27399 25891
rect 27341 25851 27399 25857
rect 27890 25848 27896 25900
rect 27948 25888 27954 25900
rect 28537 25891 28595 25897
rect 28537 25888 28549 25891
rect 27948 25860 28549 25888
rect 27948 25848 27954 25860
rect 28537 25857 28549 25860
rect 28583 25857 28595 25891
rect 28537 25851 28595 25857
rect 28813 25891 28871 25897
rect 28813 25857 28825 25891
rect 28859 25888 28871 25891
rect 28902 25888 28908 25900
rect 28859 25860 28908 25888
rect 28859 25857 28871 25860
rect 28813 25851 28871 25857
rect 28902 25848 28908 25860
rect 28960 25888 28966 25900
rect 29178 25888 29184 25900
rect 28960 25860 29184 25888
rect 28960 25848 28966 25860
rect 29178 25848 29184 25860
rect 29236 25848 29242 25900
rect 29546 25848 29552 25900
rect 29604 25888 29610 25900
rect 29897 25891 29955 25897
rect 29897 25888 29909 25891
rect 29604 25860 29909 25888
rect 29604 25848 29610 25860
rect 29897 25857 29909 25860
rect 29943 25857 29955 25891
rect 32306 25888 32312 25900
rect 32267 25860 32312 25888
rect 29897 25851 29955 25857
rect 32306 25848 32312 25860
rect 32364 25848 32370 25900
rect 33870 25888 33876 25900
rect 33831 25860 33876 25888
rect 33870 25848 33876 25860
rect 33928 25848 33934 25900
rect 34054 25888 34060 25900
rect 34015 25860 34060 25888
rect 34054 25848 34060 25860
rect 34112 25848 34118 25900
rect 25424 25792 26004 25820
rect 27249 25823 27307 25829
rect 27249 25789 27261 25823
rect 27295 25789 27307 25823
rect 27249 25783 27307 25789
rect 29641 25823 29699 25829
rect 29641 25789 29653 25823
rect 29687 25789 29699 25823
rect 29641 25783 29699 25789
rect 15194 25712 15200 25764
rect 15252 25752 15258 25764
rect 15838 25752 15844 25764
rect 15252 25724 15844 25752
rect 15252 25712 15258 25724
rect 15838 25712 15844 25724
rect 15896 25712 15902 25764
rect 25041 25755 25099 25761
rect 25041 25721 25053 25755
rect 25087 25752 25099 25755
rect 26234 25752 26240 25764
rect 25087 25724 26240 25752
rect 25087 25721 25099 25724
rect 25041 25715 25099 25721
rect 26234 25712 26240 25724
rect 26292 25752 26298 25764
rect 27264 25752 27292 25783
rect 26292 25724 27292 25752
rect 26292 25712 26298 25724
rect 17313 25687 17371 25693
rect 17313 25653 17325 25687
rect 17359 25684 17371 25687
rect 17586 25684 17592 25696
rect 17359 25656 17592 25684
rect 17359 25653 17371 25656
rect 17313 25647 17371 25653
rect 17586 25644 17592 25656
rect 17644 25644 17650 25696
rect 20993 25687 21051 25693
rect 20993 25653 21005 25687
rect 21039 25684 21051 25687
rect 21726 25684 21732 25696
rect 21039 25656 21732 25684
rect 21039 25653 21051 25656
rect 20993 25647 21051 25653
rect 21726 25644 21732 25656
rect 21784 25644 21790 25696
rect 23109 25687 23167 25693
rect 23109 25653 23121 25687
rect 23155 25684 23167 25687
rect 23290 25684 23296 25696
rect 23155 25656 23296 25684
rect 23155 25653 23167 25656
rect 23109 25647 23167 25653
rect 23290 25644 23296 25656
rect 23348 25644 23354 25696
rect 25130 25644 25136 25696
rect 25188 25684 25194 25696
rect 26973 25687 27031 25693
rect 26973 25684 26985 25687
rect 25188 25656 26985 25684
rect 25188 25644 25194 25656
rect 26973 25653 26985 25656
rect 27019 25653 27031 25687
rect 27154 25684 27160 25696
rect 27115 25656 27160 25684
rect 26973 25647 27031 25653
rect 27154 25644 27160 25656
rect 27212 25644 27218 25696
rect 29656 25684 29684 25783
rect 31570 25780 31576 25832
rect 31628 25820 31634 25832
rect 32125 25823 32183 25829
rect 32125 25820 32137 25823
rect 31628 25792 32137 25820
rect 31628 25780 31634 25792
rect 32125 25789 32137 25792
rect 32171 25789 32183 25823
rect 32125 25783 32183 25789
rect 30374 25684 30380 25696
rect 29656 25656 30380 25684
rect 30374 25644 30380 25656
rect 30432 25684 30438 25696
rect 30834 25684 30840 25696
rect 30432 25656 30840 25684
rect 30432 25644 30438 25656
rect 30834 25644 30840 25656
rect 30892 25644 30898 25696
rect 41785 25687 41843 25693
rect 41785 25653 41797 25687
rect 41831 25684 41843 25687
rect 41874 25684 41880 25696
rect 41831 25656 41880 25684
rect 41831 25653 41843 25656
rect 41785 25647 41843 25653
rect 41874 25644 41880 25656
rect 41932 25644 41938 25696
rect 1104 25594 42872 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 42872 25594
rect 1104 25520 42872 25542
rect 15197 25483 15255 25489
rect 15197 25449 15209 25483
rect 15243 25480 15255 25483
rect 15286 25480 15292 25492
rect 15243 25452 15292 25480
rect 15243 25449 15255 25452
rect 15197 25443 15255 25449
rect 15286 25440 15292 25452
rect 15344 25440 15350 25492
rect 15381 25483 15439 25489
rect 15381 25449 15393 25483
rect 15427 25449 15439 25483
rect 15381 25443 15439 25449
rect 24397 25483 24455 25489
rect 24397 25449 24409 25483
rect 24443 25480 24455 25483
rect 24578 25480 24584 25492
rect 24443 25452 24584 25480
rect 24443 25449 24455 25452
rect 24397 25443 24455 25449
rect 15396 25412 15424 25443
rect 24578 25440 24584 25452
rect 24636 25440 24642 25492
rect 25498 25480 25504 25492
rect 25459 25452 25504 25480
rect 25498 25440 25504 25452
rect 25556 25440 25562 25492
rect 28718 25440 28724 25492
rect 28776 25480 28782 25492
rect 28905 25483 28963 25489
rect 28905 25480 28917 25483
rect 28776 25452 28917 25480
rect 28776 25440 28782 25452
rect 28905 25449 28917 25452
rect 28951 25449 28963 25483
rect 30098 25480 30104 25492
rect 30059 25452 30104 25480
rect 28905 25443 28963 25449
rect 30098 25440 30104 25452
rect 30156 25440 30162 25492
rect 30466 25440 30472 25492
rect 30524 25480 30530 25492
rect 33226 25480 33232 25492
rect 30524 25452 33232 25480
rect 30524 25440 30530 25452
rect 33226 25440 33232 25452
rect 33284 25440 33290 25492
rect 25130 25412 25136 25424
rect 15304 25384 15424 25412
rect 24688 25384 25136 25412
rect 15304 25356 15332 25384
rect 15286 25304 15292 25356
rect 15344 25344 15350 25356
rect 16209 25347 16267 25353
rect 15344 25316 16160 25344
rect 15344 25304 15350 25316
rect 14550 25276 14556 25288
rect 14511 25248 14556 25276
rect 14550 25236 14556 25248
rect 14608 25276 14614 25288
rect 15378 25276 15384 25288
rect 14608 25248 15384 25276
rect 14608 25236 14614 25248
rect 15378 25236 15384 25248
rect 15436 25236 15442 25288
rect 15562 25236 15568 25288
rect 15620 25276 15626 25288
rect 16132 25276 16160 25316
rect 16209 25313 16221 25347
rect 16255 25344 16267 25347
rect 16850 25344 16856 25356
rect 16255 25316 16856 25344
rect 16255 25313 16267 25316
rect 16209 25307 16267 25313
rect 16850 25304 16856 25316
rect 16908 25304 16914 25356
rect 17586 25344 17592 25356
rect 17547 25316 17592 25344
rect 17586 25304 17592 25316
rect 17644 25304 17650 25356
rect 24302 25304 24308 25356
rect 24360 25344 24366 25356
rect 24688 25353 24716 25384
rect 25130 25372 25136 25384
rect 25188 25372 25194 25424
rect 24556 25347 24614 25353
rect 24556 25344 24568 25347
rect 24360 25316 24568 25344
rect 24360 25304 24366 25316
rect 24556 25313 24568 25316
rect 24602 25313 24614 25347
rect 24556 25307 24614 25313
rect 24673 25347 24731 25353
rect 24673 25313 24685 25347
rect 24719 25313 24731 25347
rect 24673 25307 24731 25313
rect 25041 25347 25099 25353
rect 25041 25313 25053 25347
rect 25087 25344 25099 25347
rect 25516 25344 25544 25440
rect 31110 25412 31116 25424
rect 27172 25384 31116 25412
rect 27172 25356 27200 25384
rect 31110 25372 31116 25384
rect 31168 25412 31174 25424
rect 31168 25384 32444 25412
rect 31168 25372 31174 25384
rect 25087 25316 25544 25344
rect 25869 25347 25927 25353
rect 25087 25313 25099 25316
rect 25041 25307 25099 25313
rect 25869 25313 25881 25347
rect 25915 25344 25927 25347
rect 26234 25344 26240 25356
rect 25915 25316 26240 25344
rect 25915 25313 25927 25316
rect 25869 25307 25927 25313
rect 26234 25304 26240 25316
rect 26292 25304 26298 25356
rect 26602 25344 26608 25356
rect 26563 25316 26608 25344
rect 26602 25304 26608 25316
rect 26660 25304 26666 25356
rect 26881 25347 26939 25353
rect 26881 25313 26893 25347
rect 26927 25344 26939 25347
rect 27154 25344 27160 25356
rect 26927 25316 27160 25344
rect 26927 25313 26939 25316
rect 26881 25307 26939 25313
rect 27154 25304 27160 25316
rect 27212 25304 27218 25356
rect 30650 25344 30656 25356
rect 30392 25316 30656 25344
rect 16485 25279 16543 25285
rect 16485 25276 16497 25279
rect 15620 25248 15665 25276
rect 16132 25248 16497 25276
rect 15620 25236 15626 25248
rect 16485 25245 16497 25248
rect 16531 25276 16543 25279
rect 16758 25276 16764 25288
rect 16531 25248 16764 25276
rect 16531 25245 16543 25248
rect 16485 25239 16543 25245
rect 16758 25236 16764 25248
rect 16816 25236 16822 25288
rect 17034 25236 17040 25288
rect 17092 25276 17098 25288
rect 17865 25279 17923 25285
rect 17865 25276 17877 25279
rect 17092 25248 17877 25276
rect 17092 25236 17098 25248
rect 17865 25245 17877 25248
rect 17911 25245 17923 25279
rect 17865 25239 17923 25245
rect 20165 25279 20223 25285
rect 20165 25245 20177 25279
rect 20211 25245 20223 25279
rect 20165 25239 20223 25245
rect 20349 25279 20407 25285
rect 20349 25245 20361 25279
rect 20395 25276 20407 25279
rect 20806 25276 20812 25288
rect 20395 25248 20812 25276
rect 20395 25245 20407 25248
rect 20349 25239 20407 25245
rect 14645 25211 14703 25217
rect 14645 25177 14657 25211
rect 14691 25208 14703 25211
rect 16390 25208 16396 25220
rect 14691 25180 16396 25208
rect 14691 25177 14703 25180
rect 14645 25171 14703 25177
rect 16390 25168 16396 25180
rect 16448 25168 16454 25220
rect 20180 25208 20208 25239
rect 20806 25236 20812 25248
rect 20864 25236 20870 25288
rect 25682 25276 25688 25288
rect 25643 25248 25688 25276
rect 25682 25236 25688 25248
rect 25740 25236 25746 25288
rect 28534 25276 28540 25288
rect 28495 25248 28540 25276
rect 28534 25236 28540 25248
rect 28592 25236 28598 25288
rect 30392 25285 30420 25316
rect 30650 25304 30656 25316
rect 30708 25344 30714 25356
rect 31389 25347 31447 25353
rect 31389 25344 31401 25347
rect 30708 25316 31401 25344
rect 30708 25304 30714 25316
rect 31389 25313 31401 25316
rect 31435 25313 31447 25347
rect 31389 25307 31447 25313
rect 32416 25344 32444 25384
rect 32416 25316 33548 25344
rect 32416 25288 32444 25316
rect 30377 25279 30435 25285
rect 30377 25245 30389 25279
rect 30423 25245 30435 25279
rect 30377 25239 30435 25245
rect 30466 25236 30472 25288
rect 30524 25276 30530 25288
rect 30561 25279 30619 25285
rect 30561 25276 30573 25279
rect 30524 25248 30573 25276
rect 30524 25236 30530 25248
rect 30561 25245 30573 25248
rect 30607 25245 30619 25279
rect 31294 25276 31300 25288
rect 31207 25248 31300 25276
rect 30561 25239 30619 25245
rect 31294 25236 31300 25248
rect 31352 25276 31358 25288
rect 31570 25276 31576 25288
rect 31352 25248 31432 25276
rect 31531 25248 31576 25276
rect 31352 25236 31358 25248
rect 21266 25208 21272 25220
rect 20180 25180 21272 25208
rect 21266 25168 21272 25180
rect 21324 25168 21330 25220
rect 27798 25168 27804 25220
rect 27856 25208 27862 25220
rect 28721 25211 28779 25217
rect 28721 25208 28733 25211
rect 27856 25180 28733 25208
rect 27856 25168 27862 25180
rect 28721 25177 28733 25180
rect 28767 25177 28779 25211
rect 31404 25208 31432 25248
rect 31570 25236 31576 25248
rect 31628 25236 31634 25288
rect 32398 25276 32404 25288
rect 32311 25248 32404 25276
rect 32398 25236 32404 25248
rect 32456 25236 32462 25288
rect 32677 25279 32735 25285
rect 32677 25245 32689 25279
rect 32723 25276 32735 25279
rect 33042 25276 33048 25288
rect 32723 25248 33048 25276
rect 32723 25245 32735 25248
rect 32677 25239 32735 25245
rect 33042 25236 33048 25248
rect 33100 25236 33106 25288
rect 33321 25279 33379 25285
rect 33321 25245 33333 25279
rect 33367 25276 33379 25279
rect 33410 25276 33416 25288
rect 33367 25248 33416 25276
rect 33367 25245 33379 25248
rect 33321 25239 33379 25245
rect 32493 25211 32551 25217
rect 32493 25208 32505 25211
rect 31404 25180 32505 25208
rect 28721 25171 28779 25177
rect 32493 25177 32505 25180
rect 32539 25208 32551 25211
rect 32766 25208 32772 25220
rect 32539 25180 32772 25208
rect 32539 25177 32551 25180
rect 32493 25171 32551 25177
rect 32766 25168 32772 25180
rect 32824 25208 32830 25220
rect 33336 25208 33364 25239
rect 33410 25236 33416 25248
rect 33468 25236 33474 25288
rect 33520 25285 33548 25316
rect 33505 25279 33563 25285
rect 33505 25245 33517 25279
rect 33551 25245 33563 25279
rect 33505 25239 33563 25245
rect 40034 25236 40040 25288
rect 40092 25276 40098 25288
rect 40497 25279 40555 25285
rect 40497 25276 40509 25279
rect 40092 25248 40509 25276
rect 40092 25236 40098 25248
rect 40497 25245 40509 25248
rect 40543 25245 40555 25279
rect 40497 25239 40555 25245
rect 41325 25279 41383 25285
rect 41325 25245 41337 25279
rect 41371 25276 41383 25279
rect 41506 25276 41512 25288
rect 41371 25248 41512 25276
rect 41371 25245 41383 25248
rect 41325 25239 41383 25245
rect 41506 25236 41512 25248
rect 41564 25236 41570 25288
rect 41782 25276 41788 25288
rect 41743 25248 41788 25276
rect 41782 25236 41788 25248
rect 41840 25236 41846 25288
rect 32824 25180 33364 25208
rect 32824 25168 32830 25180
rect 40218 25168 40224 25220
rect 40276 25208 40282 25220
rect 41877 25211 41935 25217
rect 41877 25208 41889 25211
rect 40276 25180 41889 25208
rect 40276 25168 40282 25180
rect 41877 25177 41889 25180
rect 41923 25177 41935 25211
rect 41877 25171 41935 25177
rect 20162 25100 20168 25152
rect 20220 25140 20226 25152
rect 20257 25143 20315 25149
rect 20257 25140 20269 25143
rect 20220 25112 20269 25140
rect 20220 25100 20226 25112
rect 20257 25109 20269 25112
rect 20303 25109 20315 25143
rect 20257 25103 20315 25109
rect 23474 25100 23480 25152
rect 23532 25140 23538 25152
rect 24765 25143 24823 25149
rect 24765 25140 24777 25143
rect 23532 25112 24777 25140
rect 23532 25100 23538 25112
rect 24765 25109 24777 25112
rect 24811 25109 24823 25143
rect 30282 25140 30288 25152
rect 30243 25112 30288 25140
rect 24765 25103 24823 25109
rect 30282 25100 30288 25112
rect 30340 25100 30346 25152
rect 30742 25100 30748 25152
rect 30800 25140 30806 25152
rect 31570 25140 31576 25152
rect 30800 25112 31576 25140
rect 30800 25100 30806 25112
rect 31570 25100 31576 25112
rect 31628 25100 31634 25152
rect 31754 25100 31760 25152
rect 31812 25140 31818 25152
rect 31812 25112 31857 25140
rect 31812 25100 31818 25112
rect 32674 25100 32680 25152
rect 32732 25140 32738 25152
rect 32861 25143 32919 25149
rect 32861 25140 32873 25143
rect 32732 25112 32873 25140
rect 32732 25100 32738 25112
rect 32861 25109 32873 25112
rect 32907 25109 32919 25143
rect 33318 25140 33324 25152
rect 33279 25112 33324 25140
rect 32861 25103 32919 25109
rect 33318 25100 33324 25112
rect 33376 25100 33382 25152
rect 40494 25100 40500 25152
rect 40552 25140 40558 25152
rect 41233 25143 41291 25149
rect 41233 25140 41245 25143
rect 40552 25112 41245 25140
rect 40552 25100 40558 25112
rect 41233 25109 41245 25112
rect 41279 25109 41291 25143
rect 41233 25103 41291 25109
rect 1104 25050 42872 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 42872 25050
rect 1104 24976 42872 24998
rect 14277 24939 14335 24945
rect 14277 24905 14289 24939
rect 14323 24936 14335 24939
rect 14550 24936 14556 24948
rect 14323 24908 14556 24936
rect 14323 24905 14335 24908
rect 14277 24899 14335 24905
rect 14550 24896 14556 24908
rect 14608 24896 14614 24948
rect 16022 24936 16028 24948
rect 15672 24908 16028 24936
rect 15672 24877 15700 24908
rect 16022 24896 16028 24908
rect 16080 24896 16086 24948
rect 25682 24945 25688 24948
rect 25669 24939 25688 24945
rect 25669 24905 25681 24939
rect 25669 24899 25688 24905
rect 25682 24896 25688 24899
rect 25740 24896 25746 24948
rect 26694 24896 26700 24948
rect 26752 24936 26758 24948
rect 27341 24939 27399 24945
rect 27341 24936 27353 24939
rect 26752 24908 27353 24936
rect 26752 24896 26758 24908
rect 27341 24905 27353 24908
rect 27387 24905 27399 24939
rect 27341 24899 27399 24905
rect 28442 24896 28448 24948
rect 28500 24936 28506 24948
rect 28629 24939 28687 24945
rect 28629 24936 28641 24939
rect 28500 24908 28641 24936
rect 28500 24896 28506 24908
rect 28629 24905 28641 24908
rect 28675 24905 28687 24939
rect 29546 24936 29552 24948
rect 29507 24908 29552 24936
rect 28629 24899 28687 24905
rect 29546 24896 29552 24908
rect 29604 24896 29610 24948
rect 31110 24896 31116 24948
rect 31168 24936 31174 24948
rect 31405 24939 31463 24945
rect 31405 24936 31417 24939
rect 31168 24908 31417 24936
rect 31168 24896 31174 24908
rect 31405 24905 31417 24908
rect 31451 24905 31463 24939
rect 31405 24899 31463 24905
rect 31570 24896 31576 24948
rect 31628 24936 31634 24948
rect 33042 24936 33048 24948
rect 31628 24908 33048 24936
rect 31628 24896 31634 24908
rect 33042 24896 33048 24908
rect 33100 24896 33106 24948
rect 15657 24871 15715 24877
rect 15657 24837 15669 24871
rect 15703 24837 15715 24871
rect 15657 24831 15715 24837
rect 15838 24828 15844 24880
rect 15896 24877 15902 24880
rect 15896 24871 15925 24877
rect 15913 24837 15925 24871
rect 15896 24831 15925 24837
rect 25869 24871 25927 24877
rect 25869 24837 25881 24871
rect 25915 24868 25927 24871
rect 27249 24871 27307 24877
rect 27249 24868 27261 24871
rect 25915 24840 27261 24868
rect 25915 24837 25927 24840
rect 25869 24831 25927 24837
rect 27249 24837 27261 24840
rect 27295 24868 27307 24871
rect 27522 24868 27528 24880
rect 27295 24840 27528 24868
rect 27295 24837 27307 24840
rect 27249 24831 27307 24837
rect 15896 24828 15902 24831
rect 27522 24828 27528 24840
rect 27580 24828 27586 24880
rect 30558 24828 30564 24880
rect 30616 24868 30622 24880
rect 31205 24871 31263 24877
rect 31205 24868 31217 24871
rect 30616 24840 31217 24868
rect 30616 24828 30622 24840
rect 31205 24837 31217 24840
rect 31251 24837 31263 24871
rect 33318 24868 33324 24880
rect 31205 24831 31263 24837
rect 32508 24840 33324 24868
rect 12894 24800 12900 24812
rect 12855 24772 12900 24800
rect 12894 24760 12900 24772
rect 12952 24760 12958 24812
rect 13164 24803 13222 24809
rect 13164 24769 13176 24803
rect 13210 24800 13222 24803
rect 13446 24800 13452 24812
rect 13210 24772 13452 24800
rect 13210 24769 13222 24772
rect 13164 24763 13222 24769
rect 13446 24760 13452 24772
rect 13504 24760 13510 24812
rect 14918 24800 14924 24812
rect 14879 24772 14924 24800
rect 14918 24760 14924 24772
rect 14976 24760 14982 24812
rect 15470 24760 15476 24812
rect 15528 24800 15534 24812
rect 15565 24803 15623 24809
rect 15565 24800 15577 24803
rect 15528 24772 15577 24800
rect 15528 24760 15534 24772
rect 15565 24769 15577 24772
rect 15611 24769 15623 24803
rect 15565 24763 15623 24769
rect 15749 24803 15807 24809
rect 15749 24769 15761 24803
rect 15795 24800 15807 24803
rect 16025 24803 16083 24809
rect 15795 24772 15884 24800
rect 15795 24769 15807 24772
rect 15749 24763 15807 24769
rect 14829 24735 14887 24741
rect 14829 24701 14841 24735
rect 14875 24732 14887 24735
rect 15856 24732 15884 24772
rect 16025 24769 16037 24803
rect 16071 24800 16083 24803
rect 16390 24800 16396 24812
rect 16071 24772 16396 24800
rect 16071 24769 16083 24772
rect 16025 24763 16083 24769
rect 16390 24760 16396 24772
rect 16448 24760 16454 24812
rect 17034 24800 17040 24812
rect 16995 24772 17040 24800
rect 17034 24760 17040 24772
rect 17092 24760 17098 24812
rect 17218 24760 17224 24812
rect 17276 24800 17282 24812
rect 17402 24800 17408 24812
rect 17276 24772 17408 24800
rect 17276 24760 17282 24772
rect 17402 24760 17408 24772
rect 17460 24760 17466 24812
rect 18690 24760 18696 24812
rect 18748 24800 18754 24812
rect 19521 24803 19579 24809
rect 19521 24800 19533 24803
rect 18748 24772 19533 24800
rect 18748 24760 18754 24772
rect 19521 24769 19533 24772
rect 19567 24769 19579 24803
rect 19521 24763 19579 24769
rect 19610 24760 19616 24812
rect 19668 24800 19674 24812
rect 19777 24803 19835 24809
rect 19777 24800 19789 24803
rect 19668 24772 19789 24800
rect 19668 24760 19674 24772
rect 19777 24769 19789 24772
rect 19823 24769 19835 24803
rect 19777 24763 19835 24769
rect 22002 24760 22008 24812
rect 22060 24800 22066 24812
rect 22189 24803 22247 24809
rect 22189 24800 22201 24803
rect 22060 24772 22201 24800
rect 22060 24760 22066 24772
rect 22189 24769 22201 24772
rect 22235 24769 22247 24803
rect 22189 24763 22247 24769
rect 23017 24803 23075 24809
rect 23017 24769 23029 24803
rect 23063 24800 23075 24803
rect 23382 24800 23388 24812
rect 23063 24772 23388 24800
rect 23063 24769 23075 24772
rect 23017 24763 23075 24769
rect 23382 24760 23388 24772
rect 23440 24760 23446 24812
rect 27154 24800 27160 24812
rect 27115 24772 27160 24800
rect 27154 24760 27160 24772
rect 27212 24760 27218 24812
rect 28813 24803 28871 24809
rect 28813 24769 28825 24803
rect 28859 24769 28871 24803
rect 29362 24800 29368 24812
rect 29323 24772 29368 24800
rect 28813 24763 28871 24769
rect 15930 24732 15936 24744
rect 14875 24704 15936 24732
rect 14875 24701 14887 24704
rect 14829 24695 14887 24701
rect 15930 24692 15936 24704
rect 15988 24692 15994 24744
rect 17126 24692 17132 24744
rect 17184 24732 17190 24744
rect 17313 24735 17371 24741
rect 17313 24732 17325 24735
rect 17184 24704 17325 24732
rect 17184 24692 17190 24704
rect 17313 24701 17325 24704
rect 17359 24701 17371 24735
rect 17313 24695 17371 24701
rect 21266 24692 21272 24744
rect 21324 24732 21330 24744
rect 22281 24735 22339 24741
rect 22281 24732 22293 24735
rect 21324 24704 22293 24732
rect 21324 24692 21330 24704
rect 22281 24701 22293 24704
rect 22327 24732 22339 24735
rect 22462 24732 22468 24744
rect 22327 24704 22468 24732
rect 22327 24701 22339 24704
rect 22281 24695 22339 24701
rect 22462 24692 22468 24704
rect 22520 24732 22526 24744
rect 25314 24732 25320 24744
rect 22520 24704 25320 24732
rect 22520 24692 22526 24704
rect 25314 24692 25320 24704
rect 25372 24692 25378 24744
rect 26602 24692 26608 24744
rect 26660 24732 26666 24744
rect 26973 24735 27031 24741
rect 26973 24732 26985 24735
rect 26660 24704 26985 24732
rect 26660 24692 26666 24704
rect 26973 24701 26985 24704
rect 27019 24701 27031 24735
rect 28828 24732 28856 24763
rect 29362 24760 29368 24772
rect 29420 24760 29426 24812
rect 30742 24732 30748 24744
rect 28828 24704 30748 24732
rect 26973 24695 27031 24701
rect 30742 24692 30748 24704
rect 30800 24692 30806 24744
rect 31220 24732 31248 24831
rect 32508 24812 32536 24840
rect 33318 24828 33324 24840
rect 33376 24828 33382 24880
rect 40218 24868 40224 24880
rect 36280 24840 36584 24868
rect 40179 24840 40224 24868
rect 31754 24760 31760 24812
rect 31812 24800 31818 24812
rect 32306 24800 32312 24812
rect 31812 24772 32312 24800
rect 31812 24760 31818 24772
rect 32306 24760 32312 24772
rect 32364 24760 32370 24812
rect 32493 24806 32551 24812
rect 32493 24772 32505 24806
rect 32539 24772 32551 24806
rect 32493 24766 32551 24772
rect 32588 24803 32646 24809
rect 32588 24769 32600 24803
rect 32634 24769 32646 24803
rect 32588 24763 32646 24769
rect 32677 24803 32735 24809
rect 32677 24769 32689 24803
rect 32723 24769 32735 24803
rect 34526 24803 34584 24809
rect 34526 24800 34538 24803
rect 32677 24763 32735 24769
rect 32968 24772 34538 24800
rect 31570 24732 31576 24744
rect 31220 24704 31576 24732
rect 31570 24692 31576 24704
rect 31628 24692 31634 24744
rect 32398 24692 32404 24744
rect 32456 24732 32462 24744
rect 32600 24732 32628 24763
rect 32456 24704 32628 24732
rect 32692 24732 32720 24763
rect 32766 24732 32772 24744
rect 32692 24704 32772 24732
rect 32456 24692 32462 24704
rect 32766 24692 32772 24704
rect 32824 24692 32830 24744
rect 32968 24741 32996 24772
rect 34526 24769 34538 24772
rect 34572 24769 34584 24803
rect 34526 24763 34584 24769
rect 34698 24760 34704 24812
rect 34756 24800 34762 24812
rect 34793 24803 34851 24809
rect 34793 24800 34805 24803
rect 34756 24772 34805 24800
rect 34756 24760 34762 24772
rect 34793 24769 34805 24772
rect 34839 24800 34851 24803
rect 36280 24800 36308 24840
rect 34839 24772 36308 24800
rect 34839 24769 34851 24772
rect 34793 24763 34851 24769
rect 36354 24760 36360 24812
rect 36412 24809 36418 24812
rect 36412 24800 36424 24809
rect 36556 24800 36584 24840
rect 40218 24828 40224 24840
rect 40276 24828 40282 24880
rect 36633 24803 36691 24809
rect 36633 24800 36645 24803
rect 36412 24772 36457 24800
rect 36556 24772 36645 24800
rect 36412 24763 36424 24772
rect 36633 24769 36645 24772
rect 36679 24769 36691 24803
rect 39298 24800 39304 24812
rect 39259 24772 39304 24800
rect 36633 24763 36691 24769
rect 36412 24760 36418 24763
rect 39298 24760 39304 24772
rect 39356 24760 39362 24812
rect 40034 24800 40040 24812
rect 39995 24772 40040 24800
rect 40034 24760 40040 24772
rect 40092 24760 40098 24812
rect 32953 24735 33011 24741
rect 32953 24701 32965 24735
rect 32999 24701 33011 24735
rect 32953 24695 33011 24701
rect 33042 24692 33048 24744
rect 33100 24732 33106 24744
rect 41230 24732 41236 24744
rect 33100 24704 33548 24732
rect 41191 24704 41236 24732
rect 33100 24692 33106 24704
rect 13906 24624 13912 24676
rect 13964 24664 13970 24676
rect 15381 24667 15439 24673
rect 15381 24664 15393 24667
rect 13964 24636 15393 24664
rect 13964 24624 13970 24636
rect 15381 24633 15393 24636
rect 15427 24633 15439 24667
rect 17497 24667 17555 24673
rect 15381 24627 15439 24633
rect 15488 24636 17264 24664
rect 13814 24556 13820 24608
rect 13872 24596 13878 24608
rect 14182 24596 14188 24608
rect 13872 24568 14188 24596
rect 13872 24556 13878 24568
rect 14182 24556 14188 24568
rect 14240 24596 14246 24608
rect 15488 24596 15516 24636
rect 14240 24568 15516 24596
rect 14240 24556 14246 24568
rect 16758 24556 16764 24608
rect 16816 24596 16822 24608
rect 17129 24599 17187 24605
rect 17129 24596 17141 24599
rect 16816 24568 17141 24596
rect 16816 24556 16822 24568
rect 17129 24565 17141 24568
rect 17175 24565 17187 24599
rect 17236 24596 17264 24636
rect 17497 24633 17509 24667
rect 17543 24664 17555 24667
rect 17954 24664 17960 24676
rect 17543 24636 17960 24664
rect 17543 24633 17555 24636
rect 17497 24627 17555 24633
rect 17954 24624 17960 24636
rect 18012 24624 18018 24676
rect 25038 24624 25044 24676
rect 25096 24664 25102 24676
rect 25501 24667 25559 24673
rect 25501 24664 25513 24667
rect 25096 24636 25513 24664
rect 25096 24624 25102 24636
rect 25501 24633 25513 24636
rect 25547 24633 25559 24667
rect 25501 24627 25559 24633
rect 27430 24624 27436 24676
rect 27488 24664 27494 24676
rect 27525 24667 27583 24673
rect 27525 24664 27537 24667
rect 27488 24636 27537 24664
rect 27488 24624 27494 24636
rect 27525 24633 27537 24636
rect 27571 24633 27583 24667
rect 27525 24627 27583 24633
rect 18598 24596 18604 24608
rect 17236 24568 18604 24596
rect 17129 24559 17187 24565
rect 18598 24556 18604 24568
rect 18656 24556 18662 24608
rect 20898 24596 20904 24608
rect 20859 24568 20904 24596
rect 20898 24556 20904 24568
rect 20956 24556 20962 24608
rect 22554 24596 22560 24608
rect 22515 24568 22560 24596
rect 22554 24556 22560 24568
rect 22612 24556 22618 24608
rect 23198 24596 23204 24608
rect 23159 24568 23204 24596
rect 23198 24556 23204 24568
rect 23256 24556 23262 24608
rect 25685 24599 25743 24605
rect 25685 24565 25697 24599
rect 25731 24596 25743 24599
rect 26234 24596 26240 24608
rect 25731 24568 26240 24596
rect 25731 24565 25743 24568
rect 25685 24559 25743 24565
rect 26234 24556 26240 24568
rect 26292 24556 26298 24608
rect 31294 24556 31300 24608
rect 31352 24596 31358 24608
rect 31389 24599 31447 24605
rect 31389 24596 31401 24599
rect 31352 24568 31401 24596
rect 31352 24556 31358 24568
rect 31389 24565 31401 24568
rect 31435 24565 31447 24599
rect 31389 24559 31447 24565
rect 31478 24556 31484 24608
rect 31536 24596 31542 24608
rect 31573 24599 31631 24605
rect 31573 24596 31585 24599
rect 31536 24568 31585 24596
rect 31536 24556 31542 24568
rect 31573 24565 31585 24568
rect 31619 24565 31631 24599
rect 31573 24559 31631 24565
rect 33226 24556 33232 24608
rect 33284 24596 33290 24608
rect 33413 24599 33471 24605
rect 33413 24596 33425 24599
rect 33284 24568 33425 24596
rect 33284 24556 33290 24568
rect 33413 24565 33425 24568
rect 33459 24565 33471 24599
rect 33520 24596 33548 24704
rect 41230 24692 41236 24704
rect 41288 24692 41294 24744
rect 35253 24599 35311 24605
rect 35253 24596 35265 24599
rect 33520 24568 35265 24596
rect 33413 24559 33471 24565
rect 35253 24565 35265 24568
rect 35299 24565 35311 24599
rect 35253 24559 35311 24565
rect 39485 24599 39543 24605
rect 39485 24565 39497 24599
rect 39531 24596 39543 24599
rect 40034 24596 40040 24608
rect 39531 24568 40040 24596
rect 39531 24565 39543 24568
rect 39485 24559 39543 24565
rect 40034 24556 40040 24568
rect 40092 24556 40098 24608
rect 1104 24506 42872 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 42872 24506
rect 1104 24432 42872 24454
rect 13446 24392 13452 24404
rect 13407 24364 13452 24392
rect 13446 24352 13452 24364
rect 13504 24352 13510 24404
rect 14826 24352 14832 24404
rect 14884 24352 14890 24404
rect 15013 24395 15071 24401
rect 15013 24361 15025 24395
rect 15059 24392 15071 24395
rect 15286 24392 15292 24404
rect 15059 24364 15292 24392
rect 15059 24361 15071 24364
rect 15013 24355 15071 24361
rect 15286 24352 15292 24364
rect 15344 24352 15350 24404
rect 15562 24392 15568 24404
rect 15523 24364 15568 24392
rect 15562 24352 15568 24364
rect 15620 24352 15626 24404
rect 17126 24392 17132 24404
rect 17087 24364 17132 24392
rect 17126 24352 17132 24364
rect 17184 24352 17190 24404
rect 19610 24392 19616 24404
rect 19571 24364 19616 24392
rect 19610 24352 19616 24364
rect 19668 24352 19674 24404
rect 20806 24392 20812 24404
rect 20767 24364 20812 24392
rect 20806 24352 20812 24364
rect 20864 24352 20870 24404
rect 23382 24392 23388 24404
rect 23343 24364 23388 24392
rect 23382 24352 23388 24364
rect 23440 24352 23446 24404
rect 29638 24352 29644 24404
rect 29696 24392 29702 24404
rect 29733 24395 29791 24401
rect 29733 24392 29745 24395
rect 29696 24364 29745 24392
rect 29696 24352 29702 24364
rect 29733 24361 29745 24364
rect 29779 24361 29791 24395
rect 29733 24355 29791 24361
rect 30561 24395 30619 24401
rect 30561 24361 30573 24395
rect 30607 24392 30619 24395
rect 30650 24392 30656 24404
rect 30607 24364 30656 24392
rect 30607 24361 30619 24364
rect 30561 24355 30619 24361
rect 30650 24352 30656 24364
rect 30708 24352 30714 24404
rect 31478 24392 31484 24404
rect 31439 24364 31484 24392
rect 31478 24352 31484 24364
rect 31536 24392 31542 24404
rect 32674 24392 32680 24404
rect 31536 24364 32352 24392
rect 32635 24364 32680 24392
rect 31536 24352 31542 24364
rect 14844 24324 14872 24352
rect 14200 24296 20300 24324
rect 3602 24216 3608 24268
rect 3660 24256 3666 24268
rect 3789 24259 3847 24265
rect 3789 24256 3801 24259
rect 3660 24228 3801 24256
rect 3660 24216 3666 24228
rect 3789 24225 3801 24228
rect 3835 24225 3847 24259
rect 5626 24256 5632 24268
rect 5587 24228 5632 24256
rect 3789 24219 3847 24225
rect 5626 24216 5632 24228
rect 5684 24216 5690 24268
rect 13814 24256 13820 24268
rect 13372 24228 13820 24256
rect 13372 24197 13400 24228
rect 13814 24216 13820 24228
rect 13872 24216 13878 24268
rect 14200 24256 14228 24296
rect 14108 24228 14228 24256
rect 14829 24259 14887 24265
rect 13357 24191 13415 24197
rect 13357 24157 13369 24191
rect 13403 24157 13415 24191
rect 13357 24151 13415 24157
rect 13541 24191 13599 24197
rect 13541 24157 13553 24191
rect 13587 24188 13599 24191
rect 13906 24188 13912 24200
rect 13587 24160 13912 24188
rect 13587 24157 13599 24160
rect 13541 24151 13599 24157
rect 13906 24148 13912 24160
rect 13964 24148 13970 24200
rect 14108 24197 14136 24228
rect 14829 24225 14841 24259
rect 14875 24256 14887 24259
rect 14918 24256 14924 24268
rect 14875 24228 14924 24256
rect 14875 24225 14887 24228
rect 14829 24219 14887 24225
rect 14918 24216 14924 24228
rect 14976 24256 14982 24268
rect 17126 24256 17132 24268
rect 14976 24228 15792 24256
rect 14976 24216 14982 24228
rect 14093 24191 14151 24197
rect 14093 24157 14105 24191
rect 14139 24157 14151 24191
rect 14093 24151 14151 24157
rect 14185 24191 14243 24197
rect 14185 24157 14197 24191
rect 14231 24188 14243 24191
rect 15105 24191 15163 24197
rect 14231 24160 14872 24188
rect 14231 24157 14243 24160
rect 14185 24151 14243 24157
rect 3418 24080 3424 24132
rect 3476 24120 3482 24132
rect 14844 24129 14872 24160
rect 15105 24157 15117 24191
rect 15151 24188 15163 24191
rect 15151 24160 15608 24188
rect 15151 24157 15163 24160
rect 15105 24151 15163 24157
rect 5445 24123 5503 24129
rect 5445 24120 5457 24123
rect 3476 24092 5457 24120
rect 3476 24080 3482 24092
rect 5445 24089 5457 24092
rect 5491 24089 5503 24123
rect 5445 24083 5503 24089
rect 14369 24123 14427 24129
rect 14369 24089 14381 24123
rect 14415 24120 14427 24123
rect 14829 24123 14887 24129
rect 14415 24092 14780 24120
rect 14415 24089 14427 24092
rect 14369 24083 14427 24089
rect 14277 24055 14335 24061
rect 14277 24021 14289 24055
rect 14323 24052 14335 24055
rect 14458 24052 14464 24064
rect 14323 24024 14464 24052
rect 14323 24021 14335 24024
rect 14277 24015 14335 24021
rect 14458 24012 14464 24024
rect 14516 24012 14522 24064
rect 14752 24052 14780 24092
rect 14829 24089 14841 24123
rect 14875 24089 14887 24123
rect 14829 24083 14887 24089
rect 15194 24052 15200 24064
rect 14752 24024 15200 24052
rect 15194 24012 15200 24024
rect 15252 24012 15258 24064
rect 15580 24052 15608 24160
rect 15764 24132 15792 24228
rect 15948 24228 17132 24256
rect 15948 24197 15976 24228
rect 17126 24216 17132 24228
rect 17184 24256 17190 24268
rect 17221 24259 17279 24265
rect 17221 24256 17233 24259
rect 17184 24228 17233 24256
rect 17184 24216 17190 24228
rect 17221 24225 17233 24228
rect 17267 24225 17279 24259
rect 17221 24219 17279 24225
rect 18138 24216 18144 24268
rect 18196 24256 18202 24268
rect 18417 24259 18475 24265
rect 18417 24256 18429 24259
rect 18196 24228 18429 24256
rect 18196 24216 18202 24228
rect 18417 24225 18429 24228
rect 18463 24225 18475 24259
rect 20162 24256 20168 24268
rect 18417 24219 18475 24225
rect 19904 24228 20168 24256
rect 15933 24191 15991 24197
rect 15933 24157 15945 24191
rect 15979 24157 15991 24191
rect 16942 24188 16948 24200
rect 16903 24160 16948 24188
rect 15933 24151 15991 24157
rect 15746 24120 15752 24132
rect 15707 24092 15752 24120
rect 15746 24080 15752 24092
rect 15804 24080 15810 24132
rect 15948 24052 15976 24151
rect 16942 24148 16948 24160
rect 17000 24148 17006 24200
rect 19904 24197 19932 24228
rect 20162 24216 20168 24228
rect 20220 24216 20226 24268
rect 17037 24191 17095 24197
rect 17037 24157 17049 24191
rect 17083 24157 17095 24191
rect 17037 24151 17095 24157
rect 18233 24191 18291 24197
rect 18233 24157 18245 24191
rect 18279 24157 18291 24191
rect 18233 24151 18291 24157
rect 19889 24191 19947 24197
rect 19889 24157 19901 24191
rect 19935 24157 19947 24191
rect 19889 24151 19947 24157
rect 19981 24191 20039 24197
rect 19981 24157 19993 24191
rect 20027 24157 20039 24191
rect 19981 24151 20039 24157
rect 16758 24080 16764 24132
rect 16816 24120 16822 24132
rect 17052 24120 17080 24151
rect 16816 24092 17080 24120
rect 18248 24120 18276 24151
rect 19426 24120 19432 24132
rect 18248 24092 19432 24120
rect 16816 24080 16822 24092
rect 19426 24080 19432 24092
rect 19484 24080 19490 24132
rect 19996 24120 20024 24151
rect 20070 24148 20076 24200
rect 20128 24188 20134 24200
rect 20272 24197 20300 24296
rect 20898 24284 20904 24336
rect 20956 24324 20962 24336
rect 21174 24324 21180 24336
rect 20956 24296 21180 24324
rect 20956 24284 20962 24296
rect 21174 24284 21180 24296
rect 21232 24324 21238 24336
rect 21545 24327 21603 24333
rect 21545 24324 21557 24327
rect 21232 24296 21557 24324
rect 21232 24284 21238 24296
rect 21545 24293 21557 24296
rect 21591 24293 21603 24327
rect 21545 24287 21603 24293
rect 26237 24327 26295 24333
rect 26237 24293 26249 24327
rect 26283 24324 26295 24327
rect 26326 24324 26332 24336
rect 26283 24296 26332 24324
rect 26283 24293 26295 24296
rect 26237 24287 26295 24293
rect 26326 24284 26332 24296
rect 26384 24284 26390 24336
rect 28997 24327 29055 24333
rect 28997 24293 29009 24327
rect 29043 24324 29055 24327
rect 29270 24324 29276 24336
rect 29043 24296 29276 24324
rect 29043 24293 29055 24296
rect 28997 24287 29055 24293
rect 29270 24284 29276 24296
rect 29328 24284 29334 24336
rect 32324 24333 32352 24364
rect 32674 24352 32680 24364
rect 32732 24352 32738 24404
rect 33321 24395 33379 24401
rect 33321 24361 33333 24395
rect 33367 24392 33379 24395
rect 33410 24392 33416 24404
rect 33367 24364 33416 24392
rect 33367 24361 33379 24364
rect 33321 24355 33379 24361
rect 33410 24352 33416 24364
rect 33468 24352 33474 24404
rect 34149 24395 34207 24401
rect 34149 24361 34161 24395
rect 34195 24392 34207 24395
rect 36354 24392 36360 24404
rect 34195 24364 36360 24392
rect 34195 24361 34207 24364
rect 34149 24355 34207 24361
rect 36354 24352 36360 24364
rect 36412 24352 36418 24404
rect 32309 24327 32367 24333
rect 32309 24293 32321 24327
rect 32355 24293 32367 24327
rect 32309 24287 32367 24293
rect 32861 24327 32919 24333
rect 32861 24293 32873 24327
rect 32907 24293 32919 24327
rect 37550 24324 37556 24336
rect 37511 24296 37556 24324
rect 32861 24287 32919 24293
rect 20622 24216 20628 24268
rect 20680 24256 20686 24268
rect 20993 24259 21051 24265
rect 20993 24256 21005 24259
rect 20680 24228 21005 24256
rect 20680 24216 20686 24228
rect 20993 24225 21005 24228
rect 21039 24225 21051 24259
rect 23750 24256 23756 24268
rect 23711 24228 23756 24256
rect 20993 24219 21051 24225
rect 23750 24216 23756 24228
rect 23808 24256 23814 24268
rect 24026 24256 24032 24268
rect 23808 24228 24032 24256
rect 23808 24216 23814 24228
rect 24026 24216 24032 24228
rect 24084 24216 24090 24268
rect 24673 24259 24731 24265
rect 24673 24225 24685 24259
rect 24719 24256 24731 24259
rect 25590 24256 25596 24268
rect 24719 24228 25596 24256
rect 24719 24225 24731 24228
rect 24673 24219 24731 24225
rect 25590 24216 25596 24228
rect 25648 24216 25654 24268
rect 26789 24259 26847 24265
rect 26789 24225 26801 24259
rect 26835 24256 26847 24259
rect 27154 24256 27160 24268
rect 26835 24228 27160 24256
rect 26835 24225 26847 24228
rect 26789 24219 26847 24225
rect 27154 24216 27160 24228
rect 27212 24256 27218 24268
rect 28534 24256 28540 24268
rect 27212 24228 28540 24256
rect 27212 24216 27218 24228
rect 28534 24216 28540 24228
rect 28592 24216 28598 24268
rect 31573 24259 31631 24265
rect 31573 24256 31585 24259
rect 30668 24228 31585 24256
rect 20257 24191 20315 24197
rect 20128 24160 20173 24188
rect 20128 24148 20134 24160
rect 20257 24157 20269 24191
rect 20303 24157 20315 24191
rect 20257 24151 20315 24157
rect 20806 24148 20812 24200
rect 20864 24188 20870 24200
rect 22097 24191 22155 24197
rect 22097 24188 22109 24191
rect 20864 24160 22109 24188
rect 20864 24148 20870 24160
rect 22097 24157 22109 24160
rect 22143 24157 22155 24191
rect 22370 24188 22376 24200
rect 22331 24160 22376 24188
rect 22097 24151 22155 24157
rect 22370 24148 22376 24160
rect 22428 24148 22434 24200
rect 22554 24148 22560 24200
rect 22612 24188 22618 24200
rect 23569 24191 23627 24197
rect 23569 24188 23581 24191
rect 22612 24160 23581 24188
rect 22612 24148 22618 24160
rect 23569 24157 23581 24160
rect 23615 24157 23627 24191
rect 24394 24188 24400 24200
rect 24355 24160 24400 24188
rect 23569 24151 23627 24157
rect 24394 24148 24400 24160
rect 24452 24148 24458 24200
rect 24486 24148 24492 24200
rect 24544 24188 24550 24200
rect 24544 24160 24589 24188
rect 24544 24148 24550 24160
rect 25682 24148 25688 24200
rect 25740 24188 25746 24200
rect 26053 24191 26111 24197
rect 26053 24188 26065 24191
rect 25740 24160 26065 24188
rect 25740 24148 25746 24160
rect 26053 24157 26065 24160
rect 26099 24157 26111 24191
rect 26053 24151 26111 24157
rect 26234 24148 26240 24200
rect 26292 24188 26298 24200
rect 26697 24191 26755 24197
rect 26697 24188 26709 24191
rect 26292 24160 26709 24188
rect 26292 24148 26298 24160
rect 26697 24157 26709 24160
rect 26743 24157 26755 24191
rect 26697 24151 26755 24157
rect 28258 24148 28264 24200
rect 28316 24188 28322 24200
rect 28718 24188 28724 24200
rect 28316 24160 28724 24188
rect 28316 24148 28322 24160
rect 28718 24148 28724 24160
rect 28776 24148 28782 24200
rect 28813 24191 28871 24197
rect 28813 24157 28825 24191
rect 28859 24188 28871 24191
rect 30374 24188 30380 24200
rect 28859 24160 30380 24188
rect 28859 24157 28871 24160
rect 28813 24151 28871 24157
rect 30374 24148 30380 24160
rect 30432 24148 30438 24200
rect 30469 24191 30527 24197
rect 30469 24157 30481 24191
rect 30515 24188 30527 24191
rect 30558 24188 30564 24200
rect 30515 24160 30564 24188
rect 30515 24157 30527 24160
rect 30469 24151 30527 24157
rect 30558 24148 30564 24160
rect 30616 24148 30622 24200
rect 30668 24197 30696 24228
rect 31573 24225 31585 24228
rect 31619 24256 31631 24259
rect 32876 24256 32904 24287
rect 37550 24284 37556 24296
rect 37608 24284 37614 24336
rect 40034 24256 40040 24268
rect 31619 24228 31754 24256
rect 32876 24228 34008 24256
rect 39995 24228 40040 24256
rect 31619 24225 31631 24228
rect 31573 24219 31631 24225
rect 31726 24200 31754 24228
rect 30653 24191 30711 24197
rect 30653 24157 30665 24191
rect 30699 24157 30711 24191
rect 31294 24188 31300 24200
rect 31255 24160 31300 24188
rect 30653 24151 30711 24157
rect 31294 24148 31300 24160
rect 31352 24148 31358 24200
rect 31726 24160 31760 24200
rect 31754 24148 31760 24160
rect 31812 24148 31818 24200
rect 33226 24148 33232 24200
rect 33284 24188 33290 24200
rect 33980 24197 34008 24228
rect 40034 24216 40040 24228
rect 40092 24216 40098 24268
rect 40402 24216 40408 24268
rect 40460 24256 40466 24268
rect 40497 24259 40555 24265
rect 40497 24256 40509 24259
rect 40460 24228 40509 24256
rect 40460 24216 40466 24228
rect 40497 24225 40509 24228
rect 40543 24225 40555 24259
rect 40497 24219 40555 24225
rect 33505 24191 33563 24197
rect 33505 24188 33517 24191
rect 33284 24160 33517 24188
rect 33284 24148 33290 24160
rect 33505 24157 33517 24160
rect 33551 24157 33563 24191
rect 33505 24151 33563 24157
rect 33965 24191 34023 24197
rect 33965 24157 33977 24191
rect 34011 24157 34023 24191
rect 33965 24151 34023 24157
rect 37737 24191 37795 24197
rect 37737 24157 37749 24191
rect 37783 24188 37795 24191
rect 38654 24188 38660 24200
rect 37783 24160 38660 24188
rect 37783 24157 37795 24160
rect 37737 24151 37795 24157
rect 38654 24148 38660 24160
rect 38712 24148 38718 24200
rect 39114 24188 39120 24200
rect 39075 24160 39120 24188
rect 39114 24148 39120 24160
rect 39172 24148 39178 24200
rect 21545 24123 21603 24129
rect 19996 24092 20852 24120
rect 20824 24064 20852 24092
rect 21545 24089 21557 24123
rect 21591 24120 21603 24123
rect 22002 24120 22008 24132
rect 21591 24092 22008 24120
rect 21591 24089 21603 24092
rect 21545 24083 21603 24089
rect 22002 24080 22008 24092
rect 22060 24080 22066 24132
rect 26970 24080 26976 24132
rect 27028 24120 27034 24132
rect 28166 24120 28172 24132
rect 27028 24092 28172 24120
rect 27028 24080 27034 24092
rect 28166 24080 28172 24092
rect 28224 24120 28230 24132
rect 28902 24120 28908 24132
rect 28224 24092 28908 24120
rect 28224 24080 28230 24092
rect 28902 24080 28908 24092
rect 28960 24120 28966 24132
rect 28997 24123 29055 24129
rect 28997 24120 29009 24123
rect 28960 24092 29009 24120
rect 28960 24080 28966 24092
rect 28997 24089 29009 24092
rect 29043 24089 29055 24123
rect 28997 24083 29055 24089
rect 29178 24080 29184 24132
rect 29236 24120 29242 24132
rect 29549 24123 29607 24129
rect 29549 24120 29561 24123
rect 29236 24092 29561 24120
rect 29236 24080 29242 24092
rect 29549 24089 29561 24092
rect 29595 24089 29607 24123
rect 29549 24083 29607 24089
rect 32306 24080 32312 24132
rect 32364 24120 32370 24132
rect 32677 24123 32735 24129
rect 32677 24120 32689 24123
rect 32364 24092 32689 24120
rect 32364 24080 32370 24092
rect 32677 24089 32689 24092
rect 32723 24089 32735 24123
rect 32677 24083 32735 24089
rect 39209 24123 39267 24129
rect 39209 24089 39221 24123
rect 39255 24120 39267 24123
rect 40221 24123 40279 24129
rect 40221 24120 40233 24123
rect 39255 24092 40233 24120
rect 39255 24089 39267 24092
rect 39209 24083 39267 24089
rect 40221 24089 40233 24092
rect 40267 24089 40279 24123
rect 40221 24083 40279 24089
rect 18046 24052 18052 24064
rect 15580 24024 15976 24052
rect 18007 24024 18052 24052
rect 18046 24012 18052 24024
rect 18104 24012 18110 24064
rect 20806 24012 20812 24064
rect 20864 24012 20870 24064
rect 21082 24012 21088 24064
rect 21140 24052 21146 24064
rect 24670 24052 24676 24064
rect 21140 24024 21185 24052
rect 24631 24024 24676 24052
rect 21140 24012 21146 24024
rect 24670 24012 24676 24024
rect 24728 24012 24734 24064
rect 28350 24012 28356 24064
rect 28408 24052 28414 24064
rect 29362 24052 29368 24064
rect 28408 24024 29368 24052
rect 28408 24012 28414 24024
rect 29362 24012 29368 24024
rect 29420 24012 29426 24064
rect 29454 24012 29460 24064
rect 29512 24052 29518 24064
rect 29749 24055 29807 24061
rect 29749 24052 29761 24055
rect 29512 24024 29761 24052
rect 29512 24012 29518 24024
rect 29749 24021 29761 24024
rect 29795 24021 29807 24055
rect 29749 24015 29807 24021
rect 29917 24055 29975 24061
rect 29917 24021 29929 24055
rect 29963 24052 29975 24055
rect 30926 24052 30932 24064
rect 29963 24024 30932 24052
rect 29963 24021 29975 24024
rect 29917 24015 29975 24021
rect 30926 24012 30932 24024
rect 30984 24012 30990 24064
rect 31110 24052 31116 24064
rect 31071 24024 31116 24052
rect 31110 24012 31116 24024
rect 31168 24012 31174 24064
rect 1104 23962 42872 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 42872 23962
rect 1104 23888 42872 23910
rect 3418 23848 3424 23860
rect 3379 23820 3424 23848
rect 3418 23808 3424 23820
rect 3476 23808 3482 23860
rect 16022 23808 16028 23860
rect 16080 23848 16086 23860
rect 16761 23851 16819 23857
rect 16761 23848 16773 23851
rect 16080 23820 16773 23848
rect 16080 23808 16086 23820
rect 16761 23817 16773 23820
rect 16807 23817 16819 23851
rect 16761 23811 16819 23817
rect 20070 23808 20076 23860
rect 20128 23848 20134 23860
rect 20717 23851 20775 23857
rect 20717 23848 20729 23851
rect 20128 23820 20729 23848
rect 20128 23808 20134 23820
rect 20717 23817 20729 23820
rect 20763 23817 20775 23851
rect 20717 23811 20775 23817
rect 21542 23808 21548 23860
rect 21600 23848 21606 23860
rect 22189 23851 22247 23857
rect 22189 23848 22201 23851
rect 21600 23820 22201 23848
rect 21600 23808 21606 23820
rect 22189 23817 22201 23820
rect 22235 23848 22247 23851
rect 22370 23848 22376 23860
rect 22235 23820 22376 23848
rect 22235 23817 22247 23820
rect 22189 23811 22247 23817
rect 22370 23808 22376 23820
rect 22428 23808 22434 23860
rect 24394 23808 24400 23860
rect 24452 23848 24458 23860
rect 24489 23851 24547 23857
rect 24489 23848 24501 23851
rect 24452 23820 24501 23848
rect 24452 23808 24458 23820
rect 24489 23817 24501 23820
rect 24535 23817 24547 23851
rect 25590 23848 25596 23860
rect 25551 23820 25596 23848
rect 24489 23811 24547 23817
rect 25590 23808 25596 23820
rect 25648 23808 25654 23860
rect 27338 23808 27344 23860
rect 27396 23848 27402 23860
rect 27396 23820 28488 23848
rect 27396 23808 27402 23820
rect 21266 23780 21272 23792
rect 20916 23752 21272 23780
rect 3326 23712 3332 23724
rect 3287 23684 3332 23712
rect 3326 23672 3332 23684
rect 3384 23672 3390 23724
rect 14458 23672 14464 23724
rect 14516 23712 14522 23724
rect 14625 23715 14683 23721
rect 14625 23712 14637 23715
rect 14516 23684 14637 23712
rect 14516 23672 14522 23684
rect 14625 23681 14637 23684
rect 14671 23681 14683 23715
rect 14625 23675 14683 23681
rect 16853 23715 16911 23721
rect 16853 23681 16865 23715
rect 16899 23712 16911 23715
rect 17034 23712 17040 23724
rect 16899 23684 17040 23712
rect 16899 23681 16911 23684
rect 16853 23675 16911 23681
rect 17034 23672 17040 23684
rect 17092 23672 17098 23724
rect 17678 23721 17684 23724
rect 17672 23675 17684 23721
rect 17736 23712 17742 23724
rect 19429 23715 19487 23721
rect 17736 23684 17772 23712
rect 17678 23672 17684 23675
rect 17736 23672 17742 23684
rect 19429 23681 19441 23715
rect 19475 23712 19487 23715
rect 20622 23712 20628 23724
rect 19475 23684 20628 23712
rect 19475 23681 19487 23684
rect 19429 23675 19487 23681
rect 14366 23644 14372 23656
rect 14327 23616 14372 23644
rect 14366 23604 14372 23616
rect 14424 23604 14430 23656
rect 16666 23604 16672 23656
rect 16724 23644 16730 23656
rect 17405 23647 17463 23653
rect 17405 23644 17417 23647
rect 16724 23616 17417 23644
rect 16724 23604 16730 23616
rect 17405 23613 17417 23616
rect 17451 23613 17463 23647
rect 17405 23607 17463 23613
rect 15746 23576 15752 23588
rect 15707 23548 15752 23576
rect 15746 23536 15752 23548
rect 15804 23536 15810 23588
rect 18785 23579 18843 23585
rect 18785 23545 18797 23579
rect 18831 23576 18843 23579
rect 19444 23576 19472 23675
rect 20622 23672 20628 23684
rect 20680 23672 20686 23724
rect 20714 23672 20720 23724
rect 20772 23712 20778 23724
rect 20916 23721 20944 23752
rect 21266 23740 21272 23752
rect 21324 23740 21330 23792
rect 23198 23740 23204 23792
rect 23256 23780 23262 23792
rect 23354 23783 23412 23789
rect 23354 23780 23366 23783
rect 23256 23752 23366 23780
rect 23256 23740 23262 23752
rect 23354 23749 23366 23752
rect 23400 23749 23412 23783
rect 23354 23743 23412 23749
rect 24670 23740 24676 23792
rect 24728 23780 24734 23792
rect 24728 23752 28304 23780
rect 24728 23740 24734 23752
rect 20901 23715 20959 23721
rect 20901 23712 20913 23715
rect 20772 23684 20913 23712
rect 20772 23672 20778 23684
rect 20901 23681 20913 23684
rect 20947 23681 20959 23715
rect 20901 23675 20959 23681
rect 20993 23715 21051 23721
rect 20993 23681 21005 23715
rect 21039 23712 21051 23715
rect 21039 23684 22048 23712
rect 21039 23681 21051 23684
rect 20993 23675 21051 23681
rect 22020 23656 22048 23684
rect 23842 23672 23848 23724
rect 23900 23712 23906 23724
rect 24949 23715 25007 23721
rect 24949 23712 24961 23715
rect 23900 23684 24961 23712
rect 23900 23672 23906 23684
rect 24949 23681 24961 23684
rect 24995 23681 25007 23715
rect 25130 23712 25136 23724
rect 25091 23684 25136 23712
rect 24949 23675 25007 23681
rect 25130 23672 25136 23684
rect 25188 23672 25194 23724
rect 25409 23715 25467 23721
rect 25409 23681 25421 23715
rect 25455 23712 25467 23715
rect 26053 23715 26111 23721
rect 26053 23712 26065 23715
rect 25455 23684 26065 23712
rect 25455 23681 25467 23684
rect 25409 23675 25467 23681
rect 26053 23681 26065 23684
rect 26099 23712 26111 23715
rect 26421 23715 26479 23721
rect 26099 23684 26372 23712
rect 26099 23681 26111 23684
rect 26053 23675 26111 23681
rect 19521 23647 19579 23653
rect 19521 23613 19533 23647
rect 19567 23644 19579 23647
rect 20806 23644 20812 23656
rect 19567 23616 20812 23644
rect 19567 23613 19579 23616
rect 19521 23607 19579 23613
rect 20806 23604 20812 23616
rect 20864 23604 20870 23656
rect 21082 23644 21088 23656
rect 20995 23616 21088 23644
rect 21082 23604 21088 23616
rect 21140 23604 21146 23656
rect 21174 23604 21180 23656
rect 21232 23644 21238 23656
rect 21232 23616 21277 23644
rect 21232 23604 21238 23616
rect 22002 23604 22008 23656
rect 22060 23644 22066 23656
rect 22281 23647 22339 23653
rect 22281 23644 22293 23647
rect 22060 23616 22293 23644
rect 22060 23604 22066 23616
rect 22281 23613 22293 23616
rect 22327 23613 22339 23647
rect 22462 23644 22468 23656
rect 22423 23616 22468 23644
rect 22281 23607 22339 23613
rect 22462 23604 22468 23616
rect 22520 23604 22526 23656
rect 23109 23647 23167 23653
rect 23109 23613 23121 23647
rect 23155 23613 23167 23647
rect 23109 23607 23167 23613
rect 19794 23576 19800 23588
rect 18831 23548 19472 23576
rect 19755 23548 19800 23576
rect 18831 23545 18843 23548
rect 18785 23539 18843 23545
rect 19794 23536 19800 23548
rect 19852 23536 19858 23588
rect 21100 23576 21128 23604
rect 20916 23548 21128 23576
rect 20916 23520 20944 23548
rect 21358 23536 21364 23588
rect 21416 23576 21422 23588
rect 23124 23576 23152 23607
rect 24854 23604 24860 23656
rect 24912 23644 24918 23656
rect 26237 23647 26295 23653
rect 26237 23644 26249 23647
rect 24912 23616 26249 23644
rect 24912 23604 24918 23616
rect 26237 23613 26249 23616
rect 26283 23613 26295 23647
rect 26344 23644 26372 23684
rect 26421 23681 26433 23715
rect 26467 23712 26479 23715
rect 26694 23712 26700 23724
rect 26467 23684 26700 23712
rect 26467 23681 26479 23684
rect 26421 23675 26479 23681
rect 26694 23672 26700 23684
rect 26752 23672 26758 23724
rect 26970 23712 26976 23724
rect 26931 23684 26976 23712
rect 26970 23672 26976 23684
rect 27028 23672 27034 23724
rect 27154 23712 27160 23724
rect 27080 23684 27160 23712
rect 27080 23644 27108 23684
rect 27154 23672 27160 23684
rect 27212 23672 27218 23724
rect 27430 23672 27436 23724
rect 27488 23712 27494 23724
rect 27525 23715 27583 23721
rect 27525 23712 27537 23715
rect 27488 23684 27537 23712
rect 27488 23672 27494 23684
rect 27525 23681 27537 23684
rect 27571 23681 27583 23715
rect 28166 23712 28172 23724
rect 28127 23684 28172 23712
rect 27525 23675 27583 23681
rect 28166 23672 28172 23684
rect 28224 23672 28230 23724
rect 28276 23718 28304 23752
rect 28332 23721 28390 23727
rect 28460 23721 28488 23820
rect 29454 23808 29460 23860
rect 29512 23848 29518 23860
rect 29733 23851 29791 23857
rect 29733 23848 29745 23851
rect 29512 23820 29745 23848
rect 29512 23808 29518 23820
rect 29733 23817 29745 23820
rect 29779 23817 29791 23851
rect 29733 23811 29791 23817
rect 31294 23808 31300 23860
rect 31352 23848 31358 23860
rect 32309 23851 32367 23857
rect 32309 23848 32321 23851
rect 31352 23820 32321 23848
rect 31352 23808 31358 23820
rect 32309 23817 32321 23820
rect 32355 23817 32367 23851
rect 32309 23811 32367 23817
rect 28718 23740 28724 23792
rect 28776 23780 28782 23792
rect 28776 23752 30696 23780
rect 28776 23740 28782 23752
rect 28332 23718 28344 23721
rect 28276 23690 28344 23718
rect 28332 23687 28344 23690
rect 28378 23687 28390 23721
rect 28332 23681 28390 23687
rect 28432 23715 28490 23721
rect 28432 23681 28444 23715
rect 28478 23681 28490 23715
rect 28432 23675 28490 23681
rect 28534 23672 28540 23724
rect 28592 23712 28598 23724
rect 29270 23712 29276 23724
rect 28592 23684 28637 23712
rect 29231 23684 29276 23712
rect 28592 23672 28598 23684
rect 29270 23672 29276 23684
rect 29328 23672 29334 23724
rect 29362 23672 29368 23724
rect 29420 23712 29426 23724
rect 30668 23721 30696 23752
rect 35268 23752 37780 23780
rect 29736 23715 29794 23721
rect 29736 23712 29748 23715
rect 29420 23684 29748 23712
rect 29420 23672 29426 23684
rect 29736 23681 29748 23684
rect 29782 23681 29794 23715
rect 29736 23675 29794 23681
rect 30653 23715 30711 23721
rect 30653 23681 30665 23715
rect 30699 23681 30711 23715
rect 30653 23675 30711 23681
rect 30745 23715 30803 23721
rect 30745 23681 30757 23715
rect 30791 23712 30803 23715
rect 30791 23684 31248 23712
rect 30791 23681 30803 23684
rect 30745 23675 30803 23681
rect 27246 23644 27252 23656
rect 26344 23616 27108 23644
rect 27207 23616 27252 23644
rect 26237 23607 26295 23613
rect 27246 23604 27252 23616
rect 27304 23604 27310 23656
rect 27338 23604 27344 23656
rect 27396 23644 27402 23656
rect 27709 23647 27767 23653
rect 27396 23616 27441 23644
rect 27396 23604 27402 23616
rect 27709 23613 27721 23647
rect 27755 23644 27767 23647
rect 29178 23644 29184 23656
rect 27755 23616 29184 23644
rect 27755 23613 27767 23616
rect 27709 23607 27767 23613
rect 29178 23604 29184 23616
rect 29236 23604 29242 23656
rect 30558 23644 30564 23656
rect 30519 23616 30564 23644
rect 30558 23604 30564 23616
rect 30616 23604 30622 23656
rect 30837 23647 30895 23653
rect 30837 23613 30849 23647
rect 30883 23644 30895 23647
rect 30926 23644 30932 23656
rect 30883 23616 30932 23644
rect 30883 23613 30895 23616
rect 30837 23607 30895 23613
rect 30926 23604 30932 23616
rect 30984 23604 30990 23656
rect 31220 23644 31248 23684
rect 31478 23672 31484 23724
rect 31536 23712 31542 23724
rect 32125 23715 32183 23721
rect 32125 23712 32137 23715
rect 31536 23684 32137 23712
rect 31536 23672 31542 23684
rect 32125 23681 32137 23684
rect 32171 23681 32183 23715
rect 32125 23675 32183 23681
rect 32214 23672 32220 23724
rect 32272 23712 32278 23724
rect 32272 23684 32317 23712
rect 32272 23672 32278 23684
rect 34698 23672 34704 23724
rect 34756 23712 34762 23724
rect 35268 23721 35296 23752
rect 35253 23715 35311 23721
rect 35253 23712 35265 23715
rect 34756 23684 35265 23712
rect 34756 23672 34762 23684
rect 35253 23681 35265 23684
rect 35299 23681 35311 23715
rect 35253 23675 35311 23681
rect 35342 23672 35348 23724
rect 35400 23712 35406 23724
rect 37752 23721 37780 23752
rect 38010 23721 38016 23724
rect 35509 23715 35567 23721
rect 35509 23712 35521 23715
rect 35400 23684 35521 23712
rect 35400 23672 35406 23684
rect 35509 23681 35521 23684
rect 35555 23681 35567 23715
rect 35509 23675 35567 23681
rect 37737 23715 37795 23721
rect 37737 23681 37749 23715
rect 37783 23681 37795 23715
rect 37737 23675 37795 23681
rect 38004 23675 38016 23721
rect 38068 23712 38074 23724
rect 38068 23684 38104 23712
rect 38010 23672 38016 23675
rect 38068 23672 38074 23684
rect 41874 23672 41880 23724
rect 41932 23712 41938 23724
rect 41932 23684 41977 23712
rect 41932 23672 41938 23684
rect 31754 23644 31760 23656
rect 31220 23616 31760 23644
rect 31754 23604 31760 23616
rect 31812 23644 31818 23656
rect 32232 23644 32260 23672
rect 31812 23616 32260 23644
rect 31812 23604 31818 23616
rect 32306 23604 32312 23656
rect 32364 23644 32370 23656
rect 32585 23647 32643 23653
rect 32585 23644 32597 23647
rect 32364 23616 32597 23644
rect 32364 23604 32370 23616
rect 32585 23613 32597 23616
rect 32631 23613 32643 23647
rect 35360 23644 35388 23672
rect 41322 23644 41328 23656
rect 32585 23607 32643 23613
rect 35268 23616 35388 23644
rect 41283 23616 41328 23644
rect 29546 23576 29552 23588
rect 21416 23548 23152 23576
rect 26252 23548 29552 23576
rect 21416 23536 21422 23548
rect 20898 23468 20904 23520
rect 20956 23468 20962 23520
rect 21821 23511 21879 23517
rect 21821 23477 21833 23511
rect 21867 23508 21879 23511
rect 21910 23508 21916 23520
rect 21867 23480 21916 23508
rect 21867 23477 21879 23480
rect 21821 23471 21879 23477
rect 21910 23468 21916 23480
rect 21968 23468 21974 23520
rect 26252 23517 26280 23548
rect 29546 23536 29552 23548
rect 29604 23536 29610 23588
rect 29638 23536 29644 23588
rect 29696 23576 29702 23588
rect 35268 23576 35296 23616
rect 41322 23604 41328 23616
rect 41380 23604 41386 23656
rect 41690 23644 41696 23656
rect 41651 23616 41696 23644
rect 41690 23604 41696 23616
rect 41748 23604 41754 23656
rect 29696 23548 30512 23576
rect 29696 23536 29702 23548
rect 26237 23511 26295 23517
rect 26237 23477 26249 23511
rect 26283 23477 26295 23511
rect 26237 23471 26295 23477
rect 26329 23511 26387 23517
rect 26329 23477 26341 23511
rect 26375 23508 26387 23511
rect 27338 23508 27344 23520
rect 26375 23480 27344 23508
rect 26375 23477 26387 23480
rect 26329 23471 26387 23477
rect 27338 23468 27344 23480
rect 27396 23468 27402 23520
rect 28813 23511 28871 23517
rect 28813 23477 28825 23511
rect 28859 23508 28871 23511
rect 29365 23511 29423 23517
rect 29365 23508 29377 23511
rect 28859 23480 29377 23508
rect 28859 23477 28871 23480
rect 28813 23471 28871 23477
rect 29365 23477 29377 23480
rect 29411 23477 29423 23511
rect 29365 23471 29423 23477
rect 29917 23511 29975 23517
rect 29917 23477 29929 23511
rect 29963 23508 29975 23511
rect 30098 23508 30104 23520
rect 29963 23480 30104 23508
rect 29963 23477 29975 23480
rect 29917 23471 29975 23477
rect 30098 23468 30104 23480
rect 30156 23468 30162 23520
rect 30374 23508 30380 23520
rect 30335 23480 30380 23508
rect 30374 23468 30380 23480
rect 30432 23468 30438 23520
rect 30484 23508 30512 23548
rect 31726 23548 35296 23576
rect 31726 23508 31754 23548
rect 30484 23480 31754 23508
rect 39022 23468 39028 23520
rect 39080 23508 39086 23520
rect 39117 23511 39175 23517
rect 39117 23508 39129 23511
rect 39080 23480 39129 23508
rect 39080 23468 39086 23480
rect 39117 23477 39129 23480
rect 39163 23477 39175 23511
rect 39117 23471 39175 23477
rect 1104 23418 42872 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 42872 23418
rect 1104 23344 42872 23366
rect 19426 23304 19432 23316
rect 19387 23276 19432 23304
rect 19426 23264 19432 23276
rect 19484 23264 19490 23316
rect 20806 23304 20812 23316
rect 20767 23276 20812 23304
rect 20806 23264 20812 23276
rect 20864 23264 20870 23316
rect 23845 23307 23903 23313
rect 23845 23273 23857 23307
rect 23891 23304 23903 23307
rect 24854 23304 24860 23316
rect 23891 23276 24860 23304
rect 23891 23273 23903 23276
rect 23845 23267 23903 23273
rect 24854 23264 24860 23276
rect 24912 23264 24918 23316
rect 26234 23264 26240 23316
rect 26292 23304 26298 23316
rect 26878 23304 26884 23316
rect 26292 23276 26884 23304
rect 26292 23264 26298 23276
rect 26878 23264 26884 23276
rect 26936 23264 26942 23316
rect 32214 23304 32220 23316
rect 29012 23276 32076 23304
rect 32175 23276 32220 23304
rect 22002 23196 22008 23248
rect 22060 23236 22066 23248
rect 22060 23208 24716 23236
rect 22060 23196 22066 23208
rect 17862 23168 17868 23180
rect 17823 23140 17868 23168
rect 17862 23128 17868 23140
rect 17920 23128 17926 23180
rect 20162 23168 20168 23180
rect 19628 23140 20168 23168
rect 1394 23060 1400 23112
rect 1452 23100 1458 23112
rect 1673 23103 1731 23109
rect 1673 23100 1685 23103
rect 1452 23072 1685 23100
rect 1452 23060 1458 23072
rect 1673 23069 1685 23072
rect 1719 23069 1731 23103
rect 18138 23100 18144 23112
rect 18099 23072 18144 23100
rect 1673 23063 1731 23069
rect 18138 23060 18144 23072
rect 18196 23060 18202 23112
rect 19628 23109 19656 23140
rect 20162 23128 20168 23140
rect 20220 23128 20226 23180
rect 22020 23168 22048 23196
rect 23382 23168 23388 23180
rect 21100 23140 22048 23168
rect 23343 23140 23388 23168
rect 19613 23103 19671 23109
rect 19613 23069 19625 23103
rect 19659 23069 19671 23103
rect 19794 23100 19800 23112
rect 19755 23072 19800 23100
rect 19613 23063 19671 23069
rect 19794 23060 19800 23072
rect 19852 23060 19858 23112
rect 19981 23103 20039 23109
rect 19981 23069 19993 23103
rect 20027 23100 20039 23103
rect 20714 23100 20720 23112
rect 20027 23072 20720 23100
rect 20027 23069 20039 23072
rect 19981 23063 20039 23069
rect 20714 23060 20720 23072
rect 20772 23060 20778 23112
rect 21100 23109 21128 23140
rect 23382 23128 23388 23140
rect 23440 23128 23446 23180
rect 24394 23168 24400 23180
rect 24355 23140 24400 23168
rect 24394 23128 24400 23140
rect 24452 23128 24458 23180
rect 24688 23177 24716 23208
rect 26326 23196 26332 23248
rect 26384 23236 26390 23248
rect 29012 23236 29040 23276
rect 32048 23236 32076 23276
rect 32214 23264 32220 23276
rect 32272 23264 32278 23316
rect 38654 23304 38660 23316
rect 38615 23276 38660 23304
rect 38654 23264 38660 23276
rect 38712 23264 38718 23316
rect 32398 23236 32404 23248
rect 26384 23208 29040 23236
rect 29288 23208 29776 23236
rect 32048 23208 32404 23236
rect 26384 23196 26390 23208
rect 24673 23171 24731 23177
rect 24673 23137 24685 23171
rect 24719 23137 24731 23171
rect 24673 23131 24731 23137
rect 28810 23128 28816 23180
rect 28868 23168 28874 23180
rect 29288 23168 29316 23208
rect 29546 23168 29552 23180
rect 28868 23140 29316 23168
rect 29507 23140 29552 23168
rect 28868 23128 28874 23140
rect 29546 23128 29552 23140
rect 29604 23128 29610 23180
rect 20809 23103 20867 23109
rect 20809 23069 20821 23103
rect 20855 23100 20867 23103
rect 21085 23103 21143 23109
rect 20855 23072 21036 23100
rect 20855 23069 20867 23072
rect 20809 23063 20867 23069
rect 19705 23035 19763 23041
rect 19705 23001 19717 23035
rect 19751 23032 19763 23035
rect 20622 23032 20628 23044
rect 19751 23004 20628 23032
rect 19751 23001 19763 23004
rect 19705 22995 19763 23001
rect 20622 22992 20628 23004
rect 20680 22992 20686 23044
rect 20898 23032 20904 23044
rect 20859 23004 20904 23032
rect 20898 22992 20904 23004
rect 20956 22992 20962 23044
rect 21008 23032 21036 23072
rect 21085 23069 21097 23103
rect 21131 23069 21143 23103
rect 22465 23103 22523 23109
rect 22465 23100 22477 23103
rect 21085 23063 21143 23069
rect 22066 23072 22477 23100
rect 21174 23032 21180 23044
rect 21008 23004 21180 23032
rect 21174 22992 21180 23004
rect 21232 23032 21238 23044
rect 22066 23032 22094 23072
rect 22465 23069 22477 23072
rect 22511 23069 22523 23103
rect 23290 23100 23296 23112
rect 23251 23072 23296 23100
rect 22465 23063 22523 23069
rect 23290 23060 23296 23072
rect 23348 23060 23354 23112
rect 23569 23103 23627 23109
rect 23569 23069 23581 23103
rect 23615 23069 23627 23103
rect 23569 23063 23627 23069
rect 23661 23103 23719 23109
rect 23661 23069 23673 23103
rect 23707 23100 23719 23103
rect 23842 23100 23848 23112
rect 23707 23072 23848 23100
rect 23707 23069 23719 23072
rect 23661 23063 23719 23069
rect 21232 23004 22094 23032
rect 22557 23035 22615 23041
rect 21232 22992 21238 23004
rect 22557 23001 22569 23035
rect 22603 23032 22615 23035
rect 23584 23032 23612 23063
rect 23842 23060 23848 23072
rect 23900 23100 23906 23112
rect 24486 23100 24492 23112
rect 23900 23072 24492 23100
rect 23900 23060 23906 23072
rect 24486 23060 24492 23072
rect 24544 23060 24550 23112
rect 29748 23109 29776 23208
rect 32398 23196 32404 23208
rect 32456 23196 32462 23248
rect 38197 23239 38255 23245
rect 38197 23205 38209 23239
rect 38243 23236 38255 23239
rect 38243 23208 39068 23236
rect 38243 23205 38255 23208
rect 38197 23199 38255 23205
rect 30101 23171 30159 23177
rect 30101 23137 30113 23171
rect 30147 23168 30159 23171
rect 30374 23168 30380 23180
rect 30147 23140 30380 23168
rect 30147 23137 30159 23140
rect 30101 23131 30159 23137
rect 30374 23128 30380 23140
rect 30432 23128 30438 23180
rect 30834 23168 30840 23180
rect 30795 23140 30840 23168
rect 30834 23128 30840 23140
rect 30892 23128 30898 23180
rect 34698 23128 34704 23180
rect 34756 23168 34762 23180
rect 39040 23177 39068 23208
rect 39390 23196 39396 23248
rect 39448 23236 39454 23248
rect 39448 23208 40816 23236
rect 39448 23196 39454 23208
rect 34885 23171 34943 23177
rect 34885 23168 34897 23171
rect 34756 23140 34897 23168
rect 34756 23128 34762 23140
rect 34885 23137 34897 23140
rect 34931 23137 34943 23171
rect 34885 23131 34943 23137
rect 39025 23171 39083 23177
rect 39025 23137 39037 23171
rect 39071 23137 39083 23171
rect 40494 23168 40500 23180
rect 40455 23140 40500 23168
rect 39025 23131 39083 23137
rect 31110 23109 31116 23112
rect 28169 23103 28227 23109
rect 28169 23069 28181 23103
rect 28215 23100 28227 23103
rect 29733 23103 29791 23109
rect 28215 23072 29500 23100
rect 28215 23069 28227 23072
rect 28169 23063 28227 23069
rect 22603 23004 23612 23032
rect 22603 23001 22615 23004
rect 22557 22995 22615 23001
rect 24210 22992 24216 23044
rect 24268 23032 24274 23044
rect 24394 23032 24400 23044
rect 24268 23004 24400 23032
rect 24268 22992 24274 23004
rect 24394 22992 24400 23004
rect 24452 22992 24458 23044
rect 26970 22992 26976 23044
rect 27028 23032 27034 23044
rect 28721 23035 28779 23041
rect 28721 23032 28733 23035
rect 27028 23004 28733 23032
rect 27028 22992 27034 23004
rect 28721 23001 28733 23004
rect 28767 23001 28779 23035
rect 29472 23032 29500 23072
rect 29733 23069 29745 23103
rect 29779 23069 29791 23103
rect 31104 23100 31116 23109
rect 31071 23072 31116 23100
rect 29733 23063 29791 23069
rect 31104 23063 31116 23072
rect 31110 23060 31116 23063
rect 31168 23060 31174 23112
rect 34900 23100 34928 23131
rect 40494 23128 40500 23140
rect 40552 23128 40558 23180
rect 40788 23177 40816 23208
rect 40773 23171 40831 23177
rect 40773 23137 40785 23171
rect 40819 23137 40831 23171
rect 40773 23131 40831 23137
rect 36817 23103 36875 23109
rect 36817 23100 36829 23103
rect 34900 23072 36829 23100
rect 36817 23069 36829 23072
rect 36863 23069 36875 23103
rect 36817 23063 36875 23069
rect 38841 23103 38899 23109
rect 38841 23069 38853 23103
rect 38887 23100 38899 23103
rect 38930 23100 38936 23112
rect 38887 23072 38936 23100
rect 38887 23069 38899 23072
rect 38841 23063 38899 23069
rect 38930 23060 38936 23072
rect 38988 23100 38994 23112
rect 39942 23100 39948 23112
rect 38988 23072 39948 23100
rect 38988 23060 38994 23072
rect 39942 23060 39948 23072
rect 40000 23060 40006 23112
rect 40310 23100 40316 23112
rect 40271 23072 40316 23100
rect 40310 23060 40316 23072
rect 40368 23060 40374 23112
rect 30009 23035 30067 23041
rect 29472 23004 29960 23032
rect 28721 22995 28779 23001
rect 28810 22964 28816 22976
rect 28771 22936 28816 22964
rect 28810 22924 28816 22936
rect 28868 22924 28874 22976
rect 29932 22964 29960 23004
rect 30009 23001 30021 23035
rect 30055 23032 30067 23035
rect 30466 23032 30472 23044
rect 30055 23004 30472 23032
rect 30055 23001 30067 23004
rect 30009 22995 30067 23001
rect 30466 22992 30472 23004
rect 30524 22992 30530 23044
rect 34882 22992 34888 23044
rect 34940 23032 34946 23044
rect 37090 23041 37096 23044
rect 35130 23035 35188 23041
rect 35130 23032 35142 23035
rect 34940 23004 35142 23032
rect 34940 22992 34946 23004
rect 35130 23001 35142 23004
rect 35176 23001 35188 23035
rect 35130 22995 35188 23001
rect 37084 22995 37096 23041
rect 37148 23032 37154 23044
rect 37148 23004 37184 23032
rect 37090 22992 37096 22995
rect 37148 22992 37154 23004
rect 39574 22964 39580 22976
rect 29932 22936 39580 22964
rect 39574 22924 39580 22936
rect 39632 22924 39638 22976
rect 1104 22874 42872 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 42872 22874
rect 1104 22800 42872 22822
rect 17678 22720 17684 22772
rect 17736 22760 17742 22772
rect 17865 22763 17923 22769
rect 17865 22760 17877 22763
rect 17736 22732 17877 22760
rect 17736 22720 17742 22732
rect 17865 22729 17877 22732
rect 17911 22729 17923 22763
rect 17865 22723 17923 22729
rect 20622 22720 20628 22772
rect 20680 22760 20686 22772
rect 25961 22763 26019 22769
rect 20680 22732 25544 22760
rect 20680 22720 20686 22732
rect 21450 22652 21456 22704
rect 21508 22692 21514 22704
rect 21508 22664 23520 22692
rect 21508 22652 21514 22664
rect 2130 22624 2136 22636
rect 2043 22596 2136 22624
rect 2130 22584 2136 22596
rect 2188 22624 2194 22636
rect 9214 22624 9220 22636
rect 2188 22596 9220 22624
rect 2188 22584 2194 22596
rect 9214 22584 9220 22596
rect 9272 22584 9278 22636
rect 18046 22624 18052 22636
rect 18007 22596 18052 22624
rect 18046 22584 18052 22596
rect 18104 22584 18110 22636
rect 18598 22624 18604 22636
rect 18559 22596 18604 22624
rect 18598 22584 18604 22596
rect 18656 22584 18662 22636
rect 20898 22584 20904 22636
rect 20956 22624 20962 22636
rect 23492 22633 23520 22664
rect 22649 22627 22707 22633
rect 22649 22624 22661 22627
rect 20956 22596 22661 22624
rect 20956 22584 20962 22596
rect 22649 22593 22661 22596
rect 22695 22593 22707 22627
rect 22649 22587 22707 22593
rect 23477 22627 23535 22633
rect 23477 22593 23489 22627
rect 23523 22593 23535 22627
rect 23477 22587 23535 22593
rect 23753 22627 23811 22633
rect 23753 22593 23765 22627
rect 23799 22593 23811 22627
rect 23753 22587 23811 22593
rect 22738 22516 22744 22568
rect 22796 22556 22802 22568
rect 22925 22559 22983 22565
rect 22925 22556 22937 22559
rect 22796 22528 22937 22556
rect 22796 22516 22802 22528
rect 22925 22525 22937 22528
rect 22971 22556 22983 22559
rect 23768 22556 23796 22587
rect 23842 22584 23848 22636
rect 23900 22624 23906 22636
rect 25516 22633 25544 22732
rect 25961 22729 25973 22763
rect 26007 22760 26019 22763
rect 27246 22760 27252 22772
rect 26007 22732 27252 22760
rect 26007 22729 26019 22732
rect 25961 22723 26019 22729
rect 27246 22720 27252 22732
rect 27304 22720 27310 22772
rect 38289 22763 38347 22769
rect 38289 22729 38301 22763
rect 38335 22760 38347 22763
rect 40310 22760 40316 22772
rect 38335 22732 40316 22760
rect 38335 22729 38347 22732
rect 38289 22723 38347 22729
rect 40310 22720 40316 22732
rect 40368 22720 40374 22772
rect 26326 22692 26332 22704
rect 25608 22664 26332 22692
rect 25608 22633 25636 22664
rect 26326 22652 26332 22664
rect 26384 22692 26390 22704
rect 28169 22695 28227 22701
rect 28169 22692 28181 22695
rect 26384 22664 28181 22692
rect 26384 22652 26390 22664
rect 28169 22661 28181 22664
rect 28215 22661 28227 22695
rect 28169 22655 28227 22661
rect 34698 22652 34704 22704
rect 34756 22692 34762 22704
rect 34756 22664 38792 22692
rect 34756 22652 34762 22664
rect 25501 22627 25559 22633
rect 23900 22596 23945 22624
rect 23900 22584 23906 22596
rect 25501 22593 25513 22627
rect 25547 22593 25559 22627
rect 25501 22587 25559 22593
rect 25593 22627 25651 22633
rect 25593 22593 25605 22627
rect 25639 22593 25651 22627
rect 25593 22587 25651 22593
rect 25777 22627 25835 22633
rect 25777 22593 25789 22627
rect 25823 22593 25835 22627
rect 26970 22624 26976 22636
rect 26931 22596 26976 22624
rect 25777 22587 25835 22593
rect 22971 22528 23796 22556
rect 22971 22525 22983 22528
rect 22925 22519 22983 22525
rect 25130 22516 25136 22568
rect 25188 22556 25194 22568
rect 25792 22556 25820 22587
rect 26970 22584 26976 22596
rect 27028 22584 27034 22636
rect 27154 22624 27160 22636
rect 27115 22596 27160 22624
rect 27154 22584 27160 22596
rect 27212 22584 27218 22636
rect 27522 22584 27528 22636
rect 27580 22624 27586 22636
rect 28350 22624 28356 22636
rect 27580 22596 27625 22624
rect 28311 22596 28356 22624
rect 27580 22584 27586 22596
rect 28350 22584 28356 22596
rect 28408 22584 28414 22636
rect 28442 22584 28448 22636
rect 28500 22624 28506 22636
rect 29086 22624 29092 22636
rect 28500 22596 28545 22624
rect 29047 22596 29092 22624
rect 28500 22584 28506 22596
rect 29086 22584 29092 22596
rect 29144 22584 29150 22636
rect 29178 22584 29184 22636
rect 29236 22624 29242 22636
rect 29457 22627 29515 22633
rect 29236 22596 29281 22624
rect 29236 22584 29242 22596
rect 29457 22593 29469 22627
rect 29503 22624 29515 22627
rect 29822 22624 29828 22636
rect 29503 22596 29828 22624
rect 29503 22593 29515 22596
rect 29457 22587 29515 22593
rect 29822 22584 29828 22596
rect 29880 22584 29886 22636
rect 30101 22627 30159 22633
rect 30101 22593 30113 22627
rect 30147 22593 30159 22627
rect 30101 22587 30159 22593
rect 30285 22627 30343 22633
rect 30285 22593 30297 22627
rect 30331 22624 30343 22627
rect 31386 22624 31392 22636
rect 30331 22596 31392 22624
rect 30331 22593 30343 22596
rect 30285 22587 30343 22593
rect 25188 22528 25820 22556
rect 27249 22559 27307 22565
rect 25188 22516 25194 22528
rect 27249 22525 27261 22559
rect 27295 22525 27307 22559
rect 27249 22519 27307 22525
rect 23382 22448 23388 22500
rect 23440 22488 23446 22500
rect 23569 22491 23627 22497
rect 23569 22488 23581 22491
rect 23440 22460 23581 22488
rect 23440 22448 23446 22460
rect 23569 22457 23581 22460
rect 23615 22457 23627 22491
rect 23569 22451 23627 22457
rect 24029 22491 24087 22497
rect 24029 22457 24041 22491
rect 24075 22488 24087 22491
rect 27264 22488 27292 22519
rect 27338 22516 27344 22568
rect 27396 22556 27402 22568
rect 27396 22528 27441 22556
rect 27396 22516 27402 22528
rect 29546 22516 29552 22568
rect 29604 22556 29610 22568
rect 30116 22556 30144 22587
rect 31386 22584 31392 22596
rect 31444 22584 31450 22636
rect 32122 22624 32128 22636
rect 32083 22596 32128 22624
rect 32122 22584 32128 22596
rect 32180 22584 32186 22636
rect 32214 22584 32220 22636
rect 32272 22624 32278 22636
rect 32309 22627 32367 22633
rect 32309 22624 32321 22627
rect 32272 22596 32321 22624
rect 32272 22584 32278 22596
rect 32309 22593 32321 22596
rect 32355 22593 32367 22627
rect 32309 22587 32367 22593
rect 32398 22584 32404 22636
rect 32456 22624 32462 22636
rect 32456 22596 32501 22624
rect 32456 22584 32462 22596
rect 34514 22584 34520 22636
rect 34572 22624 34578 22636
rect 35176 22633 35204 22664
rect 38764 22633 38792 22664
rect 34894 22627 34952 22633
rect 34894 22624 34906 22627
rect 34572 22596 34906 22624
rect 34572 22584 34578 22596
rect 34894 22593 34906 22596
rect 34940 22593 34952 22627
rect 34894 22587 34952 22593
rect 35161 22627 35219 22633
rect 35161 22593 35173 22627
rect 35207 22593 35219 22627
rect 35161 22587 35219 22593
rect 38105 22627 38163 22633
rect 38105 22593 38117 22627
rect 38151 22624 38163 22627
rect 38749 22627 38807 22633
rect 38151 22596 38700 22624
rect 38151 22593 38163 22596
rect 38105 22587 38163 22593
rect 29604 22528 30144 22556
rect 29604 22516 29610 22528
rect 24075 22460 27292 22488
rect 27709 22491 27767 22497
rect 24075 22457 24087 22460
rect 24029 22451 24087 22457
rect 27709 22457 27721 22491
rect 27755 22488 27767 22491
rect 29730 22488 29736 22500
rect 27755 22460 29736 22488
rect 27755 22457 27767 22460
rect 27709 22451 27767 22457
rect 29730 22448 29736 22460
rect 29788 22448 29794 22500
rect 1578 22380 1584 22432
rect 1636 22420 1642 22432
rect 2041 22423 2099 22429
rect 2041 22420 2053 22423
rect 1636 22392 2053 22420
rect 1636 22380 1642 22392
rect 2041 22389 2053 22392
rect 2087 22389 2099 22423
rect 2041 22383 2099 22389
rect 18785 22423 18843 22429
rect 18785 22389 18797 22423
rect 18831 22420 18843 22423
rect 19058 22420 19064 22432
rect 18831 22392 19064 22420
rect 18831 22389 18843 22392
rect 18785 22383 18843 22389
rect 19058 22380 19064 22392
rect 19116 22380 19122 22432
rect 27154 22380 27160 22432
rect 27212 22420 27218 22432
rect 28169 22423 28227 22429
rect 28169 22420 28181 22423
rect 27212 22392 28181 22420
rect 27212 22380 27218 22392
rect 28169 22389 28181 22392
rect 28215 22389 28227 22423
rect 28169 22383 28227 22389
rect 28718 22380 28724 22432
rect 28776 22420 28782 22432
rect 28905 22423 28963 22429
rect 28905 22420 28917 22423
rect 28776 22392 28917 22420
rect 28776 22380 28782 22392
rect 28905 22389 28917 22392
rect 28951 22389 28963 22423
rect 28905 22383 28963 22389
rect 29365 22423 29423 22429
rect 29365 22389 29377 22423
rect 29411 22420 29423 22423
rect 29917 22423 29975 22429
rect 29917 22420 29929 22423
rect 29411 22392 29929 22420
rect 29411 22389 29423 22392
rect 29365 22383 29423 22389
rect 29917 22389 29929 22392
rect 29963 22389 29975 22423
rect 29917 22383 29975 22389
rect 32125 22423 32183 22429
rect 32125 22389 32137 22423
rect 32171 22420 32183 22423
rect 32858 22420 32864 22432
rect 32171 22392 32864 22420
rect 32171 22389 32183 22392
rect 32125 22383 32183 22389
rect 32858 22380 32864 22392
rect 32916 22380 32922 22432
rect 38672 22420 38700 22596
rect 38749 22593 38761 22627
rect 38795 22593 38807 22627
rect 38749 22587 38807 22593
rect 38838 22584 38844 22636
rect 38896 22624 38902 22636
rect 39005 22627 39063 22633
rect 39005 22624 39017 22627
rect 38896 22596 39017 22624
rect 38896 22584 38902 22596
rect 39005 22593 39017 22596
rect 39051 22593 39063 22627
rect 39005 22587 39063 22593
rect 39942 22584 39948 22636
rect 40000 22624 40006 22636
rect 40773 22627 40831 22633
rect 40773 22624 40785 22627
rect 40000 22596 40785 22624
rect 40000 22584 40006 22596
rect 40773 22593 40785 22596
rect 40819 22593 40831 22627
rect 40773 22587 40831 22593
rect 41417 22627 41475 22633
rect 41417 22593 41429 22627
rect 41463 22624 41475 22627
rect 41966 22624 41972 22636
rect 41463 22596 41972 22624
rect 41463 22593 41475 22596
rect 41417 22587 41475 22593
rect 41966 22584 41972 22596
rect 42024 22584 42030 22636
rect 40957 22559 41015 22565
rect 40957 22525 40969 22559
rect 41003 22525 41015 22559
rect 40957 22519 41015 22525
rect 40129 22491 40187 22497
rect 40129 22457 40141 22491
rect 40175 22488 40187 22491
rect 40972 22488 41000 22519
rect 40175 22460 41000 22488
rect 40175 22457 40187 22460
rect 40129 22451 40187 22457
rect 40589 22423 40647 22429
rect 40589 22420 40601 22423
rect 38672 22392 40601 22420
rect 40589 22389 40601 22392
rect 40635 22389 40647 22423
rect 40589 22383 40647 22389
rect 40678 22380 40684 22432
rect 40736 22420 40742 22432
rect 41509 22423 41567 22429
rect 41509 22420 41521 22423
rect 40736 22392 41521 22420
rect 40736 22380 40742 22392
rect 41509 22389 41521 22392
rect 41555 22389 41567 22423
rect 41509 22383 41567 22389
rect 1104 22330 42872 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 42872 22330
rect 1104 22256 42872 22278
rect 18233 22219 18291 22225
rect 18233 22185 18245 22219
rect 18279 22216 18291 22219
rect 18598 22216 18604 22228
rect 18279 22188 18604 22216
rect 18279 22185 18291 22188
rect 18233 22179 18291 22185
rect 18598 22176 18604 22188
rect 18656 22176 18662 22228
rect 20809 22219 20867 22225
rect 20809 22185 20821 22219
rect 20855 22216 20867 22219
rect 21726 22216 21732 22228
rect 20855 22188 21732 22216
rect 20855 22185 20867 22188
rect 20809 22179 20867 22185
rect 21726 22176 21732 22188
rect 21784 22176 21790 22228
rect 22738 22216 22744 22228
rect 22699 22188 22744 22216
rect 22738 22176 22744 22188
rect 22796 22176 22802 22228
rect 24486 22216 24492 22228
rect 24447 22188 24492 22216
rect 24486 22176 24492 22188
rect 24544 22176 24550 22228
rect 26697 22219 26755 22225
rect 26697 22185 26709 22219
rect 26743 22216 26755 22219
rect 26970 22216 26976 22228
rect 26743 22188 26976 22216
rect 26743 22185 26755 22188
rect 26697 22179 26755 22185
rect 26970 22176 26976 22188
rect 27028 22176 27034 22228
rect 29638 22176 29644 22228
rect 29696 22216 29702 22228
rect 29733 22219 29791 22225
rect 29733 22216 29745 22219
rect 29696 22188 29745 22216
rect 29696 22176 29702 22188
rect 29733 22185 29745 22188
rect 29779 22185 29791 22219
rect 29733 22179 29791 22185
rect 29822 22176 29828 22228
rect 29880 22216 29886 22228
rect 31941 22219 31999 22225
rect 29880 22188 29925 22216
rect 29880 22176 29886 22188
rect 31941 22185 31953 22219
rect 31987 22216 31999 22219
rect 32122 22216 32128 22228
rect 31987 22188 32128 22216
rect 31987 22185 31999 22188
rect 31941 22179 31999 22185
rect 32122 22176 32128 22188
rect 32180 22176 32186 22228
rect 16224 22120 16528 22148
rect 16224 22092 16252 22120
rect 1394 22080 1400 22092
rect 1355 22052 1400 22080
rect 1394 22040 1400 22052
rect 1452 22040 1458 22092
rect 1578 22080 1584 22092
rect 1539 22052 1584 22080
rect 1578 22040 1584 22052
rect 1636 22040 1642 22092
rect 1854 22080 1860 22092
rect 1815 22052 1860 22080
rect 1854 22040 1860 22052
rect 1912 22040 1918 22092
rect 15654 22040 15660 22092
rect 15712 22080 15718 22092
rect 15933 22083 15991 22089
rect 15933 22080 15945 22083
rect 15712 22052 15945 22080
rect 15712 22040 15718 22052
rect 15933 22049 15945 22052
rect 15979 22049 15991 22083
rect 16206 22080 16212 22092
rect 16119 22052 16212 22080
rect 15933 22043 15991 22049
rect 16206 22040 16212 22052
rect 16264 22040 16270 22092
rect 16500 22080 16528 22120
rect 17862 22108 17868 22160
rect 17920 22148 17926 22160
rect 20714 22148 20720 22160
rect 17920 22120 19748 22148
rect 20675 22120 20720 22148
rect 17920 22108 17926 22120
rect 19720 22080 19748 22120
rect 20714 22108 20720 22120
rect 20772 22108 20778 22160
rect 23382 22108 23388 22160
rect 23440 22148 23446 22160
rect 25130 22148 25136 22160
rect 23440 22120 25136 22148
rect 23440 22108 23446 22120
rect 20625 22083 20683 22089
rect 16500 22052 18000 22080
rect 19720 22052 19840 22080
rect 17972 22024 18000 22052
rect 12894 21972 12900 22024
rect 12952 22012 12958 22024
rect 14366 22012 14372 22024
rect 12952 21984 14372 22012
rect 12952 21972 12958 21984
rect 14366 21972 14372 21984
rect 14424 22012 14430 22024
rect 15470 22012 15476 22024
rect 14424 21984 15476 22012
rect 14424 21972 14430 21984
rect 15470 21972 15476 21984
rect 15528 21972 15534 22024
rect 15838 21972 15844 22024
rect 15896 22012 15902 22024
rect 16301 22015 16359 22021
rect 16301 22012 16313 22015
rect 15896 21984 16313 22012
rect 15896 21972 15902 21984
rect 16301 21981 16313 21984
rect 16347 21981 16359 22015
rect 17954 22012 17960 22024
rect 17915 21984 17960 22012
rect 16301 21975 16359 21981
rect 17954 21972 17960 21984
rect 18012 21972 18018 22024
rect 18049 22015 18107 22021
rect 18049 21981 18061 22015
rect 18095 22012 18107 22015
rect 18138 22012 18144 22024
rect 18095 21984 18144 22012
rect 18095 21981 18107 21984
rect 18049 21975 18107 21981
rect 18138 21972 18144 21984
rect 18196 21972 18202 22024
rect 19812 22021 19840 22052
rect 20625 22049 20637 22083
rect 20671 22049 20683 22083
rect 20625 22043 20683 22049
rect 19797 22015 19855 22021
rect 19797 21981 19809 22015
rect 19843 21981 19855 22015
rect 19797 21975 19855 21981
rect 15228 21947 15286 21953
rect 15228 21913 15240 21947
rect 15274 21944 15286 21947
rect 15378 21944 15384 21956
rect 15274 21916 15384 21944
rect 15274 21913 15286 21916
rect 15228 21907 15286 21913
rect 15378 21904 15384 21916
rect 15436 21904 15442 21956
rect 20640 21888 20668 22043
rect 20898 22012 20904 22024
rect 20859 21984 20904 22012
rect 20898 21972 20904 21984
rect 20956 21972 20962 22024
rect 21358 22012 21364 22024
rect 21271 21984 21364 22012
rect 21358 21972 21364 21984
rect 21416 22012 21422 22024
rect 22002 22012 22008 22024
rect 21416 21984 22008 22012
rect 21416 21972 21422 21984
rect 22002 21972 22008 21984
rect 22060 21972 22066 22024
rect 24210 21972 24216 22024
rect 24268 22012 24274 22024
rect 24596 22021 24624 22120
rect 25130 22108 25136 22120
rect 25188 22148 25194 22160
rect 25593 22151 25651 22157
rect 25593 22148 25605 22151
rect 25188 22120 25605 22148
rect 25188 22108 25194 22120
rect 25593 22117 25605 22120
rect 25639 22117 25651 22151
rect 28350 22148 28356 22160
rect 25593 22111 25651 22117
rect 27632 22120 28356 22148
rect 24397 22015 24455 22021
rect 24397 22012 24409 22015
rect 24268 21984 24409 22012
rect 24268 21972 24274 21984
rect 24397 21981 24409 21984
rect 24443 21981 24455 22015
rect 24397 21975 24455 21981
rect 24581 22015 24639 22021
rect 24581 21981 24593 22015
rect 24627 21981 24639 22015
rect 24581 21975 24639 21981
rect 25777 22015 25835 22021
rect 25777 21981 25789 22015
rect 25823 22012 25835 22015
rect 26050 22012 26056 22024
rect 25823 21984 26056 22012
rect 25823 21981 25835 21984
rect 25777 21975 25835 21981
rect 26050 21972 26056 21984
rect 26108 22012 26114 22024
rect 27065 22015 27123 22021
rect 26108 21984 27016 22012
rect 26108 21972 26114 21984
rect 21628 21947 21686 21953
rect 21628 21913 21640 21947
rect 21674 21944 21686 21947
rect 21818 21944 21824 21956
rect 21674 21916 21824 21944
rect 21674 21913 21686 21916
rect 21628 21907 21686 21913
rect 21818 21904 21824 21916
rect 21876 21904 21882 21956
rect 25958 21944 25964 21956
rect 25919 21916 25964 21944
rect 25958 21904 25964 21916
rect 26016 21944 26022 21956
rect 26881 21947 26939 21953
rect 26881 21944 26893 21947
rect 26016 21916 26893 21944
rect 26016 21904 26022 21916
rect 26881 21913 26893 21916
rect 26927 21913 26939 21947
rect 26988 21944 27016 21984
rect 27065 21981 27077 22015
rect 27111 22012 27123 22015
rect 27632 22012 27660 22120
rect 28350 22108 28356 22120
rect 28408 22108 28414 22160
rect 28721 22151 28779 22157
rect 28721 22117 28733 22151
rect 28767 22117 28779 22151
rect 28721 22111 28779 22117
rect 27798 22080 27804 22092
rect 27759 22052 27804 22080
rect 27798 22040 27804 22052
rect 27856 22040 27862 22092
rect 28166 22040 28172 22092
rect 28224 22080 28230 22092
rect 28736 22080 28764 22111
rect 28948 22108 28954 22160
rect 29006 22148 29012 22160
rect 29546 22148 29552 22160
rect 29006 22120 29552 22148
rect 29006 22108 29012 22120
rect 29546 22108 29552 22120
rect 29604 22108 29610 22160
rect 29730 22080 29736 22092
rect 28224 22052 28764 22080
rect 29691 22052 29736 22080
rect 28224 22040 28230 22052
rect 29730 22040 29736 22052
rect 29788 22040 29794 22092
rect 29840 22080 29868 22176
rect 32033 22151 32091 22157
rect 32033 22117 32045 22151
rect 32079 22148 32091 22151
rect 32398 22148 32404 22160
rect 32079 22120 32404 22148
rect 32079 22117 32091 22120
rect 32033 22111 32091 22117
rect 32398 22108 32404 22120
rect 32456 22108 32462 22160
rect 30469 22083 30527 22089
rect 30469 22080 30481 22083
rect 29840 22052 30481 22080
rect 30469 22049 30481 22052
rect 30515 22049 30527 22083
rect 31849 22083 31907 22089
rect 31849 22080 31861 22083
rect 30469 22043 30527 22049
rect 31726 22052 31861 22080
rect 27111 21984 27660 22012
rect 27111 21981 27123 21984
rect 27065 21975 27123 21981
rect 28442 21972 28448 22024
rect 28500 22012 28506 22024
rect 28618 22015 28676 22021
rect 28618 22012 28630 22015
rect 28500 21984 28630 22012
rect 28500 21972 28506 21984
rect 28618 21981 28630 21984
rect 28664 21981 28676 22015
rect 28905 22015 28963 22021
rect 28905 22002 28917 22015
rect 28951 22002 28963 22015
rect 28618 21975 28676 21981
rect 27617 21947 27675 21953
rect 28902 21950 28908 22002
rect 28960 21950 28966 22002
rect 28994 21972 29000 22024
rect 29052 22012 29058 22024
rect 29917 22015 29975 22021
rect 29052 21984 29868 22012
rect 29052 21972 29058 21984
rect 27617 21944 27629 21947
rect 26988 21916 27629 21944
rect 26881 21907 26939 21913
rect 27617 21913 27629 21916
rect 27663 21913 27675 21947
rect 27617 21907 27675 21913
rect 29549 21947 29607 21953
rect 29549 21913 29561 21947
rect 29595 21944 29607 21947
rect 29730 21944 29736 21956
rect 29595 21916 29736 21944
rect 29595 21913 29607 21916
rect 29549 21907 29607 21913
rect 14093 21879 14151 21885
rect 14093 21845 14105 21879
rect 14139 21876 14151 21879
rect 15102 21876 15108 21888
rect 14139 21848 15108 21876
rect 14139 21845 14151 21848
rect 14093 21839 14151 21845
rect 15102 21836 15108 21848
rect 15160 21836 15166 21888
rect 19705 21879 19763 21885
rect 19705 21845 19717 21879
rect 19751 21876 19763 21879
rect 19978 21876 19984 21888
rect 19751 21848 19984 21876
rect 19751 21845 19763 21848
rect 19705 21839 19763 21845
rect 19978 21836 19984 21848
rect 20036 21836 20042 21888
rect 20622 21876 20628 21888
rect 20535 21848 20628 21876
rect 20622 21836 20628 21848
rect 20680 21876 20686 21888
rect 22922 21876 22928 21888
rect 20680 21848 22928 21876
rect 20680 21836 20686 21848
rect 22922 21836 22928 21848
rect 22980 21836 22986 21888
rect 26896 21876 26924 21907
rect 29730 21904 29736 21916
rect 29788 21904 29794 21956
rect 29840 21944 29868 21984
rect 29917 21981 29929 22015
rect 29963 22012 29975 22015
rect 30190 22012 30196 22024
rect 29963 21984 30196 22012
rect 29963 21981 29975 21984
rect 29917 21975 29975 21981
rect 30190 21972 30196 21984
rect 30248 21972 30254 22024
rect 30282 21972 30288 22024
rect 30340 22014 30346 22024
rect 30377 22015 30435 22021
rect 30377 22014 30389 22015
rect 30340 21986 30389 22014
rect 30340 21972 30346 21986
rect 30377 21981 30389 21986
rect 30423 21981 30435 22015
rect 30377 21975 30435 21981
rect 31726 21944 31754 22052
rect 31849 22049 31861 22052
rect 31895 22049 31907 22083
rect 31849 22043 31907 22049
rect 34701 22083 34759 22089
rect 34701 22049 34713 22083
rect 34747 22080 34759 22083
rect 34747 22052 35572 22080
rect 34747 22049 34759 22052
rect 34701 22043 34759 22049
rect 32125 22015 32183 22021
rect 32125 21981 32137 22015
rect 32171 22012 32183 22015
rect 32214 22012 32220 22024
rect 32171 21984 32220 22012
rect 32171 21981 32183 21984
rect 32125 21975 32183 21981
rect 32214 21972 32220 21984
rect 32272 21972 32278 22024
rect 32306 21972 32312 22024
rect 32364 22012 32370 22024
rect 32769 22015 32827 22021
rect 32769 22012 32781 22015
rect 32364 21984 32781 22012
rect 32364 21972 32370 21984
rect 32769 21981 32781 21984
rect 32815 21981 32827 22015
rect 32769 21975 32827 21981
rect 32858 21972 32864 22024
rect 32916 22012 32922 22024
rect 33025 22015 33083 22021
rect 33025 22012 33037 22015
rect 32916 21984 33037 22012
rect 32916 21972 32922 21984
rect 33025 21981 33037 21984
rect 33071 21981 33083 22015
rect 33025 21975 33083 21981
rect 29840 21916 31754 21944
rect 28166 21876 28172 21888
rect 26896 21848 28172 21876
rect 28166 21836 28172 21848
rect 28224 21836 28230 21888
rect 28629 21879 28687 21885
rect 28629 21845 28641 21879
rect 28675 21876 28687 21879
rect 29454 21876 29460 21888
rect 28675 21848 29460 21876
rect 28675 21845 28687 21848
rect 28629 21839 28687 21845
rect 29454 21836 29460 21848
rect 29512 21876 29518 21888
rect 30282 21876 30288 21888
rect 29512 21848 30288 21876
rect 29512 21836 29518 21848
rect 30282 21836 30288 21848
rect 30340 21836 30346 21888
rect 34149 21879 34207 21885
rect 34149 21845 34161 21879
rect 34195 21876 34207 21879
rect 34716 21876 34744 22043
rect 35544 22024 35572 22052
rect 38930 22040 38936 22092
rect 38988 22080 38994 22092
rect 39298 22080 39304 22092
rect 38988 22052 39160 22080
rect 39259 22052 39304 22080
rect 38988 22040 38994 22052
rect 34790 21972 34796 22024
rect 34848 22012 34854 22024
rect 34977 22015 35035 22021
rect 34977 22012 34989 22015
rect 34848 21984 34989 22012
rect 34848 21972 34854 21984
rect 34977 21981 34989 21984
rect 35023 21981 35035 22015
rect 34977 21975 35035 21981
rect 35526 21972 35532 22024
rect 35584 22012 35590 22024
rect 35989 22015 36047 22021
rect 35989 22012 36001 22015
rect 35584 21984 36001 22012
rect 35584 21972 35590 21984
rect 35989 21981 36001 21984
rect 36035 21981 36047 22015
rect 35989 21975 36047 21981
rect 36173 22015 36231 22021
rect 36173 21981 36185 22015
rect 36219 21981 36231 22015
rect 39022 22012 39028 22024
rect 38983 21984 39028 22012
rect 36173 21975 36231 21981
rect 35342 21904 35348 21956
rect 35400 21944 35406 21956
rect 35710 21944 35716 21956
rect 35400 21916 35716 21944
rect 35400 21904 35406 21916
rect 35710 21904 35716 21916
rect 35768 21944 35774 21956
rect 36188 21944 36216 21975
rect 39022 21972 39028 21984
rect 39080 21972 39086 22024
rect 39132 22021 39160 22052
rect 39298 22040 39304 22052
rect 39356 22040 39362 22092
rect 40497 22083 40555 22089
rect 40497 22049 40509 22083
rect 40543 22080 40555 22083
rect 40678 22080 40684 22092
rect 40543 22052 40684 22080
rect 40543 22049 40555 22052
rect 40497 22043 40555 22049
rect 40678 22040 40684 22052
rect 40736 22040 40742 22092
rect 42150 22080 42156 22092
rect 42111 22052 42156 22080
rect 42150 22040 42156 22052
rect 42208 22040 42214 22092
rect 39117 22015 39175 22021
rect 39117 21981 39129 22015
rect 39163 21981 39175 22015
rect 39117 21975 39175 21981
rect 39666 21972 39672 22024
rect 39724 22012 39730 22024
rect 40313 22015 40371 22021
rect 40313 22012 40325 22015
rect 39724 21984 40325 22012
rect 39724 21972 39730 21984
rect 40313 21981 40325 21984
rect 40359 21981 40371 22015
rect 40313 21975 40371 21981
rect 35768 21916 36216 21944
rect 35768 21904 35774 21916
rect 36354 21876 36360 21888
rect 34195 21848 34744 21876
rect 36315 21848 36360 21876
rect 34195 21845 34207 21848
rect 34149 21839 34207 21845
rect 36354 21836 36360 21848
rect 36412 21836 36418 21888
rect 1104 21786 42872 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 42872 21786
rect 1104 21712 42872 21734
rect 14366 21632 14372 21684
rect 14424 21672 14430 21684
rect 14645 21675 14703 21681
rect 14645 21672 14657 21675
rect 14424 21644 14657 21672
rect 14424 21632 14430 21644
rect 14645 21641 14657 21644
rect 14691 21672 14703 21675
rect 16206 21672 16212 21684
rect 14691 21644 16212 21672
rect 14691 21641 14703 21644
rect 14645 21635 14703 21641
rect 16206 21632 16212 21644
rect 16264 21632 16270 21684
rect 20898 21632 20904 21684
rect 20956 21672 20962 21684
rect 22005 21675 22063 21681
rect 22005 21672 22017 21675
rect 20956 21644 22017 21672
rect 20956 21632 20962 21644
rect 22005 21641 22017 21644
rect 22051 21641 22063 21675
rect 22922 21672 22928 21684
rect 22835 21644 22928 21672
rect 22005 21635 22063 21641
rect 22922 21632 22928 21644
rect 22980 21632 22986 21684
rect 24029 21675 24087 21681
rect 24029 21641 24041 21675
rect 24075 21672 24087 21675
rect 24118 21672 24124 21684
rect 24075 21644 24124 21672
rect 24075 21641 24087 21644
rect 24029 21635 24087 21641
rect 24118 21632 24124 21644
rect 24176 21632 24182 21684
rect 24394 21632 24400 21684
rect 24452 21672 24458 21684
rect 25409 21675 25467 21681
rect 25409 21672 25421 21675
rect 24452 21644 25421 21672
rect 24452 21632 24458 21644
rect 25409 21641 25421 21644
rect 25455 21641 25467 21675
rect 26050 21672 26056 21684
rect 26011 21644 26056 21672
rect 25409 21635 25467 21641
rect 26050 21632 26056 21644
rect 26108 21632 26114 21684
rect 28994 21672 29000 21684
rect 26160 21644 29000 21672
rect 19058 21564 19064 21616
rect 19116 21604 19122 21616
rect 19214 21607 19272 21613
rect 19214 21604 19226 21607
rect 19116 21576 19226 21604
rect 19116 21564 19122 21576
rect 19214 21573 19226 21576
rect 19260 21573 19272 21607
rect 19214 21567 19272 21573
rect 20714 21564 20720 21616
rect 20772 21604 20778 21616
rect 21821 21607 21879 21613
rect 21821 21604 21833 21607
rect 20772 21576 21833 21604
rect 20772 21564 20778 21576
rect 21821 21573 21833 21576
rect 21867 21573 21879 21607
rect 21821 21567 21879 21573
rect 21910 21564 21916 21616
rect 21968 21604 21974 21616
rect 22940 21604 22968 21632
rect 26160 21604 26188 21644
rect 28994 21632 29000 21644
rect 29052 21632 29058 21684
rect 29730 21672 29736 21684
rect 29691 21644 29736 21672
rect 29730 21632 29736 21644
rect 29788 21632 29794 21684
rect 32293 21675 32351 21681
rect 32293 21641 32305 21675
rect 32339 21672 32351 21675
rect 32398 21672 32404 21684
rect 32339 21644 32404 21672
rect 32339 21641 32351 21644
rect 32293 21635 32351 21641
rect 32398 21632 32404 21644
rect 32456 21672 32462 21684
rect 32582 21672 32588 21684
rect 32456 21644 32588 21672
rect 32456 21632 32462 21644
rect 32582 21632 32588 21644
rect 32640 21632 32646 21684
rect 38657 21675 38715 21681
rect 38657 21641 38669 21675
rect 38703 21672 38715 21675
rect 38838 21672 38844 21684
rect 38703 21644 38844 21672
rect 38703 21641 38715 21644
rect 38657 21635 38715 21641
rect 38838 21632 38844 21644
rect 38896 21632 38902 21684
rect 27614 21604 27620 21616
rect 21968 21576 22140 21604
rect 22940 21576 26188 21604
rect 27356 21576 27620 21604
rect 21968 21564 21974 21576
rect 6362 21536 6368 21548
rect 6323 21508 6368 21536
rect 6362 21496 6368 21508
rect 6420 21496 6426 21548
rect 14734 21536 14740 21548
rect 14695 21508 14740 21536
rect 14734 21496 14740 21508
rect 14792 21496 14798 21548
rect 15102 21496 15108 21548
rect 15160 21536 15166 21548
rect 15289 21539 15347 21545
rect 15289 21536 15301 21539
rect 15160 21508 15301 21536
rect 15160 21496 15166 21508
rect 15289 21505 15301 21508
rect 15335 21505 15347 21539
rect 15289 21499 15347 21505
rect 15470 21496 15476 21548
rect 15528 21536 15534 21548
rect 16666 21536 16672 21548
rect 15528 21508 16672 21536
rect 15528 21496 15534 21508
rect 16666 21496 16672 21508
rect 16724 21496 16730 21548
rect 16936 21539 16994 21545
rect 16936 21505 16948 21539
rect 16982 21536 16994 21539
rect 17218 21536 17224 21548
rect 16982 21508 17224 21536
rect 16982 21505 16994 21508
rect 16936 21499 16994 21505
rect 17218 21496 17224 21508
rect 17276 21496 17282 21548
rect 18782 21496 18788 21548
rect 18840 21536 18846 21548
rect 22112 21545 22140 21576
rect 18969 21539 19027 21545
rect 18969 21536 18981 21539
rect 18840 21508 18981 21536
rect 18840 21496 18846 21508
rect 18969 21505 18981 21508
rect 19015 21505 19027 21539
rect 18969 21499 19027 21505
rect 22097 21539 22155 21545
rect 22097 21505 22109 21539
rect 22143 21505 22155 21539
rect 22097 21499 22155 21505
rect 22741 21539 22799 21545
rect 22741 21505 22753 21539
rect 22787 21536 22799 21539
rect 23474 21536 23480 21548
rect 22787 21508 23480 21536
rect 22787 21505 22799 21508
rect 22741 21499 22799 21505
rect 23474 21496 23480 21508
rect 23532 21496 23538 21548
rect 24305 21539 24363 21545
rect 24305 21505 24317 21539
rect 24351 21536 24363 21539
rect 24394 21536 24400 21548
rect 24351 21508 24400 21536
rect 24351 21505 24363 21508
rect 24305 21499 24363 21505
rect 24394 21496 24400 21508
rect 24452 21496 24458 21548
rect 24581 21539 24639 21545
rect 24581 21505 24593 21539
rect 24627 21505 24639 21539
rect 24581 21499 24639 21505
rect 1854 21468 1860 21480
rect 1815 21440 1860 21468
rect 1854 21428 1860 21440
rect 1912 21428 1918 21480
rect 2041 21471 2099 21477
rect 2041 21437 2053 21471
rect 2087 21468 2099 21471
rect 2682 21468 2688 21480
rect 2087 21440 2688 21468
rect 2087 21437 2099 21440
rect 2041 21431 2099 21437
rect 2682 21428 2688 21440
rect 2740 21428 2746 21480
rect 2774 21428 2780 21480
rect 2832 21468 2838 21480
rect 7098 21468 7104 21480
rect 2832 21440 2877 21468
rect 7059 21440 7104 21468
rect 2832 21428 2838 21440
rect 7098 21428 7104 21440
rect 7156 21428 7162 21480
rect 15565 21471 15623 21477
rect 15565 21437 15577 21471
rect 15611 21468 15623 21471
rect 15838 21468 15844 21480
rect 15611 21440 15844 21468
rect 15611 21437 15623 21440
rect 15565 21431 15623 21437
rect 15838 21428 15844 21440
rect 15896 21428 15902 21480
rect 24121 21471 24179 21477
rect 24121 21437 24133 21471
rect 24167 21468 24179 21471
rect 24596 21468 24624 21499
rect 24670 21496 24676 21548
rect 24728 21536 24734 21548
rect 27356 21545 27384 21576
rect 27614 21564 27620 21576
rect 27672 21564 27678 21616
rect 28350 21564 28356 21616
rect 28408 21604 28414 21616
rect 30558 21604 30564 21616
rect 28408 21576 28764 21604
rect 28408 21564 28414 21576
rect 25041 21539 25099 21545
rect 25041 21536 25053 21539
rect 24728 21508 25053 21536
rect 24728 21496 24734 21508
rect 25041 21505 25053 21508
rect 25087 21505 25099 21539
rect 25041 21499 25099 21505
rect 25961 21539 26019 21545
rect 25961 21505 25973 21539
rect 26007 21505 26019 21539
rect 25961 21499 26019 21505
rect 27341 21539 27399 21545
rect 27341 21505 27353 21539
rect 27387 21505 27399 21539
rect 27522 21536 27528 21548
rect 27483 21508 27528 21536
rect 27341 21499 27399 21505
rect 24762 21468 24768 21480
rect 24167 21440 24532 21468
rect 24596 21440 24768 21468
rect 24167 21437 24179 21440
rect 24121 21431 24179 21437
rect 21818 21400 21824 21412
rect 21779 21372 21824 21400
rect 21818 21360 21824 21372
rect 21876 21360 21882 21412
rect 17586 21292 17592 21344
rect 17644 21332 17650 21344
rect 18049 21335 18107 21341
rect 18049 21332 18061 21335
rect 17644 21304 18061 21332
rect 17644 21292 17650 21304
rect 18049 21301 18061 21304
rect 18095 21301 18107 21335
rect 18049 21295 18107 21301
rect 20349 21335 20407 21341
rect 20349 21301 20361 21335
rect 20395 21332 20407 21335
rect 20806 21332 20812 21344
rect 20395 21304 20812 21332
rect 20395 21301 20407 21304
rect 20349 21295 20407 21301
rect 20806 21292 20812 21304
rect 20864 21292 20870 21344
rect 24504 21332 24532 21440
rect 24762 21428 24768 21440
rect 24820 21468 24826 21480
rect 25133 21471 25191 21477
rect 25133 21468 25145 21471
rect 24820 21440 25145 21468
rect 24820 21428 24826 21440
rect 25133 21437 25145 21440
rect 25179 21437 25191 21471
rect 25133 21431 25191 21437
rect 24578 21360 24584 21412
rect 24636 21400 24642 21412
rect 25976 21400 26004 21499
rect 27522 21496 27528 21508
rect 27580 21496 27586 21548
rect 28166 21496 28172 21548
rect 28224 21536 28230 21548
rect 28534 21536 28540 21548
rect 28224 21508 28540 21536
rect 28224 21496 28230 21508
rect 28534 21496 28540 21508
rect 28592 21496 28598 21548
rect 28736 21545 28764 21576
rect 29288 21576 30564 21604
rect 29288 21548 29316 21576
rect 30558 21564 30564 21576
rect 30616 21564 30622 21616
rect 32493 21607 32551 21613
rect 32493 21573 32505 21607
rect 32539 21604 32551 21607
rect 33042 21604 33048 21616
rect 32539 21576 33048 21604
rect 32539 21573 32551 21576
rect 32493 21567 32551 21573
rect 33042 21564 33048 21576
rect 33100 21564 33106 21616
rect 35621 21607 35679 21613
rect 35621 21573 35633 21607
rect 35667 21604 35679 21607
rect 41874 21604 41880 21616
rect 35667 21576 36216 21604
rect 41835 21576 41880 21604
rect 35667 21573 35679 21576
rect 35621 21567 35679 21573
rect 28721 21539 28779 21545
rect 28721 21505 28733 21539
rect 28767 21505 28779 21539
rect 29270 21536 29276 21548
rect 29183 21508 29276 21536
rect 28721 21499 28779 21505
rect 29270 21496 29276 21508
rect 29328 21496 29334 21548
rect 29549 21539 29607 21545
rect 29549 21505 29561 21539
rect 29595 21536 29607 21539
rect 30650 21536 30656 21548
rect 29595 21508 30656 21536
rect 29595 21505 29607 21508
rect 29549 21499 29607 21505
rect 30650 21496 30656 21508
rect 30708 21496 30714 21548
rect 35526 21536 35532 21548
rect 35487 21508 35532 21536
rect 35526 21496 35532 21508
rect 35584 21496 35590 21548
rect 35710 21536 35716 21548
rect 35671 21508 35716 21536
rect 35710 21496 35716 21508
rect 35768 21496 35774 21548
rect 36188 21545 36216 21576
rect 41874 21564 41880 21576
rect 41932 21564 41938 21616
rect 36173 21539 36231 21545
rect 36173 21505 36185 21539
rect 36219 21505 36231 21539
rect 36354 21536 36360 21548
rect 36315 21508 36360 21536
rect 36173 21499 36231 21505
rect 36354 21496 36360 21508
rect 36412 21496 36418 21548
rect 38473 21539 38531 21545
rect 38473 21536 38485 21539
rect 38028 21508 38485 21536
rect 27709 21471 27767 21477
rect 27709 21437 27721 21471
rect 27755 21468 27767 21471
rect 28442 21468 28448 21480
rect 27755 21440 28448 21468
rect 27755 21437 27767 21440
rect 27709 21431 27767 21437
rect 28442 21428 28448 21440
rect 28500 21468 28506 21480
rect 33686 21468 33692 21480
rect 28500 21440 33692 21468
rect 28500 21428 28506 21440
rect 33686 21428 33692 21440
rect 33744 21428 33750 21480
rect 37274 21428 37280 21480
rect 37332 21468 37338 21480
rect 38028 21477 38056 21508
rect 38473 21505 38485 21508
rect 38519 21505 38531 21539
rect 38473 21499 38531 21505
rect 39577 21539 39635 21545
rect 39577 21505 39589 21539
rect 39623 21536 39635 21539
rect 39666 21536 39672 21548
rect 39623 21508 39672 21536
rect 39623 21505 39635 21508
rect 39577 21499 39635 21505
rect 39666 21496 39672 21508
rect 39724 21496 39730 21548
rect 37553 21471 37611 21477
rect 37553 21468 37565 21471
rect 37332 21440 37565 21468
rect 37332 21428 37338 21440
rect 37553 21437 37565 21440
rect 37599 21437 37611 21471
rect 37553 21431 37611 21437
rect 38013 21471 38071 21477
rect 38013 21437 38025 21471
rect 38059 21437 38071 21471
rect 38013 21431 38071 21437
rect 39298 21428 39304 21480
rect 39356 21468 39362 21480
rect 40037 21471 40095 21477
rect 40037 21468 40049 21471
rect 39356 21440 40049 21468
rect 39356 21428 39362 21440
rect 40037 21437 40049 21440
rect 40083 21437 40095 21471
rect 40037 21431 40095 21437
rect 40221 21471 40279 21477
rect 40221 21437 40233 21471
rect 40267 21468 40279 21471
rect 40954 21468 40960 21480
rect 40267 21440 40960 21468
rect 40267 21437 40279 21440
rect 40221 21431 40279 21437
rect 40954 21428 40960 21440
rect 41012 21428 41018 21480
rect 24636 21372 26004 21400
rect 24636 21360 24642 21372
rect 27890 21360 27896 21412
rect 27948 21400 27954 21412
rect 29365 21403 29423 21409
rect 29365 21400 29377 21403
rect 27948 21372 29377 21400
rect 27948 21360 27954 21372
rect 29365 21369 29377 21372
rect 29411 21369 29423 21403
rect 29365 21363 29423 21369
rect 29457 21403 29515 21409
rect 29457 21369 29469 21403
rect 29503 21400 29515 21403
rect 30282 21400 30288 21412
rect 29503 21372 30288 21400
rect 29503 21369 29515 21372
rect 29457 21363 29515 21369
rect 30282 21360 30288 21372
rect 30340 21360 30346 21412
rect 32125 21403 32183 21409
rect 32125 21369 32137 21403
rect 32171 21400 32183 21403
rect 32490 21400 32496 21412
rect 32171 21372 32496 21400
rect 32171 21369 32183 21372
rect 32125 21363 32183 21369
rect 32490 21360 32496 21372
rect 32548 21360 32554 21412
rect 37921 21403 37979 21409
rect 37921 21369 37933 21403
rect 37967 21400 37979 21403
rect 38470 21400 38476 21412
rect 37967 21372 38476 21400
rect 37967 21369 37979 21372
rect 37921 21363 37979 21369
rect 38470 21360 38476 21372
rect 38528 21360 38534 21412
rect 24670 21332 24676 21344
rect 24504 21304 24676 21332
rect 24670 21292 24676 21304
rect 24728 21292 24734 21344
rect 25130 21332 25136 21344
rect 25091 21304 25136 21332
rect 25130 21292 25136 21304
rect 25188 21292 25194 21344
rect 28721 21335 28779 21341
rect 28721 21301 28733 21335
rect 28767 21332 28779 21335
rect 29270 21332 29276 21344
rect 28767 21304 29276 21332
rect 28767 21301 28779 21304
rect 28721 21295 28779 21301
rect 29270 21292 29276 21304
rect 29328 21292 29334 21344
rect 32214 21292 32220 21344
rect 32272 21332 32278 21344
rect 32309 21335 32367 21341
rect 32309 21332 32321 21335
rect 32272 21304 32321 21332
rect 32272 21292 32278 21304
rect 32309 21301 32321 21304
rect 32355 21332 32367 21335
rect 34790 21332 34796 21344
rect 32355 21304 34796 21332
rect 32355 21301 32367 21304
rect 32309 21295 32367 21301
rect 34790 21292 34796 21304
rect 34848 21292 34854 21344
rect 36170 21332 36176 21344
rect 36131 21304 36176 21332
rect 36170 21292 36176 21304
rect 36228 21292 36234 21344
rect 1104 21242 42872 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 42872 21242
rect 1104 21168 42872 21190
rect 1854 21088 1860 21140
rect 1912 21128 1918 21140
rect 1949 21131 2007 21137
rect 1949 21128 1961 21131
rect 1912 21100 1961 21128
rect 1912 21088 1918 21100
rect 1949 21097 1961 21100
rect 1995 21097 2007 21131
rect 2682 21128 2688 21140
rect 2643 21100 2688 21128
rect 1949 21091 2007 21097
rect 2682 21088 2688 21100
rect 2740 21088 2746 21140
rect 7466 21128 7472 21140
rect 7427 21100 7472 21128
rect 7466 21088 7472 21100
rect 7524 21128 7530 21140
rect 8110 21128 8116 21140
rect 7524 21100 8116 21128
rect 7524 21088 7530 21100
rect 8110 21088 8116 21100
rect 8168 21088 8174 21140
rect 15378 21088 15384 21140
rect 15436 21128 15442 21140
rect 15473 21131 15531 21137
rect 15473 21128 15485 21131
rect 15436 21100 15485 21128
rect 15436 21088 15442 21100
rect 15473 21097 15485 21100
rect 15519 21097 15531 21131
rect 17218 21128 17224 21140
rect 17179 21100 17224 21128
rect 15473 21091 15531 21097
rect 17218 21088 17224 21100
rect 17276 21088 17282 21140
rect 20806 21128 20812 21140
rect 17328 21100 17816 21128
rect 20767 21100 20812 21128
rect 16206 21060 16212 21072
rect 15764 21032 16212 21060
rect 13449 20995 13507 21001
rect 13449 20961 13461 20995
rect 13495 20992 13507 20995
rect 13495 20964 14596 20992
rect 13495 20961 13507 20964
rect 13449 20955 13507 20961
rect 2777 20927 2835 20933
rect 2777 20893 2789 20927
rect 2823 20924 2835 20927
rect 3326 20924 3332 20936
rect 2823 20896 3332 20924
rect 2823 20893 2835 20896
rect 2777 20887 2835 20893
rect 3326 20884 3332 20896
rect 3384 20924 3390 20936
rect 5718 20924 5724 20936
rect 3384 20896 5488 20924
rect 5631 20896 5724 20924
rect 3384 20884 3390 20896
rect 5460 20868 5488 20896
rect 5718 20884 5724 20896
rect 5776 20924 5782 20936
rect 6181 20927 6239 20933
rect 6181 20924 6193 20927
rect 5776 20896 6193 20924
rect 5776 20884 5782 20896
rect 6181 20893 6193 20896
rect 6227 20924 6239 20927
rect 6362 20924 6368 20936
rect 6227 20896 6368 20924
rect 6227 20893 6239 20896
rect 6181 20887 6239 20893
rect 6362 20884 6368 20896
rect 6420 20884 6426 20936
rect 13357 20927 13415 20933
rect 13357 20893 13369 20927
rect 13403 20893 13415 20927
rect 13357 20887 13415 20893
rect 13541 20927 13599 20933
rect 13541 20893 13553 20927
rect 13587 20924 13599 20927
rect 14366 20924 14372 20936
rect 13587 20896 14372 20924
rect 13587 20893 13599 20896
rect 13541 20887 13599 20893
rect 5442 20856 5448 20868
rect 5403 20828 5448 20856
rect 5442 20816 5448 20828
rect 5500 20816 5506 20868
rect 13372 20856 13400 20887
rect 14366 20884 14372 20896
rect 14424 20884 14430 20936
rect 14568 20933 14596 20964
rect 14461 20927 14519 20933
rect 14461 20893 14473 20927
rect 14507 20893 14519 20927
rect 14461 20887 14519 20893
rect 14553 20927 14611 20933
rect 14553 20893 14565 20927
rect 14599 20893 14611 20927
rect 14553 20887 14611 20893
rect 14476 20856 14504 20887
rect 14642 20884 14648 20936
rect 14700 20924 14706 20936
rect 14737 20927 14795 20933
rect 14737 20924 14749 20927
rect 14700 20896 14749 20924
rect 14700 20884 14706 20896
rect 14737 20893 14749 20896
rect 14783 20893 14795 20927
rect 15654 20924 15660 20936
rect 15615 20896 15660 20924
rect 14737 20887 14795 20893
rect 15654 20884 15660 20896
rect 15712 20884 15718 20936
rect 15764 20924 15792 21032
rect 16206 21020 16212 21032
rect 16264 21060 16270 21072
rect 16850 21060 16856 21072
rect 16264 21032 16856 21060
rect 16264 21020 16270 21032
rect 16850 21020 16856 21032
rect 16908 21060 16914 21072
rect 17328 21060 17356 21100
rect 17678 21060 17684 21072
rect 16908 21032 17356 21060
rect 17639 21032 17684 21060
rect 16908 21020 16914 21032
rect 17678 21020 17684 21032
rect 17736 21020 17742 21072
rect 17788 21060 17816 21100
rect 20806 21088 20812 21100
rect 20864 21088 20870 21140
rect 24394 21088 24400 21140
rect 24452 21128 24458 21140
rect 25130 21128 25136 21140
rect 24452 21100 25136 21128
rect 24452 21088 24458 21100
rect 25130 21088 25136 21100
rect 25188 21088 25194 21140
rect 28626 21088 28632 21140
rect 28684 21088 28690 21140
rect 28905 21131 28963 21137
rect 28905 21097 28917 21131
rect 28951 21128 28963 21131
rect 29086 21128 29092 21140
rect 28951 21100 29092 21128
rect 28951 21097 28963 21100
rect 28905 21091 28963 21097
rect 29086 21088 29092 21100
rect 29144 21088 29150 21140
rect 31021 21131 31079 21137
rect 31021 21128 31033 21131
rect 30392 21100 31033 21128
rect 21818 21060 21824 21072
rect 17788 21032 21824 21060
rect 21818 21020 21824 21032
rect 21876 21020 21882 21072
rect 27065 21063 27123 21069
rect 27065 21029 27077 21063
rect 27111 21060 27123 21063
rect 27338 21060 27344 21072
rect 27111 21032 27344 21060
rect 27111 21029 27123 21032
rect 27065 21023 27123 21029
rect 27338 21020 27344 21032
rect 27396 21020 27402 21072
rect 28442 21020 28448 21072
rect 28500 21060 28506 21072
rect 28644 21060 28672 21088
rect 30392 21060 30420 21100
rect 31021 21097 31033 21100
rect 31067 21097 31079 21131
rect 32398 21128 32404 21140
rect 31021 21091 31079 21097
rect 31220 21100 32404 21128
rect 28500 21032 30420 21060
rect 30653 21063 30711 21069
rect 28500 21020 28506 21032
rect 30653 21029 30665 21063
rect 30699 21060 30711 21063
rect 31220 21060 31248 21100
rect 32398 21088 32404 21100
rect 32456 21088 32462 21140
rect 33686 21088 33692 21140
rect 33744 21128 33750 21140
rect 34514 21128 34520 21140
rect 33744 21100 34520 21128
rect 33744 21088 33750 21100
rect 34514 21088 34520 21100
rect 34572 21128 34578 21140
rect 37182 21128 37188 21140
rect 34572 21100 35020 21128
rect 37143 21100 37188 21128
rect 34572 21088 34578 21100
rect 33042 21060 33048 21072
rect 30699 21032 31248 21060
rect 32955 21032 33048 21060
rect 30699 21029 30711 21032
rect 30653 21023 30711 21029
rect 33042 21020 33048 21032
rect 33100 21060 33106 21072
rect 34992 21060 35020 21100
rect 37182 21088 37188 21100
rect 37240 21088 37246 21140
rect 38010 21088 38016 21140
rect 38068 21128 38074 21140
rect 38105 21131 38163 21137
rect 38105 21128 38117 21131
rect 38068 21100 38117 21128
rect 38068 21088 38074 21100
rect 38105 21097 38117 21100
rect 38151 21097 38163 21131
rect 39298 21128 39304 21140
rect 39259 21100 39304 21128
rect 38105 21091 38163 21097
rect 39298 21088 39304 21100
rect 39356 21088 39362 21140
rect 40954 21128 40960 21140
rect 40915 21100 40960 21128
rect 40954 21088 40960 21100
rect 41012 21088 41018 21140
rect 41601 21131 41659 21137
rect 41601 21097 41613 21131
rect 41647 21128 41659 21131
rect 41690 21128 41696 21140
rect 41647 21100 41696 21128
rect 41647 21097 41659 21100
rect 41601 21091 41659 21097
rect 41690 21088 41696 21100
rect 41748 21088 41754 21140
rect 36265 21063 36323 21069
rect 33100 21032 33824 21060
rect 34992 21032 35112 21060
rect 33100 21020 33106 21032
rect 15838 20952 15844 21004
rect 15896 20992 15902 21004
rect 16117 20995 16175 21001
rect 16117 20992 16129 20995
rect 15896 20964 16129 20992
rect 15896 20952 15902 20964
rect 16117 20961 16129 20964
rect 16163 20992 16175 20995
rect 16163 20964 17816 20992
rect 16163 20961 16175 20964
rect 16117 20955 16175 20961
rect 16574 20924 16580 20936
rect 15764 20896 15884 20924
rect 16535 20896 16580 20924
rect 15010 20856 15016 20868
rect 13372 20828 14412 20856
rect 14476 20828 15016 20856
rect 14090 20788 14096 20800
rect 14051 20760 14096 20788
rect 14090 20748 14096 20760
rect 14148 20748 14154 20800
rect 14384 20788 14412 20828
rect 15010 20816 15016 20828
rect 15068 20856 15074 20868
rect 15856 20865 15884 20896
rect 16574 20884 16580 20896
rect 16632 20884 16638 20936
rect 16850 20884 16856 20936
rect 16908 20924 16914 20936
rect 17037 20927 17095 20933
rect 16908 20896 16952 20924
rect 16908 20884 16914 20896
rect 17037 20893 17049 20927
rect 17083 20924 17095 20927
rect 17126 20924 17132 20936
rect 17083 20896 17132 20924
rect 17083 20893 17095 20896
rect 17037 20887 17095 20893
rect 17126 20884 17132 20896
rect 17184 20884 17190 20936
rect 15749 20859 15807 20865
rect 15749 20856 15761 20859
rect 15068 20828 15761 20856
rect 15068 20816 15074 20828
rect 15749 20825 15761 20828
rect 15795 20825 15807 20859
rect 15749 20819 15807 20825
rect 15841 20859 15899 20865
rect 15841 20825 15853 20859
rect 15887 20825 15899 20859
rect 15841 20819 15899 20825
rect 15979 20859 16037 20865
rect 15979 20825 15991 20859
rect 16025 20856 16037 20859
rect 16298 20856 16304 20868
rect 16025 20828 16304 20856
rect 16025 20825 16037 20828
rect 15979 20819 16037 20825
rect 15562 20788 15568 20800
rect 14384 20760 15568 20788
rect 15562 20748 15568 20760
rect 15620 20748 15626 20800
rect 15764 20788 15792 20819
rect 16298 20816 16304 20828
rect 16356 20856 16362 20868
rect 16715 20859 16773 20865
rect 16715 20856 16727 20859
rect 16356 20828 16727 20856
rect 16356 20816 16362 20828
rect 16715 20825 16727 20828
rect 16761 20825 16773 20859
rect 16715 20819 16773 20825
rect 16945 20859 17003 20865
rect 16945 20825 16957 20859
rect 16991 20825 17003 20859
rect 16945 20819 17003 20825
rect 16960 20788 16988 20819
rect 17586 20816 17592 20868
rect 17644 20856 17650 20868
rect 17681 20859 17739 20865
rect 17681 20856 17693 20859
rect 17644 20828 17693 20856
rect 17644 20816 17650 20828
rect 17681 20825 17693 20828
rect 17727 20825 17739 20859
rect 17788 20856 17816 20964
rect 20714 20952 20720 21004
rect 20772 20992 20778 21004
rect 20901 20995 20959 21001
rect 20901 20992 20913 20995
rect 20772 20964 20913 20992
rect 20772 20952 20778 20964
rect 20901 20961 20913 20964
rect 20947 20961 20959 20995
rect 20901 20955 20959 20961
rect 25501 20995 25559 21001
rect 25501 20961 25513 20995
rect 25547 20992 25559 20995
rect 25958 20992 25964 21004
rect 25547 20964 25964 20992
rect 25547 20961 25559 20964
rect 25501 20955 25559 20961
rect 25958 20952 25964 20964
rect 26016 20952 26022 21004
rect 33686 20992 33692 21004
rect 33647 20964 33692 20992
rect 33686 20952 33692 20964
rect 33744 20952 33750 21004
rect 33796 20992 33824 21032
rect 33796 20964 35020 20992
rect 17954 20924 17960 20936
rect 17915 20896 17960 20924
rect 17954 20884 17960 20896
rect 18012 20884 18018 20936
rect 19245 20927 19303 20933
rect 19245 20893 19257 20927
rect 19291 20893 19303 20927
rect 19245 20887 19303 20893
rect 19429 20927 19487 20933
rect 19429 20893 19441 20927
rect 19475 20893 19487 20927
rect 19429 20887 19487 20893
rect 19613 20927 19671 20933
rect 19613 20893 19625 20927
rect 19659 20924 19671 20927
rect 20257 20927 20315 20933
rect 20257 20924 20269 20927
rect 19659 20896 20269 20924
rect 19659 20893 19671 20896
rect 19613 20887 19671 20893
rect 20257 20893 20269 20896
rect 20303 20893 20315 20927
rect 21082 20924 21088 20936
rect 21043 20896 21088 20924
rect 20257 20887 20315 20893
rect 17865 20859 17923 20865
rect 17865 20856 17877 20859
rect 17788 20828 17877 20856
rect 17681 20819 17739 20825
rect 17865 20825 17877 20828
rect 17911 20856 17923 20859
rect 19260 20856 19288 20887
rect 17911 20828 19288 20856
rect 19444 20856 19472 20887
rect 21082 20884 21088 20896
rect 21140 20884 21146 20936
rect 21913 20927 21971 20933
rect 21913 20893 21925 20927
rect 21959 20924 21971 20927
rect 23474 20924 23480 20936
rect 21959 20896 23480 20924
rect 21959 20893 21971 20896
rect 21913 20887 21971 20893
rect 23474 20884 23480 20896
rect 23532 20884 23538 20936
rect 24578 20924 24584 20936
rect 24539 20896 24584 20924
rect 24578 20884 24584 20896
rect 24636 20884 24642 20936
rect 25038 20884 25044 20936
rect 25096 20924 25102 20936
rect 25225 20927 25283 20933
rect 25225 20924 25237 20927
rect 25096 20896 25237 20924
rect 25096 20884 25102 20896
rect 25225 20893 25237 20896
rect 25271 20893 25283 20927
rect 27062 20924 27068 20936
rect 27023 20896 27068 20924
rect 25225 20887 25283 20893
rect 27062 20884 27068 20896
rect 27120 20884 27126 20936
rect 27249 20927 27307 20933
rect 27249 20893 27261 20927
rect 27295 20924 27307 20927
rect 27614 20924 27620 20936
rect 27295 20896 27620 20924
rect 27295 20893 27307 20896
rect 27249 20887 27307 20893
rect 27614 20884 27620 20896
rect 27672 20924 27678 20936
rect 27672 20896 27844 20924
rect 27672 20884 27678 20896
rect 19978 20856 19984 20868
rect 19444 20828 19984 20856
rect 17911 20825 17923 20828
rect 17865 20819 17923 20825
rect 19978 20816 19984 20828
rect 20036 20816 20042 20868
rect 20806 20856 20812 20868
rect 20767 20828 20812 20856
rect 20806 20816 20812 20828
rect 20864 20816 20870 20868
rect 24765 20859 24823 20865
rect 24765 20825 24777 20859
rect 24811 20856 24823 20859
rect 24854 20856 24860 20868
rect 24811 20828 24860 20856
rect 24811 20825 24823 20828
rect 24765 20819 24823 20825
rect 24854 20816 24860 20828
rect 24912 20816 24918 20868
rect 26694 20856 26700 20868
rect 26655 20828 26700 20856
rect 26694 20816 26700 20828
rect 26752 20816 26758 20868
rect 27709 20859 27767 20865
rect 27709 20856 27721 20859
rect 27632 20828 27721 20856
rect 27632 20800 27660 20828
rect 27709 20825 27721 20828
rect 27755 20825 27767 20859
rect 27816 20856 27844 20896
rect 27890 20884 27896 20936
rect 27948 20924 27954 20936
rect 28718 20924 28724 20936
rect 27948 20896 27993 20924
rect 28679 20896 28724 20924
rect 27948 20884 27954 20896
rect 28718 20884 28724 20896
rect 28776 20884 28782 20936
rect 28810 20884 28816 20936
rect 28868 20924 28874 20936
rect 28905 20927 28963 20933
rect 28905 20924 28917 20927
rect 28868 20896 28917 20924
rect 28868 20884 28874 20896
rect 28905 20893 28917 20896
rect 28951 20893 28963 20927
rect 28905 20887 28963 20893
rect 31665 20927 31723 20933
rect 31665 20893 31677 20927
rect 31711 20924 31723 20927
rect 32306 20924 32312 20936
rect 31711 20896 32312 20924
rect 31711 20893 31723 20896
rect 31665 20887 31723 20893
rect 32306 20884 32312 20896
rect 32364 20884 32370 20936
rect 33796 20933 33824 20964
rect 33781 20927 33839 20933
rect 33781 20893 33793 20927
rect 33827 20893 33839 20927
rect 33781 20887 33839 20893
rect 34701 20927 34759 20933
rect 34701 20893 34713 20927
rect 34747 20924 34759 20927
rect 34790 20924 34796 20936
rect 34747 20896 34796 20924
rect 34747 20893 34759 20896
rect 34701 20887 34759 20893
rect 34790 20884 34796 20896
rect 34848 20884 34854 20936
rect 34992 20933 35020 20964
rect 35084 20933 35112 21032
rect 36265 21029 36277 21063
rect 36311 21060 36323 21063
rect 36311 21032 36860 21060
rect 36311 21029 36323 21032
rect 36265 21023 36323 21029
rect 35989 20995 36047 21001
rect 35989 20961 36001 20995
rect 36035 20992 36047 20995
rect 36354 20992 36360 21004
rect 36035 20964 36360 20992
rect 36035 20961 36047 20964
rect 35989 20955 36047 20961
rect 36354 20952 36360 20964
rect 36412 20952 36418 21004
rect 36832 21001 36860 21032
rect 36817 20995 36875 21001
rect 36817 20961 36829 20995
rect 36863 20961 36875 20995
rect 36817 20955 36875 20961
rect 37001 20995 37059 21001
rect 37001 20961 37013 20995
rect 37047 20992 37059 20995
rect 37182 20992 37188 21004
rect 37047 20964 37188 20992
rect 37047 20961 37059 20964
rect 37001 20955 37059 20961
rect 34977 20927 35035 20933
rect 34977 20893 34989 20927
rect 35023 20893 35035 20927
rect 34977 20887 35035 20893
rect 35069 20927 35127 20933
rect 35069 20893 35081 20927
rect 35115 20893 35127 20927
rect 35897 20927 35955 20933
rect 35897 20924 35909 20927
rect 35069 20887 35127 20893
rect 35176 20896 35909 20924
rect 28077 20859 28135 20865
rect 28077 20856 28089 20859
rect 27816 20828 28089 20856
rect 27709 20819 27767 20825
rect 28077 20825 28089 20828
rect 28123 20856 28135 20859
rect 28166 20856 28172 20868
rect 28123 20828 28172 20856
rect 28123 20825 28135 20828
rect 28077 20819 28135 20825
rect 28166 20816 28172 20828
rect 28224 20816 28230 20868
rect 31021 20859 31079 20865
rect 31021 20825 31033 20859
rect 31067 20856 31079 20859
rect 31067 20828 31524 20856
rect 31067 20825 31079 20828
rect 31021 20819 31079 20825
rect 20070 20788 20076 20800
rect 15764 20760 16988 20788
rect 20031 20760 20076 20788
rect 20070 20748 20076 20760
rect 20128 20748 20134 20800
rect 21266 20788 21272 20800
rect 21227 20760 21272 20788
rect 21266 20748 21272 20760
rect 21324 20748 21330 20800
rect 21818 20788 21824 20800
rect 21779 20760 21824 20788
rect 21818 20748 21824 20760
rect 21876 20748 21882 20800
rect 27614 20788 27620 20800
rect 27527 20760 27620 20788
rect 27614 20748 27620 20760
rect 27672 20788 27678 20800
rect 30282 20788 30288 20800
rect 27672 20760 30288 20788
rect 27672 20748 27678 20760
rect 30282 20748 30288 20760
rect 30340 20748 30346 20800
rect 31205 20791 31263 20797
rect 31205 20757 31217 20791
rect 31251 20788 31263 20791
rect 31386 20788 31392 20800
rect 31251 20760 31392 20788
rect 31251 20757 31263 20760
rect 31205 20751 31263 20757
rect 31386 20748 31392 20760
rect 31444 20748 31450 20800
rect 31496 20788 31524 20828
rect 31570 20816 31576 20868
rect 31628 20856 31634 20868
rect 31910 20859 31968 20865
rect 31910 20856 31922 20859
rect 31628 20828 31922 20856
rect 31628 20816 31634 20828
rect 31910 20825 31922 20828
rect 31956 20825 31968 20859
rect 34882 20856 34888 20868
rect 34843 20828 34888 20856
rect 31910 20819 31968 20825
rect 34882 20816 34888 20828
rect 34940 20816 34946 20868
rect 32122 20788 32128 20800
rect 31496 20760 32128 20788
rect 32122 20748 32128 20760
rect 32180 20748 32186 20800
rect 34054 20748 34060 20800
rect 34112 20788 34118 20800
rect 34149 20791 34207 20797
rect 34149 20788 34161 20791
rect 34112 20760 34161 20788
rect 34112 20748 34118 20760
rect 34149 20757 34161 20760
rect 34195 20788 34207 20791
rect 35176 20788 35204 20896
rect 35897 20893 35909 20896
rect 35943 20924 35955 20927
rect 36262 20924 36268 20936
rect 35943 20896 36268 20924
rect 35943 20893 35955 20896
rect 35897 20887 35955 20893
rect 36262 20884 36268 20896
rect 36320 20884 36326 20936
rect 36832 20868 36860 20955
rect 37182 20952 37188 20964
rect 37240 20992 37246 21004
rect 37240 20964 37780 20992
rect 37240 20952 37246 20964
rect 36906 20884 36912 20936
rect 36964 20924 36970 20936
rect 37752 20933 37780 20964
rect 38746 20952 38752 21004
rect 38804 20992 38810 21004
rect 38804 20964 40264 20992
rect 38804 20952 38810 20964
rect 37645 20927 37703 20933
rect 36964 20896 37009 20924
rect 36964 20884 36970 20896
rect 37645 20893 37657 20927
rect 37691 20893 37703 20927
rect 37645 20887 37703 20893
rect 37737 20927 37795 20933
rect 37737 20893 37749 20927
rect 37783 20893 37795 20927
rect 37918 20924 37924 20936
rect 37879 20896 37924 20924
rect 37737 20887 37795 20893
rect 36814 20856 36820 20868
rect 36727 20828 36820 20856
rect 36814 20816 36820 20828
rect 36872 20856 36878 20868
rect 37660 20856 37688 20887
rect 37918 20884 37924 20896
rect 37976 20884 37982 20936
rect 40236 20933 40264 20964
rect 39117 20927 39175 20933
rect 39117 20893 39129 20927
rect 39163 20924 39175 20927
rect 40037 20927 40095 20933
rect 40037 20924 40049 20927
rect 39163 20896 40049 20924
rect 39163 20893 39175 20896
rect 39117 20887 39175 20893
rect 40037 20893 40049 20896
rect 40083 20893 40095 20927
rect 40037 20887 40095 20893
rect 40221 20927 40279 20933
rect 40221 20893 40233 20927
rect 40267 20893 40279 20927
rect 40221 20887 40279 20893
rect 40310 20884 40316 20936
rect 40368 20924 40374 20936
rect 40862 20924 40868 20936
rect 40368 20896 40413 20924
rect 40823 20896 40868 20924
rect 40368 20884 40374 20896
rect 40862 20884 40868 20896
rect 40920 20884 40926 20936
rect 41506 20924 41512 20936
rect 41467 20896 41512 20924
rect 41506 20884 41512 20896
rect 41564 20884 41570 20936
rect 37826 20856 37832 20868
rect 36872 20828 37832 20856
rect 36872 20816 36878 20828
rect 37826 20816 37832 20828
rect 37884 20816 37890 20868
rect 34195 20760 35204 20788
rect 35253 20791 35311 20797
rect 34195 20757 34207 20760
rect 34149 20751 34207 20757
rect 35253 20757 35265 20791
rect 35299 20788 35311 20791
rect 35342 20788 35348 20800
rect 35299 20760 35348 20788
rect 35299 20757 35311 20760
rect 35253 20751 35311 20757
rect 35342 20748 35348 20760
rect 35400 20748 35406 20800
rect 1104 20698 42872 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 42872 20698
rect 1104 20624 42872 20646
rect 5718 20584 5724 20596
rect 5679 20556 5724 20584
rect 5718 20544 5724 20556
rect 5776 20544 5782 20596
rect 16945 20587 17003 20593
rect 14476 20556 15240 20584
rect 10318 20516 10324 20528
rect 5552 20488 10324 20516
rect 5552 20460 5580 20488
rect 10318 20476 10324 20488
rect 10376 20476 10382 20528
rect 13164 20519 13222 20525
rect 13164 20485 13176 20519
rect 13210 20516 13222 20519
rect 14090 20516 14096 20528
rect 13210 20488 14096 20516
rect 13210 20485 13222 20488
rect 13164 20479 13222 20485
rect 14090 20476 14096 20488
rect 14148 20476 14154 20528
rect 5534 20448 5540 20460
rect 5495 20420 5540 20448
rect 5534 20408 5540 20420
rect 5592 20408 5598 20460
rect 6362 20448 6368 20460
rect 6323 20420 6368 20448
rect 6362 20408 6368 20420
rect 6420 20408 6426 20460
rect 8110 20408 8116 20460
rect 8168 20448 8174 20460
rect 14476 20448 14504 20556
rect 14826 20516 14832 20528
rect 14787 20488 14832 20516
rect 14826 20476 14832 20488
rect 14884 20476 14890 20528
rect 15212 20516 15240 20556
rect 16945 20553 16957 20587
rect 16991 20584 17003 20587
rect 17126 20584 17132 20596
rect 16991 20556 17132 20584
rect 16991 20553 17003 20556
rect 16945 20547 17003 20553
rect 17126 20544 17132 20556
rect 17184 20544 17190 20596
rect 20993 20587 21051 20593
rect 20993 20553 21005 20587
rect 21039 20584 21051 20587
rect 21082 20584 21088 20596
rect 21039 20556 21088 20584
rect 21039 20553 21051 20556
rect 20993 20547 21051 20553
rect 21082 20544 21088 20556
rect 21140 20544 21146 20596
rect 24210 20584 24216 20596
rect 24171 20556 24216 20584
rect 24210 20544 24216 20556
rect 24268 20544 24274 20596
rect 24762 20584 24768 20596
rect 24723 20556 24768 20584
rect 24762 20544 24768 20556
rect 24820 20544 24826 20596
rect 27522 20584 27528 20596
rect 24964 20556 25360 20584
rect 27483 20556 27528 20584
rect 19880 20519 19938 20525
rect 15059 20485 15117 20491
rect 15212 20488 19334 20516
rect 15059 20482 15071 20485
rect 8168 20420 14504 20448
rect 15044 20451 15071 20482
rect 15105 20451 15117 20485
rect 15044 20445 15117 20451
rect 15657 20451 15715 20457
rect 8168 20408 8174 20420
rect 7193 20383 7251 20389
rect 7193 20349 7205 20383
rect 7239 20380 7251 20383
rect 7650 20380 7656 20392
rect 7239 20352 7656 20380
rect 7239 20349 7251 20352
rect 7193 20343 7251 20349
rect 7650 20340 7656 20352
rect 7708 20340 7714 20392
rect 12894 20380 12900 20392
rect 12855 20352 12900 20380
rect 12894 20340 12900 20352
rect 12952 20340 12958 20392
rect 15044 20380 15072 20445
rect 15657 20417 15669 20451
rect 15703 20417 15715 20451
rect 15657 20411 15715 20417
rect 15672 20380 15700 20411
rect 16022 20408 16028 20460
rect 16080 20448 16086 20460
rect 16853 20451 16911 20457
rect 16853 20448 16865 20451
rect 16080 20420 16865 20448
rect 16080 20408 16086 20420
rect 16853 20417 16865 20420
rect 16899 20417 16911 20451
rect 16853 20411 16911 20417
rect 17037 20451 17095 20457
rect 17037 20417 17049 20451
rect 17083 20448 17095 20451
rect 17678 20448 17684 20460
rect 17083 20420 17684 20448
rect 17083 20417 17095 20420
rect 17037 20411 17095 20417
rect 17678 20408 17684 20420
rect 17736 20408 17742 20460
rect 18693 20451 18751 20457
rect 18693 20417 18705 20451
rect 18739 20417 18751 20451
rect 19306 20448 19334 20488
rect 19880 20485 19892 20519
rect 19926 20516 19938 20519
rect 20070 20516 20076 20528
rect 19926 20488 20076 20516
rect 19926 20485 19938 20488
rect 19880 20479 19938 20485
rect 20070 20476 20076 20488
rect 20128 20476 20134 20528
rect 24228 20516 24256 20544
rect 24964 20516 24992 20556
rect 24228 20488 24992 20516
rect 25038 20476 25044 20528
rect 25096 20516 25102 20528
rect 25225 20519 25283 20525
rect 25225 20516 25237 20519
rect 25096 20488 25237 20516
rect 25096 20476 25102 20488
rect 25225 20485 25237 20488
rect 25271 20485 25283 20519
rect 25225 20479 25283 20485
rect 23934 20448 23940 20460
rect 19306 20420 23940 20448
rect 18693 20411 18751 20417
rect 14752 20352 15700 20380
rect 15749 20383 15807 20389
rect 14752 20324 14780 20352
rect 15749 20349 15761 20383
rect 15795 20380 15807 20383
rect 16114 20380 16120 20392
rect 15795 20352 16120 20380
rect 15795 20349 15807 20352
rect 15749 20343 15807 20349
rect 16114 20340 16120 20352
rect 16172 20340 16178 20392
rect 17586 20340 17592 20392
rect 17644 20380 17650 20392
rect 17954 20380 17960 20392
rect 17644 20352 17960 20380
rect 17644 20340 17650 20352
rect 17954 20340 17960 20352
rect 18012 20380 18018 20392
rect 18509 20383 18567 20389
rect 18509 20380 18521 20383
rect 18012 20352 18521 20380
rect 18012 20340 18018 20352
rect 18509 20349 18521 20352
rect 18555 20349 18567 20383
rect 18708 20380 18736 20411
rect 23934 20408 23940 20420
rect 23992 20408 23998 20460
rect 24118 20448 24124 20460
rect 24079 20420 24124 20448
rect 24118 20408 24124 20420
rect 24176 20408 24182 20460
rect 24302 20448 24308 20460
rect 24263 20420 24308 20448
rect 24302 20408 24308 20420
rect 24360 20408 24366 20460
rect 24854 20408 24860 20460
rect 24912 20448 24918 20460
rect 24949 20451 25007 20457
rect 24949 20448 24961 20451
rect 24912 20420 24961 20448
rect 24912 20408 24918 20420
rect 24949 20417 24961 20420
rect 24995 20448 25007 20451
rect 25332 20448 25360 20556
rect 27522 20544 27528 20556
rect 27580 20544 27586 20596
rect 28721 20587 28779 20593
rect 28721 20553 28733 20587
rect 28767 20553 28779 20587
rect 28721 20547 28779 20553
rect 27065 20519 27123 20525
rect 27065 20485 27077 20519
rect 27111 20516 27123 20519
rect 27614 20516 27620 20528
rect 27111 20488 27620 20516
rect 27111 20485 27123 20488
rect 27065 20479 27123 20485
rect 26237 20451 26295 20457
rect 26237 20448 26249 20451
rect 24995 20420 25268 20448
rect 25332 20420 26249 20448
rect 24995 20417 25007 20420
rect 24949 20411 25007 20417
rect 18708 20352 19012 20380
rect 18509 20343 18567 20349
rect 14277 20315 14335 20321
rect 14277 20281 14289 20315
rect 14323 20312 14335 20315
rect 14734 20312 14740 20324
rect 14323 20284 14740 20312
rect 14323 20281 14335 20284
rect 14277 20275 14335 20281
rect 14734 20272 14740 20284
rect 14792 20272 14798 20324
rect 15197 20315 15255 20321
rect 15197 20281 15209 20315
rect 15243 20312 15255 20315
rect 16574 20312 16580 20324
rect 15243 20284 16580 20312
rect 15243 20281 15255 20284
rect 15197 20275 15255 20281
rect 16574 20272 16580 20284
rect 16632 20272 16638 20324
rect 1394 20204 1400 20256
rect 1452 20244 1458 20256
rect 1673 20247 1731 20253
rect 1673 20244 1685 20247
rect 1452 20216 1685 20244
rect 1452 20204 1458 20216
rect 1673 20213 1685 20216
rect 1719 20213 1731 20247
rect 1673 20207 1731 20213
rect 15013 20247 15071 20253
rect 15013 20213 15025 20247
rect 15059 20244 15071 20247
rect 15102 20244 15108 20256
rect 15059 20216 15108 20244
rect 15059 20213 15071 20216
rect 15013 20207 15071 20213
rect 15102 20204 15108 20216
rect 15160 20204 15166 20256
rect 15838 20244 15844 20256
rect 15799 20216 15844 20244
rect 15838 20204 15844 20216
rect 15896 20204 15902 20256
rect 16025 20247 16083 20253
rect 16025 20213 16037 20247
rect 16071 20244 16083 20247
rect 17218 20244 17224 20256
rect 16071 20216 17224 20244
rect 16071 20213 16083 20216
rect 16025 20207 16083 20213
rect 17218 20204 17224 20216
rect 17276 20204 17282 20256
rect 18874 20244 18880 20256
rect 18835 20216 18880 20244
rect 18874 20204 18880 20216
rect 18932 20204 18938 20256
rect 18984 20244 19012 20352
rect 19334 20340 19340 20392
rect 19392 20380 19398 20392
rect 19613 20383 19671 20389
rect 19613 20380 19625 20383
rect 19392 20352 19625 20380
rect 19392 20340 19398 20352
rect 19613 20349 19625 20352
rect 19659 20349 19671 20383
rect 19613 20343 19671 20349
rect 25133 20383 25191 20389
rect 25133 20349 25145 20383
rect 25179 20349 25191 20383
rect 25240 20380 25268 20420
rect 26237 20417 26249 20420
rect 26283 20448 26295 20451
rect 26694 20448 26700 20460
rect 26283 20420 26700 20448
rect 26283 20417 26295 20420
rect 26237 20411 26295 20417
rect 26694 20408 26700 20420
rect 26752 20408 26758 20460
rect 27080 20380 27108 20479
rect 27614 20476 27620 20488
rect 27672 20476 27678 20528
rect 28736 20516 28764 20547
rect 29638 20544 29644 20596
rect 29696 20584 29702 20596
rect 30006 20584 30012 20596
rect 29696 20556 30012 20584
rect 29696 20544 29702 20556
rect 30006 20544 30012 20556
rect 30064 20544 30070 20596
rect 31570 20584 31576 20596
rect 31531 20556 31576 20584
rect 31570 20544 31576 20556
rect 31628 20544 31634 20596
rect 32122 20584 32128 20596
rect 32083 20556 32128 20584
rect 32122 20544 32128 20556
rect 32180 20544 32186 20596
rect 32214 20544 32220 20596
rect 32272 20584 32278 20596
rect 32493 20587 32551 20593
rect 32493 20584 32505 20587
rect 32272 20556 32505 20584
rect 32272 20544 32278 20556
rect 32493 20553 32505 20556
rect 32539 20553 32551 20587
rect 32493 20547 32551 20553
rect 33965 20587 34023 20593
rect 33965 20553 33977 20587
rect 34011 20584 34023 20587
rect 34882 20584 34888 20596
rect 34011 20556 34888 20584
rect 34011 20553 34023 20556
rect 33965 20547 34023 20553
rect 34882 20544 34888 20556
rect 34940 20544 34946 20596
rect 40221 20587 40279 20593
rect 34992 20556 38332 20584
rect 31846 20516 31852 20528
rect 28736 20488 30052 20516
rect 28166 20448 28172 20460
rect 28127 20420 28172 20448
rect 28166 20408 28172 20420
rect 28224 20408 28230 20460
rect 28537 20451 28595 20457
rect 28537 20417 28549 20451
rect 28583 20448 28595 20451
rect 28718 20448 28724 20460
rect 28583 20420 28724 20448
rect 28583 20417 28595 20420
rect 28537 20411 28595 20417
rect 25240 20352 27108 20380
rect 25133 20343 25191 20349
rect 24854 20272 24860 20324
rect 24912 20312 24918 20324
rect 25148 20312 25176 20343
rect 27246 20340 27252 20392
rect 27304 20380 27310 20392
rect 28552 20380 28580 20411
rect 28718 20408 28724 20420
rect 28776 20408 28782 20460
rect 29917 20451 29975 20457
rect 29917 20417 29929 20451
rect 29963 20417 29975 20451
rect 30024 20448 30052 20488
rect 30944 20488 31852 20516
rect 30944 20457 30972 20488
rect 31846 20476 31852 20488
rect 31904 20476 31910 20528
rect 33042 20516 33048 20528
rect 32324 20488 33048 20516
rect 30745 20451 30803 20457
rect 30745 20448 30757 20451
rect 30024 20420 30757 20448
rect 29917 20411 29975 20417
rect 27304 20352 28580 20380
rect 27304 20340 27310 20352
rect 25774 20312 25780 20324
rect 24912 20284 25780 20312
rect 24912 20272 24918 20284
rect 25774 20272 25780 20284
rect 25832 20312 25838 20324
rect 27433 20315 27491 20321
rect 27433 20312 27445 20315
rect 25832 20284 27445 20312
rect 25832 20272 25838 20284
rect 27433 20281 27445 20284
rect 27479 20312 27491 20315
rect 27890 20312 27896 20324
rect 27479 20284 27896 20312
rect 27479 20281 27491 20284
rect 27433 20275 27491 20281
rect 27890 20272 27896 20284
rect 27948 20272 27954 20324
rect 29932 20312 29960 20411
rect 30116 20389 30144 20420
rect 30745 20417 30757 20420
rect 30791 20417 30803 20451
rect 30745 20411 30803 20417
rect 30929 20451 30987 20457
rect 30929 20417 30941 20451
rect 30975 20417 30987 20451
rect 31386 20448 31392 20460
rect 31347 20420 31392 20448
rect 30929 20411 30987 20417
rect 31386 20408 31392 20420
rect 31444 20408 31450 20460
rect 32324 20457 32352 20488
rect 33042 20476 33048 20488
rect 33100 20476 33106 20528
rect 32309 20451 32367 20457
rect 32309 20417 32321 20451
rect 32355 20417 32367 20451
rect 32309 20411 32367 20417
rect 32582 20408 32588 20460
rect 32640 20448 32646 20460
rect 33873 20451 33931 20457
rect 32640 20420 32685 20448
rect 32640 20408 32646 20420
rect 33873 20417 33885 20451
rect 33919 20417 33931 20451
rect 34054 20448 34060 20460
rect 34015 20420 34060 20448
rect 33873 20411 33931 20417
rect 30101 20383 30159 20389
rect 30101 20349 30113 20383
rect 30147 20380 30159 20383
rect 30190 20380 30196 20392
rect 30147 20352 30196 20380
rect 30147 20349 30159 20352
rect 30101 20343 30159 20349
rect 30190 20340 30196 20352
rect 30248 20340 30254 20392
rect 30282 20340 30288 20392
rect 30340 20380 30346 20392
rect 33888 20380 33916 20411
rect 34054 20408 34060 20420
rect 34112 20408 34118 20460
rect 30340 20352 33916 20380
rect 30340 20340 30346 20352
rect 33870 20312 33876 20324
rect 29932 20284 33876 20312
rect 33870 20272 33876 20284
rect 33928 20272 33934 20324
rect 19978 20244 19984 20256
rect 18984 20216 19984 20244
rect 19978 20204 19984 20216
rect 20036 20204 20042 20256
rect 25222 20244 25228 20256
rect 25183 20216 25228 20244
rect 25222 20204 25228 20216
rect 25280 20204 25286 20256
rect 26326 20204 26332 20256
rect 26384 20244 26390 20256
rect 26421 20247 26479 20253
rect 26421 20244 26433 20247
rect 26384 20216 26433 20244
rect 26384 20204 26390 20216
rect 26421 20213 26433 20216
rect 26467 20244 26479 20247
rect 27154 20244 27160 20256
rect 26467 20216 27160 20244
rect 26467 20213 26479 20216
rect 26421 20207 26479 20213
rect 27154 20204 27160 20216
rect 27212 20204 27218 20256
rect 28534 20244 28540 20256
rect 28495 20216 28540 20244
rect 28534 20204 28540 20216
rect 28592 20204 28598 20256
rect 29546 20244 29552 20256
rect 29507 20216 29552 20244
rect 29546 20204 29552 20216
rect 29604 20204 29610 20256
rect 30374 20204 30380 20256
rect 30432 20244 30438 20256
rect 30745 20247 30803 20253
rect 30745 20244 30757 20247
rect 30432 20216 30757 20244
rect 30432 20204 30438 20216
rect 30745 20213 30757 20216
rect 30791 20213 30803 20247
rect 30745 20207 30803 20213
rect 32214 20204 32220 20256
rect 32272 20244 32278 20256
rect 34992 20244 35020 20556
rect 36262 20516 36268 20528
rect 36223 20488 36268 20516
rect 36262 20476 36268 20488
rect 36320 20476 36326 20528
rect 37182 20476 37188 20528
rect 37240 20516 37246 20528
rect 37240 20488 38240 20516
rect 37240 20476 37246 20488
rect 36170 20408 36176 20460
rect 36228 20448 36234 20460
rect 36906 20448 36912 20460
rect 36228 20420 36912 20448
rect 36228 20408 36234 20420
rect 36906 20408 36912 20420
rect 36964 20448 36970 20460
rect 37090 20448 37096 20460
rect 36964 20420 37096 20448
rect 36964 20408 36970 20420
rect 37090 20408 37096 20420
rect 37148 20448 37154 20460
rect 37737 20451 37795 20457
rect 37737 20448 37749 20451
rect 37148 20420 37749 20448
rect 37148 20408 37154 20420
rect 37737 20417 37749 20420
rect 37783 20417 37795 20451
rect 37737 20411 37795 20417
rect 37826 20408 37832 20460
rect 37884 20448 37890 20460
rect 38212 20457 38240 20488
rect 37921 20451 37979 20457
rect 37921 20448 37933 20451
rect 37884 20420 37933 20448
rect 37884 20408 37890 20420
rect 37921 20417 37933 20420
rect 37967 20417 37979 20451
rect 37921 20411 37979 20417
rect 38197 20451 38255 20457
rect 38197 20417 38209 20451
rect 38243 20417 38255 20451
rect 38304 20448 38332 20556
rect 40221 20553 40233 20587
rect 40267 20584 40279 20587
rect 40310 20584 40316 20596
rect 40267 20556 40316 20584
rect 40267 20553 40279 20556
rect 40221 20547 40279 20553
rect 40310 20544 40316 20556
rect 40368 20544 40374 20596
rect 38381 20519 38439 20525
rect 38381 20485 38393 20519
rect 38427 20516 38439 20519
rect 39086 20519 39144 20525
rect 39086 20516 39098 20519
rect 38427 20488 39098 20516
rect 38427 20485 38439 20488
rect 38381 20479 38439 20485
rect 39086 20485 39098 20488
rect 39132 20485 39144 20519
rect 39086 20479 39144 20485
rect 41386 20488 41644 20516
rect 40957 20451 41015 20457
rect 40957 20448 40969 20451
rect 38304 20420 40969 20448
rect 38197 20411 38255 20417
rect 40957 20417 40969 20420
rect 41003 20417 41015 20451
rect 40957 20411 41015 20417
rect 35894 20340 35900 20392
rect 35952 20380 35958 20392
rect 35952 20352 37504 20380
rect 35952 20340 35958 20352
rect 36170 20272 36176 20324
rect 36228 20312 36234 20324
rect 36633 20315 36691 20321
rect 36633 20312 36645 20315
rect 36228 20284 36645 20312
rect 36228 20272 36234 20284
rect 36633 20281 36645 20284
rect 36679 20281 36691 20315
rect 36633 20275 36691 20281
rect 32272 20216 35020 20244
rect 36725 20247 36783 20253
rect 32272 20204 32278 20216
rect 36725 20213 36737 20247
rect 36771 20244 36783 20247
rect 37274 20244 37280 20256
rect 36771 20216 37280 20244
rect 36771 20213 36783 20216
rect 36725 20207 36783 20213
rect 37274 20204 37280 20216
rect 37332 20204 37338 20256
rect 37476 20244 37504 20352
rect 37550 20340 37556 20392
rect 37608 20380 37614 20392
rect 38841 20383 38899 20389
rect 38841 20380 38853 20383
rect 37608 20352 38853 20380
rect 37608 20340 37614 20352
rect 38841 20349 38853 20352
rect 38887 20349 38899 20383
rect 38841 20343 38899 20349
rect 41386 20312 41414 20488
rect 41616 20457 41644 20488
rect 41601 20451 41659 20457
rect 41601 20417 41613 20451
rect 41647 20417 41659 20451
rect 41601 20411 41659 20417
rect 40144 20284 41414 20312
rect 40144 20244 40172 20284
rect 37476 20216 40172 20244
rect 40218 20204 40224 20256
rect 40276 20244 40282 20256
rect 41049 20247 41107 20253
rect 41049 20244 41061 20247
rect 40276 20216 41061 20244
rect 40276 20204 40282 20216
rect 41049 20213 41061 20216
rect 41095 20213 41107 20247
rect 41690 20244 41696 20256
rect 41651 20216 41696 20244
rect 41049 20207 41107 20213
rect 41690 20204 41696 20216
rect 41748 20204 41754 20256
rect 1104 20154 42872 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 42872 20154
rect 1104 20080 42872 20102
rect 5442 20000 5448 20052
rect 5500 20040 5506 20052
rect 39114 20040 39120 20052
rect 5500 20012 39120 20040
rect 5500 20000 5506 20012
rect 39114 20000 39120 20012
rect 39172 20040 39178 20052
rect 40862 20040 40868 20052
rect 39172 20012 40868 20040
rect 39172 20000 39178 20012
rect 40862 20000 40868 20012
rect 40920 20000 40926 20052
rect 16666 19932 16672 19984
rect 16724 19972 16730 19984
rect 17770 19972 17776 19984
rect 16724 19944 17776 19972
rect 16724 19932 16730 19944
rect 17770 19932 17776 19944
rect 17828 19972 17834 19984
rect 18417 19975 18475 19981
rect 18417 19972 18429 19975
rect 17828 19944 18429 19972
rect 17828 19932 17834 19944
rect 18417 19941 18429 19944
rect 18463 19972 18475 19975
rect 18782 19972 18788 19984
rect 18463 19944 18788 19972
rect 18463 19941 18475 19944
rect 18417 19935 18475 19941
rect 18782 19932 18788 19944
rect 18840 19972 18846 19984
rect 20714 19972 20720 19984
rect 18840 19944 19334 19972
rect 20675 19944 20720 19972
rect 18840 19932 18846 19944
rect 1394 19904 1400 19916
rect 1355 19876 1400 19904
rect 1394 19864 1400 19876
rect 1452 19864 1458 19916
rect 1854 19904 1860 19916
rect 1815 19876 1860 19904
rect 1854 19864 1860 19876
rect 1912 19864 1918 19916
rect 6730 19904 6736 19916
rect 6691 19876 6736 19904
rect 6730 19864 6736 19876
rect 6788 19864 6794 19916
rect 11606 19904 11612 19916
rect 11519 19876 11612 19904
rect 11606 19864 11612 19876
rect 11664 19904 11670 19916
rect 13354 19904 13360 19916
rect 11664 19876 13360 19904
rect 11664 19864 11670 19876
rect 13354 19864 13360 19876
rect 13412 19864 13418 19916
rect 15749 19907 15807 19913
rect 15749 19873 15761 19907
rect 15795 19904 15807 19907
rect 16574 19904 16580 19916
rect 15795 19876 16580 19904
rect 15795 19873 15807 19876
rect 15749 19867 15807 19873
rect 16574 19864 16580 19876
rect 16632 19864 16638 19916
rect 19306 19848 19334 19944
rect 20714 19932 20720 19944
rect 20772 19932 20778 19984
rect 24118 19932 24124 19984
rect 24176 19972 24182 19984
rect 24489 19975 24547 19981
rect 24489 19972 24501 19975
rect 24176 19944 24501 19972
rect 24176 19932 24182 19944
rect 24489 19941 24501 19944
rect 24535 19941 24547 19975
rect 26878 19972 26884 19984
rect 24489 19935 24547 19941
rect 24596 19944 26884 19972
rect 24596 19904 24624 19944
rect 26878 19932 26884 19944
rect 26936 19932 26942 19984
rect 28258 19972 28264 19984
rect 27080 19944 28264 19972
rect 23676 19876 24624 19904
rect 24857 19907 24915 19913
rect 6181 19839 6239 19845
rect 6181 19805 6193 19839
rect 6227 19836 6239 19839
rect 6362 19836 6368 19848
rect 6227 19808 6368 19836
rect 6227 19805 6239 19808
rect 6181 19799 6239 19805
rect 6362 19796 6368 19808
rect 6420 19796 6426 19848
rect 10318 19836 10324 19848
rect 10279 19808 10324 19836
rect 10318 19796 10324 19808
rect 10376 19796 10382 19848
rect 10505 19839 10563 19845
rect 10505 19805 10517 19839
rect 10551 19836 10563 19839
rect 11057 19839 11115 19845
rect 11057 19836 11069 19839
rect 10551 19808 11069 19836
rect 10551 19805 10563 19808
rect 10505 19799 10563 19805
rect 11057 19805 11069 19808
rect 11103 19836 11115 19839
rect 11238 19836 11244 19848
rect 11103 19808 11244 19836
rect 11103 19805 11115 19808
rect 11057 19799 11115 19805
rect 11238 19796 11244 19808
rect 11296 19796 11302 19848
rect 15838 19796 15844 19848
rect 15896 19836 15902 19848
rect 16022 19836 16028 19848
rect 15896 19808 16028 19836
rect 15896 19796 15902 19808
rect 16022 19796 16028 19808
rect 16080 19796 16086 19848
rect 19306 19836 19340 19848
rect 19247 19808 19340 19836
rect 19334 19796 19340 19808
rect 19392 19796 19398 19848
rect 21729 19839 21787 19845
rect 21729 19836 21741 19839
rect 19444 19808 21741 19836
rect 19444 19780 19472 19808
rect 21729 19805 21741 19808
rect 21775 19805 21787 19839
rect 21729 19799 21787 19805
rect 22373 19839 22431 19845
rect 22373 19805 22385 19839
rect 22419 19805 22431 19839
rect 22373 19799 22431 19805
rect 1581 19771 1639 19777
rect 1581 19737 1593 19771
rect 1627 19768 1639 19771
rect 2038 19768 2044 19780
rect 1627 19740 2044 19768
rect 1627 19737 1639 19740
rect 1581 19731 1639 19737
rect 2038 19728 2044 19740
rect 2096 19728 2102 19780
rect 18601 19771 18659 19777
rect 18601 19737 18613 19771
rect 18647 19768 18659 19771
rect 19426 19768 19432 19780
rect 18647 19740 19432 19768
rect 18647 19737 18659 19740
rect 18601 19731 18659 19737
rect 19426 19728 19432 19740
rect 19484 19728 19490 19780
rect 19604 19771 19662 19777
rect 19604 19737 19616 19771
rect 19650 19737 19662 19771
rect 19604 19731 19662 19737
rect 21913 19771 21971 19777
rect 21913 19737 21925 19771
rect 21959 19768 21971 19771
rect 22002 19768 22008 19780
rect 21959 19740 22008 19768
rect 21959 19737 21971 19740
rect 21913 19731 21971 19737
rect 2590 19660 2596 19712
rect 2648 19700 2654 19712
rect 11606 19700 11612 19712
rect 2648 19672 11612 19700
rect 2648 19660 2654 19672
rect 11606 19660 11612 19672
rect 11664 19660 11670 19712
rect 19334 19660 19340 19712
rect 19392 19700 19398 19712
rect 19628 19700 19656 19731
rect 22002 19728 22008 19740
rect 22060 19768 22066 19780
rect 22388 19768 22416 19799
rect 22060 19740 22416 19768
rect 22640 19771 22698 19777
rect 22060 19728 22066 19740
rect 22640 19737 22652 19771
rect 22686 19768 22698 19771
rect 22738 19768 22744 19780
rect 22686 19740 22744 19768
rect 22686 19737 22698 19740
rect 22640 19731 22698 19737
rect 22738 19728 22744 19740
rect 22796 19728 22802 19780
rect 19392 19672 19656 19700
rect 19392 19660 19398 19672
rect 21634 19660 21640 19712
rect 21692 19700 21698 19712
rect 23676 19700 23704 19876
rect 24857 19873 24869 19907
rect 24903 19904 24915 19907
rect 25498 19904 25504 19916
rect 24903 19876 25504 19904
rect 24903 19873 24915 19876
rect 24857 19867 24915 19873
rect 25498 19864 25504 19876
rect 25556 19864 25562 19916
rect 25774 19904 25780 19916
rect 25735 19876 25780 19904
rect 25774 19864 25780 19876
rect 25832 19864 25838 19916
rect 26326 19864 26332 19916
rect 26384 19904 26390 19916
rect 27080 19913 27108 19944
rect 28258 19932 28264 19944
rect 28316 19932 28322 19984
rect 30377 19975 30435 19981
rect 30377 19941 30389 19975
rect 30423 19972 30435 19975
rect 30650 19972 30656 19984
rect 30423 19944 30656 19972
rect 30423 19941 30435 19944
rect 30377 19935 30435 19941
rect 30650 19932 30656 19944
rect 30708 19932 30714 19984
rect 32493 19975 32551 19981
rect 32493 19941 32505 19975
rect 32539 19972 32551 19975
rect 32582 19972 32588 19984
rect 32539 19944 32588 19972
rect 32539 19941 32551 19944
rect 32493 19935 32551 19941
rect 32582 19932 32588 19944
rect 32640 19932 32646 19984
rect 37274 19932 37280 19984
rect 37332 19972 37338 19984
rect 37332 19944 38700 19972
rect 37332 19932 37338 19944
rect 27065 19907 27123 19913
rect 27065 19904 27077 19907
rect 26384 19876 27077 19904
rect 26384 19864 26390 19876
rect 27065 19873 27077 19876
rect 27111 19873 27123 19907
rect 27338 19904 27344 19916
rect 27299 19876 27344 19904
rect 27065 19867 27123 19873
rect 27338 19864 27344 19876
rect 27396 19904 27402 19916
rect 28077 19907 28135 19913
rect 27396 19876 27936 19904
rect 27396 19864 27402 19876
rect 24578 19796 24584 19848
rect 24636 19836 24642 19848
rect 24673 19839 24731 19845
rect 24673 19836 24685 19839
rect 24636 19808 24685 19836
rect 24636 19796 24642 19808
rect 24673 19805 24685 19808
rect 24719 19805 24731 19839
rect 24673 19799 24731 19805
rect 24762 19796 24768 19848
rect 24820 19836 24826 19848
rect 24820 19808 24865 19836
rect 24820 19796 24826 19808
rect 24946 19796 24952 19848
rect 25004 19836 25010 19848
rect 25004 19808 25049 19836
rect 25004 19796 25010 19808
rect 25222 19796 25228 19848
rect 25280 19836 25286 19848
rect 26973 19839 27031 19845
rect 26973 19836 26985 19839
rect 25280 19808 26985 19836
rect 25280 19796 25286 19808
rect 26973 19805 26985 19808
rect 27019 19836 27031 19839
rect 27246 19836 27252 19848
rect 27019 19808 27252 19836
rect 27019 19805 27031 19808
rect 26973 19799 27031 19805
rect 27246 19796 27252 19808
rect 27304 19796 27310 19848
rect 27908 19845 27936 19876
rect 28077 19873 28089 19907
rect 28123 19904 28135 19907
rect 28350 19904 28356 19916
rect 28123 19876 28356 19904
rect 28123 19873 28135 19876
rect 28077 19867 28135 19873
rect 28350 19864 28356 19876
rect 28408 19904 28414 19916
rect 34698 19904 34704 19916
rect 28408 19876 34704 19904
rect 28408 19864 28414 19876
rect 34698 19864 34704 19876
rect 34756 19904 34762 19916
rect 34793 19907 34851 19913
rect 34793 19904 34805 19907
rect 34756 19876 34805 19904
rect 34756 19864 34762 19876
rect 34793 19873 34805 19876
rect 34839 19873 34851 19907
rect 34793 19867 34851 19873
rect 36899 19907 36957 19913
rect 36899 19873 36911 19907
rect 36945 19904 36957 19907
rect 37090 19904 37096 19916
rect 36945 19876 37096 19904
rect 36945 19873 36957 19876
rect 36899 19867 36957 19873
rect 37090 19864 37096 19876
rect 37148 19864 37154 19916
rect 38565 19907 38623 19913
rect 38565 19904 38577 19907
rect 37936 19876 38577 19904
rect 37936 19848 37964 19876
rect 38565 19873 38577 19876
rect 38611 19873 38623 19907
rect 38565 19867 38623 19873
rect 27893 19839 27951 19845
rect 27893 19805 27905 19839
rect 27939 19805 27951 19839
rect 30098 19836 30104 19848
rect 30059 19808 30104 19836
rect 27893 19799 27951 19805
rect 30098 19796 30104 19808
rect 30156 19796 30162 19848
rect 30190 19796 30196 19848
rect 30248 19836 30254 19848
rect 30374 19836 30380 19848
rect 30248 19808 30293 19836
rect 30335 19808 30380 19836
rect 30248 19796 30254 19808
rect 30374 19796 30380 19808
rect 30432 19796 30438 19848
rect 32309 19839 32367 19845
rect 32309 19805 32321 19839
rect 32355 19836 32367 19839
rect 32398 19836 32404 19848
rect 32355 19808 32404 19836
rect 32355 19805 32367 19808
rect 32309 19799 32367 19805
rect 32398 19796 32404 19808
rect 32456 19796 32462 19848
rect 32585 19839 32643 19845
rect 32585 19805 32597 19839
rect 32631 19836 32643 19839
rect 33594 19836 33600 19848
rect 32631 19808 33600 19836
rect 32631 19805 32643 19808
rect 32585 19799 32643 19805
rect 33594 19796 33600 19808
rect 33652 19836 33658 19848
rect 34885 19839 34943 19845
rect 34885 19836 34897 19839
rect 33652 19808 34897 19836
rect 33652 19796 33658 19808
rect 34885 19805 34897 19808
rect 34931 19805 34943 19839
rect 36814 19836 36820 19848
rect 36775 19808 36820 19836
rect 34885 19799 34943 19805
rect 36814 19796 36820 19808
rect 36872 19796 36878 19848
rect 37001 19839 37059 19845
rect 37001 19805 37013 19839
rect 37047 19836 37059 19839
rect 37182 19836 37188 19848
rect 37047 19808 37188 19836
rect 37047 19805 37059 19808
rect 37001 19799 37059 19805
rect 37182 19796 37188 19808
rect 37240 19836 37246 19848
rect 37553 19839 37611 19845
rect 37553 19836 37565 19839
rect 37240 19808 37565 19836
rect 37240 19796 37246 19808
rect 37553 19805 37565 19808
rect 37599 19805 37611 19839
rect 37553 19799 37611 19805
rect 37829 19839 37887 19845
rect 37829 19805 37841 19839
rect 37875 19836 37887 19839
rect 37918 19836 37924 19848
rect 37875 19808 37924 19836
rect 37875 19805 37887 19808
rect 37829 19799 37887 19805
rect 37918 19796 37924 19808
rect 37976 19796 37982 19848
rect 38470 19836 38476 19848
rect 38431 19808 38476 19836
rect 38470 19796 38476 19808
rect 38528 19796 38534 19848
rect 38672 19845 38700 19944
rect 39132 19845 39160 20000
rect 40497 19907 40555 19913
rect 40497 19873 40509 19907
rect 40543 19904 40555 19907
rect 41690 19904 41696 19916
rect 40543 19876 41696 19904
rect 40543 19873 40555 19876
rect 40497 19867 40555 19873
rect 41690 19864 41696 19876
rect 41748 19864 41754 19916
rect 38657 19839 38715 19845
rect 38657 19805 38669 19839
rect 38703 19805 38715 19839
rect 38657 19799 38715 19805
rect 39117 19839 39175 19845
rect 39117 19805 39129 19839
rect 39163 19805 39175 19839
rect 40310 19836 40316 19848
rect 40271 19808 40316 19836
rect 39117 19799 39175 19805
rect 40310 19796 40316 19808
rect 40368 19796 40374 19848
rect 23934 19728 23940 19780
rect 23992 19768 23998 19780
rect 35894 19768 35900 19780
rect 23992 19740 35900 19768
rect 23992 19728 23998 19740
rect 35894 19728 35900 19740
rect 35952 19728 35958 19780
rect 37090 19728 37096 19780
rect 37148 19768 37154 19780
rect 37645 19771 37703 19777
rect 37645 19768 37657 19771
rect 37148 19740 37657 19768
rect 37148 19728 37154 19740
rect 37645 19737 37657 19740
rect 37691 19737 37703 19771
rect 42150 19768 42156 19780
rect 42111 19740 42156 19768
rect 37645 19731 37703 19737
rect 42150 19728 42156 19740
rect 42208 19728 42214 19780
rect 21692 19672 23704 19700
rect 23753 19703 23811 19709
rect 21692 19660 21698 19672
rect 23753 19669 23765 19703
rect 23799 19700 23811 19703
rect 24578 19700 24584 19712
rect 23799 19672 24584 19700
rect 23799 19669 23811 19672
rect 23753 19663 23811 19669
rect 24578 19660 24584 19672
rect 24636 19660 24642 19712
rect 32125 19703 32183 19709
rect 32125 19669 32137 19703
rect 32171 19700 32183 19703
rect 32490 19700 32496 19712
rect 32171 19672 32496 19700
rect 32171 19669 32183 19672
rect 32125 19663 32183 19669
rect 32490 19660 32496 19672
rect 32548 19660 32554 19712
rect 34974 19660 34980 19712
rect 35032 19700 35038 19712
rect 35253 19703 35311 19709
rect 35253 19700 35265 19703
rect 35032 19672 35265 19700
rect 35032 19660 35038 19672
rect 35253 19669 35265 19672
rect 35299 19669 35311 19703
rect 36630 19700 36636 19712
rect 36591 19672 36636 19700
rect 35253 19663 35311 19669
rect 36630 19660 36636 19672
rect 36688 19660 36694 19712
rect 38010 19700 38016 19712
rect 37971 19672 38016 19700
rect 38010 19660 38016 19672
rect 38068 19660 38074 19712
rect 39209 19703 39267 19709
rect 39209 19669 39221 19703
rect 39255 19700 39267 19703
rect 40402 19700 40408 19712
rect 39255 19672 40408 19700
rect 39255 19669 39267 19672
rect 39209 19663 39267 19669
rect 40402 19660 40408 19672
rect 40460 19660 40466 19712
rect 1104 19610 42872 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 42872 19610
rect 1104 19536 42872 19558
rect 2038 19496 2044 19508
rect 1999 19468 2044 19496
rect 2038 19456 2044 19468
rect 2096 19456 2102 19508
rect 8938 19456 8944 19508
rect 8996 19496 9002 19508
rect 16206 19496 16212 19508
rect 8996 19468 12020 19496
rect 8996 19456 9002 19468
rect 11992 19437 12020 19468
rect 15856 19468 16212 19496
rect 11977 19431 12035 19437
rect 10520 19400 11284 19428
rect 2130 19360 2136 19372
rect 2091 19332 2136 19360
rect 2130 19320 2136 19332
rect 2188 19320 2194 19372
rect 10520 19369 10548 19400
rect 11256 19372 11284 19400
rect 11977 19397 11989 19431
rect 12023 19428 12035 19431
rect 12158 19428 12164 19440
rect 12023 19400 12164 19428
rect 12023 19397 12035 19400
rect 11977 19391 12035 19397
rect 12158 19388 12164 19400
rect 12216 19388 12222 19440
rect 15010 19388 15016 19440
rect 15068 19428 15074 19440
rect 15856 19437 15884 19468
rect 16206 19456 16212 19468
rect 16264 19456 16270 19508
rect 19334 19456 19340 19508
rect 19392 19496 19398 19508
rect 19613 19499 19671 19505
rect 19613 19496 19625 19499
rect 19392 19468 19625 19496
rect 19392 19456 19398 19468
rect 19613 19465 19625 19468
rect 19659 19465 19671 19499
rect 19613 19459 19671 19465
rect 23753 19499 23811 19505
rect 23753 19465 23765 19499
rect 23799 19465 23811 19499
rect 24302 19496 24308 19508
rect 24263 19468 24308 19496
rect 23753 19459 23811 19465
rect 15749 19431 15807 19437
rect 15749 19428 15761 19431
rect 15068 19400 15761 19428
rect 15068 19388 15074 19400
rect 15749 19397 15761 19400
rect 15795 19397 15807 19431
rect 15749 19391 15807 19397
rect 15841 19431 15899 19437
rect 15841 19397 15853 19431
rect 15887 19397 15899 19431
rect 15841 19391 15899 19397
rect 15979 19431 16037 19437
rect 15979 19397 15991 19431
rect 16025 19428 16037 19431
rect 16298 19428 16304 19440
rect 16025 19400 16304 19428
rect 16025 19397 16037 19400
rect 15979 19391 16037 19397
rect 16298 19388 16304 19400
rect 16356 19388 16362 19440
rect 10505 19363 10563 19369
rect 10505 19329 10517 19363
rect 10551 19329 10563 19363
rect 10505 19323 10563 19329
rect 10686 19320 10692 19372
rect 10744 19360 10750 19372
rect 10781 19363 10839 19369
rect 10781 19360 10793 19363
rect 10744 19332 10793 19360
rect 10744 19320 10750 19332
rect 10781 19329 10793 19332
rect 10827 19329 10839 19363
rect 10781 19323 10839 19329
rect 11238 19320 11244 19372
rect 11296 19360 11302 19372
rect 11609 19363 11667 19369
rect 11609 19360 11621 19363
rect 11296 19332 11621 19360
rect 11296 19320 11302 19332
rect 11609 19329 11621 19332
rect 11655 19329 11667 19363
rect 12894 19360 12900 19372
rect 12855 19332 12900 19360
rect 11609 19323 11667 19329
rect 12894 19320 12900 19332
rect 12952 19320 12958 19372
rect 13164 19363 13222 19369
rect 13164 19329 13176 19363
rect 13210 19360 13222 19363
rect 15473 19363 15531 19369
rect 15473 19360 15485 19363
rect 13210 19332 15485 19360
rect 13210 19329 13222 19332
rect 13164 19323 13222 19329
rect 15473 19329 15485 19332
rect 15519 19329 15531 19363
rect 15654 19360 15660 19372
rect 15615 19332 15660 19360
rect 15473 19323 15531 19329
rect 15654 19320 15660 19332
rect 15712 19320 15718 19372
rect 16114 19360 16120 19372
rect 16075 19332 16120 19360
rect 16114 19320 16120 19332
rect 16172 19320 16178 19372
rect 16853 19363 16911 19369
rect 16853 19360 16865 19363
rect 16500 19332 16865 19360
rect 15838 19252 15844 19304
rect 15896 19292 15902 19304
rect 16500 19292 16528 19332
rect 16853 19329 16865 19332
rect 16899 19329 16911 19363
rect 16853 19323 16911 19329
rect 17770 19320 17776 19372
rect 17828 19369 17834 19372
rect 18046 19369 18052 19372
rect 17828 19360 17838 19369
rect 17828 19332 17873 19360
rect 17828 19323 17838 19332
rect 18040 19323 18052 19369
rect 18104 19360 18110 19372
rect 18104 19332 18140 19360
rect 17828 19320 17834 19323
rect 18046 19320 18052 19323
rect 18104 19320 18110 19332
rect 18874 19320 18880 19372
rect 18932 19360 18938 19372
rect 19797 19363 19855 19369
rect 19797 19360 19809 19363
rect 18932 19332 19809 19360
rect 18932 19320 18938 19332
rect 19797 19329 19809 19332
rect 19843 19329 19855 19363
rect 19797 19323 19855 19329
rect 22002 19320 22008 19372
rect 22060 19360 22066 19372
rect 22373 19363 22431 19369
rect 22373 19360 22385 19363
rect 22060 19332 22385 19360
rect 22060 19320 22066 19332
rect 22373 19329 22385 19332
rect 22419 19329 22431 19363
rect 22373 19323 22431 19329
rect 22462 19320 22468 19372
rect 22520 19360 22526 19372
rect 22629 19363 22687 19369
rect 22629 19360 22641 19363
rect 22520 19332 22641 19360
rect 22520 19320 22526 19332
rect 22629 19329 22641 19332
rect 22675 19329 22687 19363
rect 23768 19360 23796 19459
rect 24302 19456 24308 19468
rect 24360 19456 24366 19508
rect 24946 19496 24952 19508
rect 24412 19468 24952 19496
rect 24412 19428 24440 19468
rect 24946 19456 24952 19468
rect 25004 19456 25010 19508
rect 25222 19496 25228 19508
rect 25183 19468 25228 19496
rect 25222 19456 25228 19468
rect 25280 19456 25286 19508
rect 27062 19496 27068 19508
rect 27023 19468 27068 19496
rect 27062 19456 27068 19468
rect 27120 19456 27126 19508
rect 32398 19496 32404 19508
rect 32359 19468 32404 19496
rect 32398 19456 32404 19468
rect 32456 19456 32462 19508
rect 37182 19456 37188 19508
rect 37240 19496 37246 19508
rect 37645 19499 37703 19505
rect 37645 19496 37657 19499
rect 37240 19468 37657 19496
rect 37240 19456 37246 19468
rect 37645 19465 37657 19468
rect 37691 19465 37703 19499
rect 37645 19459 37703 19465
rect 24228 19400 24440 19428
rect 24228 19369 24256 19400
rect 26878 19388 26884 19440
rect 26936 19428 26942 19440
rect 32214 19428 32220 19440
rect 26936 19400 32220 19428
rect 26936 19388 26942 19400
rect 32214 19388 32220 19400
rect 32272 19388 32278 19440
rect 32493 19431 32551 19437
rect 32493 19397 32505 19431
rect 32539 19428 32551 19431
rect 33594 19428 33600 19440
rect 32539 19400 33600 19428
rect 32539 19397 32551 19400
rect 32493 19391 32551 19397
rect 33594 19388 33600 19400
rect 33652 19388 33658 19440
rect 40218 19428 40224 19440
rect 40179 19400 40224 19428
rect 40218 19388 40224 19400
rect 40276 19388 40282 19440
rect 24213 19363 24271 19369
rect 24213 19360 24225 19363
rect 23768 19332 24225 19360
rect 22629 19323 22687 19329
rect 24213 19329 24225 19332
rect 24259 19329 24271 19363
rect 24213 19323 24271 19329
rect 24486 19320 24492 19372
rect 24544 19360 24550 19372
rect 24762 19360 24768 19372
rect 24544 19332 24768 19360
rect 24544 19320 24550 19332
rect 24762 19320 24768 19332
rect 24820 19360 24826 19372
rect 25133 19363 25191 19369
rect 25133 19360 25145 19363
rect 24820 19332 25145 19360
rect 24820 19320 24826 19332
rect 25133 19329 25145 19332
rect 25179 19329 25191 19363
rect 25133 19323 25191 19329
rect 25498 19320 25504 19372
rect 25556 19360 25562 19372
rect 25777 19363 25835 19369
rect 25777 19360 25789 19363
rect 25556 19332 25789 19360
rect 25556 19320 25562 19332
rect 25777 19329 25789 19332
rect 25823 19329 25835 19363
rect 25961 19363 26019 19369
rect 25961 19360 25973 19363
rect 25777 19323 25835 19329
rect 25884 19332 25973 19360
rect 15896 19264 16528 19292
rect 16669 19295 16727 19301
rect 15896 19252 15902 19264
rect 16669 19261 16681 19295
rect 16715 19292 16727 19295
rect 24578 19292 24584 19304
rect 16715 19264 17172 19292
rect 24539 19264 24584 19292
rect 16715 19261 16727 19264
rect 16669 19255 16727 19261
rect 14274 19156 14280 19168
rect 14235 19128 14280 19156
rect 14274 19116 14280 19128
rect 14332 19116 14338 19168
rect 16942 19116 16948 19168
rect 17000 19156 17006 19168
rect 17037 19159 17095 19165
rect 17037 19156 17049 19159
rect 17000 19128 17049 19156
rect 17000 19116 17006 19128
rect 17037 19125 17049 19128
rect 17083 19125 17095 19159
rect 17144 19156 17172 19264
rect 24578 19252 24584 19264
rect 24636 19292 24642 19304
rect 25884 19292 25912 19332
rect 25961 19329 25973 19332
rect 26007 19329 26019 19363
rect 25961 19323 26019 19329
rect 27157 19363 27215 19369
rect 27157 19329 27169 19363
rect 27203 19360 27215 19363
rect 27338 19360 27344 19372
rect 27203 19332 27344 19360
rect 27203 19329 27215 19332
rect 27157 19323 27215 19329
rect 27338 19320 27344 19332
rect 27396 19320 27402 19372
rect 28718 19360 28724 19372
rect 28679 19332 28724 19360
rect 28718 19320 28724 19332
rect 28776 19320 28782 19372
rect 29181 19363 29239 19369
rect 29181 19329 29193 19363
rect 29227 19360 29239 19363
rect 29546 19360 29552 19372
rect 29227 19332 29552 19360
rect 29227 19329 29239 19332
rect 29181 19323 29239 19329
rect 29546 19320 29552 19332
rect 29604 19360 29610 19372
rect 29825 19363 29883 19369
rect 29825 19360 29837 19363
rect 29604 19332 29837 19360
rect 29604 19320 29610 19332
rect 29825 19329 29837 19332
rect 29871 19360 29883 19363
rect 29914 19360 29920 19372
rect 29871 19332 29920 19360
rect 29871 19329 29883 19332
rect 29825 19323 29883 19329
rect 29914 19320 29920 19332
rect 29972 19320 29978 19372
rect 30009 19363 30067 19369
rect 30009 19329 30021 19363
rect 30055 19360 30067 19363
rect 30466 19360 30472 19372
rect 30055 19332 30472 19360
rect 30055 19329 30067 19332
rect 30009 19323 30067 19329
rect 24636 19264 25912 19292
rect 28905 19295 28963 19301
rect 24636 19252 24642 19264
rect 28905 19261 28917 19295
rect 28951 19292 28963 19295
rect 30024 19292 30052 19323
rect 30466 19320 30472 19332
rect 30524 19320 30530 19372
rect 32582 19360 32588 19372
rect 32543 19332 32588 19360
rect 32582 19320 32588 19332
rect 32640 19320 32646 19372
rect 34885 19363 34943 19369
rect 34885 19329 34897 19363
rect 34931 19360 34943 19363
rect 35342 19360 35348 19372
rect 34931 19332 35348 19360
rect 34931 19329 34943 19332
rect 34885 19323 34943 19329
rect 35342 19320 35348 19332
rect 35400 19320 35406 19372
rect 37461 19363 37519 19369
rect 37461 19329 37473 19363
rect 37507 19360 37519 19363
rect 38470 19360 38476 19372
rect 37507 19332 38476 19360
rect 37507 19329 37519 19332
rect 37461 19323 37519 19329
rect 28951 19264 30052 19292
rect 28951 19261 28963 19264
rect 28905 19255 28963 19261
rect 30098 19252 30104 19304
rect 30156 19292 30162 19304
rect 32122 19292 32128 19304
rect 30156 19264 30201 19292
rect 32083 19264 32128 19292
rect 30156 19252 30162 19264
rect 32122 19252 32128 19264
rect 32180 19252 32186 19304
rect 34974 19292 34980 19304
rect 34935 19264 34980 19292
rect 34974 19252 34980 19264
rect 35032 19252 35038 19304
rect 37476 19292 37504 19323
rect 38470 19320 38476 19332
rect 38528 19320 38534 19372
rect 40034 19360 40040 19372
rect 39995 19332 40040 19360
rect 40034 19320 40040 19332
rect 40092 19320 40098 19372
rect 41230 19292 41236 19304
rect 35268 19264 37504 19292
rect 41191 19264 41236 19292
rect 24302 19184 24308 19236
rect 24360 19224 24366 19236
rect 24670 19224 24676 19236
rect 24360 19196 24676 19224
rect 24360 19184 24366 19196
rect 24670 19184 24676 19196
rect 24728 19184 24734 19236
rect 25777 19227 25835 19233
rect 25777 19193 25789 19227
rect 25823 19224 25835 19227
rect 26326 19224 26332 19236
rect 25823 19196 26332 19224
rect 25823 19193 25835 19196
rect 25777 19187 25835 19193
rect 26326 19184 26332 19196
rect 26384 19184 26390 19236
rect 28994 19224 29000 19236
rect 28953 19196 29000 19224
rect 28994 19184 29000 19196
rect 29052 19233 29058 19236
rect 29052 19227 29101 19233
rect 29052 19193 29055 19227
rect 29089 19224 29101 19227
rect 30116 19224 30144 19252
rect 35268 19233 35296 19264
rect 41230 19252 41236 19264
rect 41288 19252 41294 19304
rect 29089 19196 30144 19224
rect 35253 19227 35311 19233
rect 29089 19193 29101 19196
rect 29052 19187 29101 19193
rect 35253 19193 35265 19227
rect 35299 19193 35311 19227
rect 35253 19187 35311 19193
rect 39577 19227 39635 19233
rect 39577 19193 39589 19227
rect 39623 19224 39635 19227
rect 40310 19224 40316 19236
rect 39623 19196 40316 19224
rect 39623 19193 39635 19196
rect 39577 19187 39635 19193
rect 29052 19184 29058 19187
rect 40310 19184 40316 19196
rect 40368 19184 40374 19236
rect 18690 19156 18696 19168
rect 17144 19128 18696 19156
rect 17037 19119 17095 19125
rect 18690 19116 18696 19128
rect 18748 19156 18754 19168
rect 19153 19159 19211 19165
rect 19153 19156 19165 19159
rect 18748 19128 19165 19156
rect 18748 19116 18754 19128
rect 19153 19125 19165 19128
rect 19199 19125 19211 19159
rect 19153 19119 19211 19125
rect 24397 19159 24455 19165
rect 24397 19125 24409 19159
rect 24443 19156 24455 19159
rect 24854 19156 24860 19168
rect 24443 19128 24860 19156
rect 24443 19125 24455 19128
rect 24397 19119 24455 19125
rect 24854 19116 24860 19128
rect 24912 19116 24918 19168
rect 28810 19156 28816 19168
rect 28771 19128 28816 19156
rect 28810 19116 28816 19128
rect 28868 19116 28874 19168
rect 29641 19159 29699 19165
rect 29641 19125 29653 19159
rect 29687 19156 29699 19159
rect 29822 19156 29828 19168
rect 29687 19128 29828 19156
rect 29687 19125 29699 19128
rect 29641 19119 29699 19125
rect 29822 19116 29828 19128
rect 29880 19116 29886 19168
rect 1104 19066 42872 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 42872 19066
rect 1104 18992 42872 19014
rect 17957 18955 18015 18961
rect 17957 18921 17969 18955
rect 18003 18952 18015 18955
rect 18046 18952 18052 18964
rect 18003 18924 18052 18952
rect 18003 18921 18015 18924
rect 17957 18915 18015 18921
rect 18046 18912 18052 18924
rect 18104 18912 18110 18964
rect 19426 18912 19432 18964
rect 19484 18952 19490 18964
rect 20257 18955 20315 18961
rect 20257 18952 20269 18955
rect 19484 18924 20269 18952
rect 19484 18912 19490 18924
rect 20257 18921 20269 18924
rect 20303 18921 20315 18955
rect 20257 18915 20315 18921
rect 20806 18912 20812 18964
rect 20864 18952 20870 18964
rect 26234 18952 26240 18964
rect 20864 18924 26240 18952
rect 20864 18912 20870 18924
rect 26234 18912 26240 18924
rect 26292 18912 26298 18964
rect 33594 18952 33600 18964
rect 33555 18924 33600 18952
rect 33594 18912 33600 18924
rect 33652 18912 33658 18964
rect 13541 18887 13599 18893
rect 13541 18853 13553 18887
rect 13587 18884 13599 18887
rect 14642 18884 14648 18896
rect 13587 18856 14648 18884
rect 13587 18853 13599 18856
rect 13541 18847 13599 18853
rect 14642 18844 14648 18856
rect 14700 18884 14706 18896
rect 15010 18884 15016 18896
rect 14700 18856 15016 18884
rect 14700 18844 14706 18856
rect 15010 18844 15016 18856
rect 15068 18844 15074 18896
rect 19613 18887 19671 18893
rect 19613 18853 19625 18887
rect 19659 18884 19671 18887
rect 20070 18884 20076 18896
rect 19659 18856 20076 18884
rect 19659 18853 19671 18856
rect 19613 18847 19671 18853
rect 20070 18844 20076 18856
rect 20128 18844 20134 18896
rect 22738 18884 22744 18896
rect 22699 18856 22744 18884
rect 22738 18844 22744 18856
rect 22796 18844 22802 18896
rect 25498 18844 25504 18896
rect 25556 18884 25562 18896
rect 25777 18887 25835 18893
rect 25777 18884 25789 18887
rect 25556 18856 25789 18884
rect 25556 18844 25562 18856
rect 25777 18853 25789 18856
rect 25823 18853 25835 18887
rect 25777 18847 25835 18853
rect 14274 18776 14280 18828
rect 14332 18816 14338 18828
rect 14553 18819 14611 18825
rect 14553 18816 14565 18819
rect 14332 18788 14565 18816
rect 14332 18776 14338 18788
rect 14553 18785 14565 18788
rect 14599 18816 14611 18819
rect 14918 18816 14924 18828
rect 14599 18788 14924 18816
rect 14599 18785 14611 18788
rect 14553 18779 14611 18785
rect 14918 18776 14924 18788
rect 14976 18816 14982 18828
rect 15381 18819 15439 18825
rect 15381 18816 15393 18819
rect 14976 18788 15393 18816
rect 14976 18776 14982 18788
rect 15381 18785 15393 18788
rect 15427 18785 15439 18819
rect 15381 18779 15439 18785
rect 15657 18819 15715 18825
rect 15657 18785 15669 18819
rect 15703 18816 15715 18819
rect 16114 18816 16120 18828
rect 15703 18788 16120 18816
rect 15703 18785 15715 18788
rect 15657 18779 15715 18785
rect 16114 18776 16120 18788
rect 16172 18776 16178 18828
rect 16298 18776 16304 18828
rect 16356 18816 16362 18828
rect 24397 18819 24455 18825
rect 24397 18816 24409 18819
rect 16356 18788 17816 18816
rect 16356 18776 16362 18788
rect 11057 18751 11115 18757
rect 11057 18717 11069 18751
rect 11103 18748 11115 18751
rect 11238 18748 11244 18760
rect 11103 18720 11244 18748
rect 11103 18717 11115 18720
rect 11057 18711 11115 18717
rect 11238 18708 11244 18720
rect 11296 18708 11302 18760
rect 14737 18751 14795 18757
rect 14737 18717 14749 18751
rect 14783 18748 14795 18751
rect 15010 18748 15016 18760
rect 14783 18720 15016 18748
rect 14783 18717 14795 18720
rect 14737 18711 14795 18717
rect 15010 18708 15016 18720
rect 15068 18708 15074 18760
rect 16942 18748 16948 18760
rect 16903 18720 16948 18748
rect 16942 18708 16948 18720
rect 17000 18708 17006 18760
rect 17402 18748 17408 18760
rect 17363 18720 17408 18748
rect 17402 18708 17408 18720
rect 17460 18708 17466 18760
rect 17788 18757 17816 18788
rect 22066 18788 24409 18816
rect 22066 18760 22094 18788
rect 24397 18785 24409 18788
rect 24443 18785 24455 18819
rect 24397 18779 24455 18785
rect 28810 18776 28816 18828
rect 28868 18816 28874 18828
rect 29733 18819 29791 18825
rect 29733 18816 29745 18819
rect 28868 18788 29745 18816
rect 28868 18776 28874 18788
rect 29733 18785 29745 18788
rect 29779 18785 29791 18819
rect 29733 18779 29791 18785
rect 30006 18776 30012 18828
rect 30064 18816 30070 18828
rect 30193 18819 30251 18825
rect 30193 18816 30205 18819
rect 30064 18788 30205 18816
rect 30064 18776 30070 18788
rect 30193 18785 30205 18788
rect 30239 18785 30251 18819
rect 40402 18816 40408 18828
rect 40363 18788 40408 18816
rect 30193 18779 30251 18785
rect 40402 18776 40408 18788
rect 40460 18776 40466 18828
rect 17773 18751 17831 18757
rect 17773 18717 17785 18751
rect 17819 18717 17831 18751
rect 20898 18748 20904 18760
rect 20859 18720 20904 18748
rect 17773 18711 17831 18717
rect 20898 18708 20904 18720
rect 20956 18748 20962 18760
rect 22002 18748 22008 18760
rect 20956 18720 22008 18748
rect 20956 18708 20962 18720
rect 22002 18708 22008 18720
rect 22060 18720 22094 18760
rect 22060 18708 22066 18720
rect 22278 18708 22284 18760
rect 22336 18748 22342 18760
rect 22925 18751 22983 18757
rect 22925 18748 22937 18751
rect 22336 18720 22937 18748
rect 22336 18708 22342 18720
rect 22925 18717 22937 18720
rect 22971 18717 22983 18751
rect 22925 18711 22983 18717
rect 28629 18751 28687 18757
rect 28629 18717 28641 18751
rect 28675 18748 28687 18751
rect 28994 18748 29000 18760
rect 28675 18720 29000 18748
rect 28675 18717 28687 18720
rect 28629 18711 28687 18717
rect 28994 18708 29000 18720
rect 29052 18708 29058 18760
rect 29822 18708 29828 18760
rect 29880 18748 29886 18760
rect 29880 18720 29925 18748
rect 29880 18708 29886 18720
rect 30466 18708 30472 18760
rect 30524 18748 30530 18760
rect 30653 18751 30711 18757
rect 30653 18748 30665 18751
rect 30524 18720 30665 18748
rect 30524 18708 30530 18720
rect 30653 18717 30665 18720
rect 30699 18717 30711 18751
rect 30653 18711 30711 18717
rect 30837 18751 30895 18757
rect 30837 18717 30849 18751
rect 30883 18717 30895 18751
rect 30837 18711 30895 18717
rect 32217 18751 32275 18757
rect 32217 18717 32229 18751
rect 32263 18748 32275 18751
rect 32306 18748 32312 18760
rect 32263 18720 32312 18748
rect 32263 18717 32275 18720
rect 32217 18711 32275 18717
rect 11609 18683 11667 18689
rect 11609 18649 11621 18683
rect 11655 18680 11667 18683
rect 11698 18680 11704 18692
rect 11655 18652 11704 18680
rect 11655 18649 11667 18652
rect 11609 18643 11667 18649
rect 11698 18640 11704 18652
rect 11756 18640 11762 18692
rect 13357 18683 13415 18689
rect 13357 18649 13369 18683
rect 13403 18680 13415 18683
rect 13630 18680 13636 18692
rect 13403 18652 13636 18680
rect 13403 18649 13415 18652
rect 13357 18643 13415 18649
rect 13630 18640 13636 18652
rect 13688 18640 13694 18692
rect 16666 18680 16672 18692
rect 16627 18652 16672 18680
rect 16666 18640 16672 18652
rect 16724 18640 16730 18692
rect 17586 18680 17592 18692
rect 17547 18652 17592 18680
rect 17586 18640 17592 18652
rect 17644 18640 17650 18692
rect 17681 18683 17739 18689
rect 17681 18649 17693 18683
rect 17727 18680 17739 18683
rect 18874 18680 18880 18692
rect 17727 18652 18880 18680
rect 17727 18649 17739 18652
rect 17681 18643 17739 18649
rect 18874 18640 18880 18652
rect 18932 18680 18938 18692
rect 19245 18683 19303 18689
rect 19245 18680 19257 18683
rect 18932 18652 19257 18680
rect 18932 18640 18938 18652
rect 19245 18649 19257 18652
rect 19291 18649 19303 18683
rect 19245 18643 19303 18649
rect 20349 18683 20407 18689
rect 20349 18649 20361 18683
rect 20395 18680 20407 18683
rect 20806 18680 20812 18692
rect 20395 18652 20812 18680
rect 20395 18649 20407 18652
rect 20349 18643 20407 18649
rect 20806 18640 20812 18652
rect 20864 18640 20870 18692
rect 20990 18640 20996 18692
rect 21048 18680 21054 18692
rect 21146 18683 21204 18689
rect 21146 18680 21158 18683
rect 21048 18652 21158 18680
rect 21048 18640 21054 18652
rect 21146 18649 21158 18652
rect 21192 18649 21204 18683
rect 21146 18643 21204 18649
rect 23566 18640 23572 18692
rect 23624 18680 23630 18692
rect 24642 18683 24700 18689
rect 24642 18680 24654 18683
rect 23624 18652 24654 18680
rect 23624 18640 23630 18652
rect 24642 18649 24654 18652
rect 24688 18649 24700 18683
rect 24642 18643 24700 18649
rect 28813 18683 28871 18689
rect 28813 18649 28825 18683
rect 28859 18680 28871 18683
rect 29914 18680 29920 18692
rect 28859 18652 29920 18680
rect 28859 18649 28871 18652
rect 28813 18643 28871 18649
rect 29914 18640 29920 18652
rect 29972 18640 29978 18692
rect 30006 18640 30012 18692
rect 30064 18680 30070 18692
rect 30101 18683 30159 18689
rect 30101 18680 30113 18683
rect 30064 18652 30113 18680
rect 30064 18640 30070 18652
rect 30101 18649 30113 18652
rect 30147 18680 30159 18683
rect 30852 18680 30880 18711
rect 32306 18708 32312 18720
rect 32364 18708 32370 18760
rect 32490 18757 32496 18760
rect 32484 18748 32496 18757
rect 32451 18720 32496 18748
rect 32484 18711 32496 18720
rect 32490 18708 32496 18711
rect 32548 18708 32554 18760
rect 38930 18748 38936 18760
rect 38891 18720 38936 18748
rect 38930 18708 38936 18720
rect 38988 18708 38994 18760
rect 39022 18708 39028 18760
rect 39080 18748 39086 18760
rect 39080 18720 39125 18748
rect 39080 18708 39086 18720
rect 39574 18708 39580 18760
rect 39632 18748 39638 18760
rect 40221 18751 40279 18757
rect 40221 18748 40233 18751
rect 39632 18720 40233 18748
rect 39632 18708 39638 18720
rect 40221 18717 40233 18720
rect 40267 18717 40279 18751
rect 40221 18711 40279 18717
rect 42058 18680 42064 18692
rect 30147 18652 30880 18680
rect 42019 18652 42064 18680
rect 30147 18649 30159 18652
rect 30101 18643 30159 18649
rect 42058 18640 42064 18652
rect 42116 18640 42122 18692
rect 14921 18615 14979 18621
rect 14921 18581 14933 18615
rect 14967 18612 14979 18615
rect 15930 18612 15936 18624
rect 14967 18584 15936 18612
rect 14967 18581 14979 18584
rect 14921 18575 14979 18581
rect 15930 18572 15936 18584
rect 15988 18572 15994 18624
rect 19705 18615 19763 18621
rect 19705 18581 19717 18615
rect 19751 18612 19763 18615
rect 19978 18612 19984 18624
rect 19751 18584 19984 18612
rect 19751 18581 19763 18584
rect 19705 18575 19763 18581
rect 19978 18572 19984 18584
rect 20036 18572 20042 18624
rect 22281 18615 22339 18621
rect 22281 18581 22293 18615
rect 22327 18612 22339 18615
rect 24486 18612 24492 18624
rect 22327 18584 24492 18612
rect 22327 18581 22339 18584
rect 22281 18575 22339 18581
rect 24486 18572 24492 18584
rect 24544 18572 24550 18624
rect 28997 18615 29055 18621
rect 28997 18581 29009 18615
rect 29043 18612 29055 18615
rect 29086 18612 29092 18624
rect 29043 18584 29092 18612
rect 29043 18581 29055 18584
rect 28997 18575 29055 18581
rect 29086 18572 29092 18584
rect 29144 18572 29150 18624
rect 29549 18615 29607 18621
rect 29549 18581 29561 18615
rect 29595 18612 29607 18615
rect 29638 18612 29644 18624
rect 29595 18584 29644 18612
rect 29595 18581 29607 18584
rect 29549 18575 29607 18581
rect 29638 18572 29644 18584
rect 29696 18572 29702 18624
rect 30742 18612 30748 18624
rect 30703 18584 30748 18612
rect 30742 18572 30748 18584
rect 30800 18572 30806 18624
rect 39209 18615 39267 18621
rect 39209 18581 39221 18615
rect 39255 18612 39267 18615
rect 39390 18612 39396 18624
rect 39255 18584 39396 18612
rect 39255 18581 39267 18584
rect 39209 18575 39267 18581
rect 39390 18572 39396 18584
rect 39448 18572 39454 18624
rect 1104 18522 42872 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 42872 18522
rect 1104 18448 42872 18470
rect 16206 18368 16212 18420
rect 16264 18408 16270 18420
rect 22278 18408 22284 18420
rect 16264 18380 17724 18408
rect 22239 18380 22284 18408
rect 16264 18368 16270 18380
rect 12894 18340 12900 18352
rect 11532 18312 12900 18340
rect 11532 18216 11560 18312
rect 12894 18300 12900 18312
rect 12952 18300 12958 18352
rect 16117 18343 16175 18349
rect 16117 18309 16129 18343
rect 16163 18340 16175 18343
rect 17589 18343 17647 18349
rect 17589 18340 17601 18343
rect 16163 18312 17601 18340
rect 16163 18309 16175 18312
rect 16117 18303 16175 18309
rect 17589 18309 17601 18312
rect 17635 18309 17647 18343
rect 17589 18303 17647 18309
rect 11784 18275 11842 18281
rect 11784 18241 11796 18275
rect 11830 18272 11842 18275
rect 13722 18272 13728 18284
rect 11830 18244 13728 18272
rect 11830 18241 11842 18244
rect 11784 18235 11842 18241
rect 13722 18232 13728 18244
rect 13780 18232 13786 18284
rect 15197 18275 15255 18281
rect 15197 18272 15209 18275
rect 14476 18244 15209 18272
rect 11514 18204 11520 18216
rect 11475 18176 11520 18204
rect 11514 18164 11520 18176
rect 11572 18164 11578 18216
rect 14476 18213 14504 18244
rect 15197 18241 15209 18244
rect 15243 18241 15255 18275
rect 15838 18272 15844 18284
rect 15802 18244 15844 18272
rect 15197 18235 15255 18241
rect 15838 18232 15844 18244
rect 15896 18232 15902 18284
rect 15930 18232 15936 18284
rect 15988 18272 15994 18284
rect 15988 18244 16033 18272
rect 15988 18232 15994 18244
rect 16574 18232 16580 18284
rect 16632 18272 16638 18284
rect 16669 18275 16727 18281
rect 16669 18272 16681 18275
rect 16632 18244 16681 18272
rect 16632 18232 16638 18244
rect 16669 18241 16681 18244
rect 16715 18241 16727 18275
rect 16669 18235 16727 18241
rect 16853 18275 16911 18281
rect 16853 18241 16865 18275
rect 16899 18241 16911 18275
rect 16853 18235 16911 18241
rect 14461 18207 14519 18213
rect 14461 18173 14473 18207
rect 14507 18173 14519 18207
rect 14918 18204 14924 18216
rect 14879 18176 14924 18204
rect 14461 18167 14519 18173
rect 12897 18139 12955 18145
rect 12897 18105 12909 18139
rect 12943 18136 12955 18139
rect 14476 18136 14504 18167
rect 14918 18164 14924 18176
rect 14976 18164 14982 18216
rect 15010 18164 15016 18216
rect 15068 18204 15074 18216
rect 16868 18204 16896 18235
rect 16942 18232 16948 18284
rect 17000 18272 17006 18284
rect 17696 18281 17724 18380
rect 22278 18368 22284 18380
rect 22336 18368 22342 18420
rect 28629 18411 28687 18417
rect 28629 18377 28641 18411
rect 28675 18408 28687 18411
rect 28718 18408 28724 18420
rect 28675 18380 28724 18408
rect 28675 18377 28687 18380
rect 28629 18371 28687 18377
rect 28718 18368 28724 18380
rect 28776 18368 28782 18420
rect 30006 18408 30012 18420
rect 28966 18380 30012 18408
rect 28966 18340 28994 18380
rect 28736 18312 28994 18340
rect 17497 18275 17555 18281
rect 17497 18272 17509 18275
rect 17000 18244 17509 18272
rect 17000 18232 17006 18244
rect 17497 18241 17509 18244
rect 17543 18241 17555 18275
rect 17497 18235 17555 18241
rect 17681 18275 17739 18281
rect 17681 18241 17693 18275
rect 17727 18272 17739 18275
rect 18046 18272 18052 18284
rect 17727 18244 18052 18272
rect 17727 18241 17739 18244
rect 17681 18235 17739 18241
rect 18046 18232 18052 18244
rect 18104 18232 18110 18284
rect 18601 18275 18659 18281
rect 18601 18241 18613 18275
rect 18647 18272 18659 18275
rect 18690 18272 18696 18284
rect 18647 18244 18696 18272
rect 18647 18241 18659 18244
rect 18601 18235 18659 18241
rect 18616 18204 18644 18235
rect 18690 18232 18696 18244
rect 18748 18232 18754 18284
rect 18874 18272 18880 18284
rect 18835 18244 18880 18272
rect 18874 18232 18880 18244
rect 18932 18232 18938 18284
rect 19978 18272 19984 18284
rect 19939 18244 19984 18272
rect 19978 18232 19984 18244
rect 20036 18232 20042 18284
rect 28626 18232 28632 18284
rect 28684 18272 28690 18284
rect 28736 18281 28764 18312
rect 29086 18300 29092 18352
rect 29144 18340 29150 18352
rect 29454 18349 29460 18352
rect 29144 18312 29224 18340
rect 29144 18300 29150 18312
rect 29196 18281 29224 18312
rect 29449 18303 29460 18349
rect 29512 18340 29518 18352
rect 29512 18312 29549 18340
rect 29454 18300 29460 18303
rect 29512 18300 29518 18312
rect 29625 18281 29653 18380
rect 30006 18368 30012 18380
rect 30064 18368 30070 18420
rect 38930 18408 38936 18420
rect 38891 18380 38936 18408
rect 38930 18368 38936 18380
rect 38988 18368 38994 18420
rect 39574 18408 39580 18420
rect 39535 18380 39580 18408
rect 39574 18368 39580 18380
rect 39632 18368 39638 18420
rect 30098 18300 30104 18352
rect 30156 18340 30162 18352
rect 32217 18343 32275 18349
rect 32217 18340 32229 18343
rect 30156 18312 32229 18340
rect 30156 18300 30162 18312
rect 32217 18309 32229 18312
rect 32263 18309 32275 18343
rect 32217 18303 32275 18309
rect 32306 18300 32312 18352
rect 32364 18340 32370 18352
rect 32401 18343 32459 18349
rect 32401 18340 32413 18343
rect 32364 18312 32413 18340
rect 32364 18300 32370 18312
rect 32401 18309 32413 18312
rect 32447 18340 32459 18343
rect 37820 18343 37878 18349
rect 32447 18312 36400 18340
rect 32447 18309 32459 18312
rect 32401 18303 32459 18309
rect 28721 18275 28779 18281
rect 28721 18272 28733 18275
rect 28684 18244 28733 18272
rect 28684 18232 28690 18244
rect 28721 18241 28733 18244
rect 28767 18241 28779 18275
rect 28721 18235 28779 18241
rect 29181 18275 29239 18281
rect 29181 18241 29193 18275
rect 29227 18241 29239 18275
rect 29181 18235 29239 18241
rect 29365 18275 29423 18281
rect 29365 18241 29377 18275
rect 29411 18272 29423 18275
rect 29595 18275 29653 18281
rect 29411 18244 29500 18272
rect 29411 18241 29423 18244
rect 29365 18235 29423 18241
rect 15068 18176 18644 18204
rect 15068 18164 15074 18176
rect 21634 18164 21640 18216
rect 21692 18204 21698 18216
rect 21821 18207 21879 18213
rect 21821 18204 21833 18207
rect 21692 18176 21833 18204
rect 21692 18164 21698 18176
rect 21821 18173 21833 18176
rect 21867 18173 21879 18207
rect 29472 18204 29500 18244
rect 29595 18241 29607 18275
rect 29641 18241 29653 18275
rect 30650 18272 30656 18284
rect 30611 18244 30656 18272
rect 29595 18235 29653 18241
rect 30650 18232 30656 18244
rect 30708 18272 30714 18284
rect 33428 18281 33456 18312
rect 36372 18284 36400 18312
rect 37820 18309 37832 18343
rect 37866 18340 37878 18343
rect 38010 18340 38016 18352
rect 37866 18312 38016 18340
rect 37866 18309 37878 18312
rect 37820 18303 37878 18309
rect 38010 18300 38016 18312
rect 38068 18300 38074 18352
rect 33413 18275 33471 18281
rect 30708 18244 31754 18272
rect 30708 18232 30714 18244
rect 30561 18207 30619 18213
rect 30561 18204 30573 18207
rect 29472 18176 30573 18204
rect 21821 18167 21879 18173
rect 30561 18173 30573 18176
rect 30607 18204 30619 18207
rect 30742 18204 30748 18216
rect 30607 18176 30748 18204
rect 30607 18173 30619 18176
rect 30561 18167 30619 18173
rect 30742 18164 30748 18176
rect 30800 18164 30806 18216
rect 31726 18204 31754 18244
rect 33413 18241 33425 18275
rect 33459 18241 33471 18275
rect 33669 18275 33727 18281
rect 33669 18272 33681 18275
rect 33413 18235 33471 18241
rect 33520 18244 33681 18272
rect 33520 18204 33548 18244
rect 33669 18241 33681 18244
rect 33715 18241 33727 18275
rect 33669 18235 33727 18241
rect 36354 18232 36360 18284
rect 36412 18272 36418 18284
rect 37550 18272 37556 18284
rect 36412 18244 37556 18272
rect 36412 18232 36418 18244
rect 37550 18232 37556 18244
rect 37608 18232 37614 18284
rect 39390 18272 39396 18284
rect 39351 18244 39396 18272
rect 39390 18232 39396 18244
rect 39448 18232 39454 18284
rect 41322 18204 41328 18216
rect 31726 18176 33548 18204
rect 41283 18176 41328 18204
rect 41322 18164 41328 18176
rect 41380 18164 41386 18216
rect 41690 18204 41696 18216
rect 41651 18176 41696 18204
rect 41690 18164 41696 18176
rect 41748 18164 41754 18216
rect 41874 18204 41880 18216
rect 41835 18176 41880 18204
rect 41874 18164 41880 18176
rect 41932 18164 41938 18216
rect 12943 18108 14504 18136
rect 14936 18136 14964 18164
rect 15194 18136 15200 18148
rect 14936 18108 15200 18136
rect 12943 18105 12955 18108
rect 12897 18099 12955 18105
rect 15194 18096 15200 18108
rect 15252 18096 15258 18148
rect 15654 18096 15660 18148
rect 15712 18136 15718 18148
rect 16117 18139 16175 18145
rect 16117 18136 16129 18139
rect 15712 18108 16129 18136
rect 15712 18096 15718 18108
rect 16117 18105 16129 18108
rect 16163 18105 16175 18139
rect 16117 18099 16175 18105
rect 20070 18096 20076 18148
rect 20128 18136 20134 18148
rect 22189 18139 22247 18145
rect 22189 18136 22201 18139
rect 20128 18108 22201 18136
rect 20128 18096 20134 18108
rect 22189 18105 22201 18108
rect 22235 18136 22247 18139
rect 32122 18136 32128 18148
rect 22235 18108 32128 18136
rect 22235 18105 22247 18108
rect 22189 18099 22247 18105
rect 32122 18096 32128 18108
rect 32180 18096 32186 18148
rect 13538 18028 13544 18080
rect 13596 18068 13602 18080
rect 14231 18071 14289 18077
rect 14231 18068 14243 18071
rect 13596 18040 14243 18068
rect 13596 18028 13602 18040
rect 14231 18037 14243 18040
rect 14277 18068 14289 18071
rect 14734 18068 14740 18080
rect 14277 18040 14740 18068
rect 14277 18037 14289 18040
rect 14231 18031 14289 18037
rect 14734 18028 14740 18040
rect 14792 18028 14798 18080
rect 15102 18028 15108 18080
rect 15160 18068 15166 18080
rect 15381 18071 15439 18077
rect 15381 18068 15393 18071
rect 15160 18040 15393 18068
rect 15160 18028 15166 18040
rect 15381 18037 15393 18040
rect 15427 18037 15439 18071
rect 15381 18031 15439 18037
rect 16482 18028 16488 18080
rect 16540 18068 16546 18080
rect 17037 18071 17095 18077
rect 17037 18068 17049 18071
rect 16540 18040 17049 18068
rect 16540 18028 16546 18040
rect 17037 18037 17049 18040
rect 17083 18037 17095 18071
rect 20162 18068 20168 18080
rect 20123 18040 20168 18068
rect 17037 18031 17095 18037
rect 20162 18028 20168 18040
rect 20220 18028 20226 18080
rect 29730 18068 29736 18080
rect 29691 18040 29736 18068
rect 29730 18028 29736 18040
rect 29788 18028 29794 18080
rect 31018 18068 31024 18080
rect 30979 18040 31024 18068
rect 31018 18028 31024 18040
rect 31076 18028 31082 18080
rect 34790 18068 34796 18080
rect 34751 18040 34796 18068
rect 34790 18028 34796 18040
rect 34848 18028 34854 18080
rect 1104 17978 42872 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 42872 17978
rect 1104 17904 42872 17926
rect 13722 17824 13728 17876
rect 13780 17864 13786 17876
rect 14093 17867 14151 17873
rect 14093 17864 14105 17867
rect 13780 17836 14105 17864
rect 13780 17824 13786 17836
rect 14093 17833 14105 17836
rect 14139 17833 14151 17867
rect 14093 17827 14151 17833
rect 14458 17824 14464 17876
rect 14516 17864 14522 17876
rect 14516 17836 14780 17864
rect 14516 17824 14522 17836
rect 13541 17799 13599 17805
rect 13541 17765 13553 17799
rect 13587 17796 13599 17799
rect 14366 17796 14372 17808
rect 13587 17768 14372 17796
rect 13587 17765 13599 17768
rect 13541 17759 13599 17765
rect 14366 17756 14372 17768
rect 14424 17756 14430 17808
rect 14752 17796 14780 17836
rect 14918 17824 14924 17876
rect 14976 17864 14982 17876
rect 15197 17867 15255 17873
rect 15197 17864 15209 17867
rect 14976 17836 15209 17864
rect 14976 17824 14982 17836
rect 15197 17833 15209 17836
rect 15243 17833 15255 17867
rect 15197 17827 15255 17833
rect 15378 17824 15384 17876
rect 15436 17864 15442 17876
rect 15436 17836 15976 17864
rect 15436 17824 15442 17836
rect 15948 17808 15976 17836
rect 16114 17824 16120 17876
rect 16172 17864 16178 17876
rect 16669 17867 16727 17873
rect 16669 17864 16681 17867
rect 16172 17836 16681 17864
rect 16172 17824 16178 17836
rect 16669 17833 16681 17836
rect 16715 17833 16727 17867
rect 16669 17827 16727 17833
rect 16853 17867 16911 17873
rect 16853 17833 16865 17867
rect 16899 17864 16911 17867
rect 17586 17864 17592 17876
rect 16899 17836 17592 17864
rect 16899 17833 16911 17836
rect 16853 17827 16911 17833
rect 17586 17824 17592 17836
rect 17644 17824 17650 17876
rect 26234 17824 26240 17876
rect 26292 17864 26298 17876
rect 30006 17864 30012 17876
rect 26292 17836 30012 17864
rect 26292 17824 26298 17836
rect 30006 17824 30012 17836
rect 30064 17824 30070 17876
rect 40034 17824 40040 17876
rect 40092 17864 40098 17876
rect 40681 17867 40739 17873
rect 40681 17864 40693 17867
rect 40092 17836 40693 17864
rect 40092 17824 40098 17836
rect 40681 17833 40693 17836
rect 40727 17833 40739 17867
rect 40681 17827 40739 17833
rect 41417 17867 41475 17873
rect 41417 17833 41429 17867
rect 41463 17864 41475 17867
rect 41690 17864 41696 17876
rect 41463 17836 41696 17864
rect 41463 17833 41475 17836
rect 41417 17827 41475 17833
rect 41690 17824 41696 17836
rect 41748 17824 41754 17876
rect 41874 17824 41880 17876
rect 41932 17864 41938 17876
rect 41969 17867 42027 17873
rect 41969 17864 41981 17867
rect 41932 17836 41981 17864
rect 41932 17824 41938 17836
rect 41969 17833 41981 17836
rect 42015 17833 42027 17867
rect 41969 17827 42027 17833
rect 14752 17768 15792 17796
rect 14642 17728 14648 17740
rect 14384 17700 14648 17728
rect 1946 17620 1952 17672
rect 2004 17660 2010 17672
rect 2041 17663 2099 17669
rect 2041 17660 2053 17663
rect 2004 17632 2053 17660
rect 2004 17620 2010 17632
rect 2041 17629 2053 17632
rect 2087 17629 2099 17663
rect 2041 17623 2099 17629
rect 2961 17663 3019 17669
rect 2961 17629 2973 17663
rect 3007 17660 3019 17663
rect 11057 17663 11115 17669
rect 11057 17660 11069 17663
rect 3007 17632 11069 17660
rect 3007 17629 3019 17632
rect 2961 17623 3019 17629
rect 11057 17629 11069 17632
rect 11103 17660 11115 17663
rect 11146 17660 11152 17672
rect 11103 17632 11152 17660
rect 11103 17629 11115 17632
rect 11057 17623 11115 17629
rect 11146 17620 11152 17632
rect 11204 17620 11210 17672
rect 11238 17620 11244 17672
rect 11296 17660 11302 17672
rect 11517 17663 11575 17669
rect 11517 17660 11529 17663
rect 11296 17632 11529 17660
rect 11296 17620 11302 17632
rect 11517 17629 11529 17632
rect 11563 17629 11575 17663
rect 13262 17660 13268 17672
rect 13223 17632 13268 17660
rect 11517 17623 11575 17629
rect 13262 17620 13268 17632
rect 13320 17620 13326 17672
rect 14090 17620 14096 17672
rect 14148 17660 14154 17672
rect 14384 17669 14412 17700
rect 14642 17688 14648 17700
rect 14700 17688 14706 17740
rect 15764 17728 15792 17768
rect 15930 17756 15936 17808
rect 15988 17796 15994 17808
rect 19337 17799 19395 17805
rect 19337 17796 19349 17799
rect 15988 17768 19349 17796
rect 15988 17756 15994 17768
rect 19337 17765 19349 17768
rect 19383 17765 19395 17799
rect 19337 17759 19395 17765
rect 29454 17756 29460 17808
rect 29512 17796 29518 17808
rect 30745 17799 30803 17805
rect 30745 17796 30757 17799
rect 29512 17768 30757 17796
rect 29512 17756 29518 17768
rect 30745 17765 30757 17768
rect 30791 17765 30803 17799
rect 30745 17759 30803 17765
rect 17954 17728 17960 17740
rect 15764 17700 16804 17728
rect 14277 17663 14335 17669
rect 14277 17660 14289 17663
rect 14148 17632 14289 17660
rect 14148 17620 14154 17632
rect 14277 17629 14289 17632
rect 14323 17629 14335 17663
rect 14277 17623 14335 17629
rect 14369 17663 14427 17669
rect 14369 17629 14381 17663
rect 14415 17629 14427 17663
rect 14734 17660 14740 17672
rect 14695 17632 14740 17660
rect 14369 17623 14427 17629
rect 14734 17620 14740 17632
rect 14792 17620 14798 17672
rect 15335 17629 15393 17635
rect 15335 17604 15347 17629
rect 13538 17592 13544 17604
rect 13499 17564 13544 17592
rect 13538 17552 13544 17564
rect 13596 17552 13602 17604
rect 13722 17552 13728 17604
rect 13780 17592 13786 17604
rect 14458 17592 14464 17604
rect 13780 17564 14464 17592
rect 13780 17552 13786 17564
rect 14458 17552 14464 17564
rect 14516 17552 14522 17604
rect 14550 17552 14556 17604
rect 14608 17601 14614 17604
rect 14608 17595 14637 17601
rect 14625 17561 14637 17595
rect 14608 17555 14637 17561
rect 14608 17552 14614 17555
rect 15286 17552 15292 17604
rect 15344 17595 15347 17604
rect 15381 17626 15393 17629
rect 15381 17595 15408 17626
rect 15580 17601 15700 17626
rect 15344 17564 15408 17595
rect 15565 17598 15700 17601
rect 15565 17595 15623 17598
rect 15344 17552 15350 17564
rect 15565 17561 15577 17595
rect 15611 17561 15623 17595
rect 15672 17592 15700 17598
rect 15746 17592 15752 17604
rect 15672 17564 15752 17592
rect 15565 17555 15623 17561
rect 15746 17552 15752 17564
rect 15804 17552 15810 17604
rect 16482 17592 16488 17604
rect 16443 17564 16488 17592
rect 16482 17552 16488 17564
rect 16540 17552 16546 17604
rect 16666 17552 16672 17604
rect 16724 17601 16730 17604
rect 16724 17595 16743 17601
rect 16731 17561 16743 17595
rect 16776 17592 16804 17700
rect 17788 17700 17960 17728
rect 17788 17669 17816 17700
rect 17954 17688 17960 17700
rect 18012 17688 18018 17740
rect 18966 17728 18972 17740
rect 18064 17700 18972 17728
rect 17773 17663 17831 17669
rect 17773 17629 17785 17663
rect 17819 17629 17831 17663
rect 17773 17623 17831 17629
rect 17862 17620 17868 17672
rect 17920 17660 17926 17672
rect 18064 17669 18092 17700
rect 18966 17688 18972 17700
rect 19024 17728 19030 17740
rect 19245 17731 19303 17737
rect 19245 17728 19257 17731
rect 19024 17700 19257 17728
rect 19024 17688 19030 17700
rect 19245 17697 19257 17700
rect 19291 17697 19303 17731
rect 19245 17691 19303 17697
rect 28997 17731 29055 17737
rect 28997 17697 29009 17731
rect 29043 17728 29055 17731
rect 29362 17728 29368 17740
rect 29043 17700 29368 17728
rect 29043 17697 29055 17700
rect 28997 17691 29055 17697
rect 29362 17688 29368 17700
rect 29420 17728 29426 17740
rect 31297 17731 31355 17737
rect 31297 17728 31309 17731
rect 29420 17700 31309 17728
rect 29420 17688 29426 17700
rect 31297 17697 31309 17700
rect 31343 17697 31355 17731
rect 36354 17728 36360 17740
rect 36315 17700 36360 17728
rect 31297 17691 31355 17697
rect 36354 17688 36360 17700
rect 36412 17688 36418 17740
rect 39022 17728 39028 17740
rect 38488 17700 39028 17728
rect 38488 17672 38516 17700
rect 39022 17688 39028 17700
rect 39080 17688 39086 17740
rect 18049 17663 18107 17669
rect 17920 17632 17965 17660
rect 17920 17620 17926 17632
rect 18049 17629 18061 17663
rect 18095 17629 18107 17663
rect 18049 17623 18107 17629
rect 18141 17663 18199 17669
rect 18141 17629 18153 17663
rect 18187 17660 18199 17663
rect 18322 17660 18328 17672
rect 18187 17632 18328 17660
rect 18187 17629 18199 17632
rect 18141 17623 18199 17629
rect 18322 17620 18328 17632
rect 18380 17620 18386 17672
rect 19521 17663 19579 17669
rect 19521 17629 19533 17663
rect 19567 17660 19579 17663
rect 20070 17660 20076 17672
rect 19567 17632 20076 17660
rect 19567 17629 19579 17632
rect 19521 17623 19579 17629
rect 20070 17620 20076 17632
rect 20128 17620 20134 17672
rect 20257 17663 20315 17669
rect 20257 17629 20269 17663
rect 20303 17660 20315 17663
rect 20898 17660 20904 17672
rect 20303 17632 20904 17660
rect 20303 17629 20315 17632
rect 20257 17623 20315 17629
rect 20898 17620 20904 17632
rect 20956 17660 20962 17672
rect 22465 17663 22523 17669
rect 22465 17660 22477 17663
rect 20956 17632 22477 17660
rect 20956 17620 20962 17632
rect 22465 17629 22477 17632
rect 22511 17629 22523 17663
rect 22465 17623 22523 17629
rect 27157 17663 27215 17669
rect 27157 17629 27169 17663
rect 27203 17660 27215 17663
rect 27798 17660 27804 17672
rect 27203 17632 27804 17660
rect 27203 17629 27215 17632
rect 27157 17623 27215 17629
rect 27798 17620 27804 17632
rect 27856 17620 27862 17672
rect 28718 17620 28724 17672
rect 28776 17669 28782 17672
rect 28776 17660 28788 17669
rect 28776 17632 28821 17660
rect 28776 17623 28788 17632
rect 28776 17620 28782 17623
rect 29914 17620 29920 17672
rect 29972 17660 29978 17672
rect 30653 17663 30711 17669
rect 30653 17660 30665 17663
rect 29972 17632 30665 17660
rect 29972 17620 29978 17632
rect 30653 17629 30665 17632
rect 30699 17629 30711 17663
rect 30653 17623 30711 17629
rect 31018 17620 31024 17672
rect 31076 17660 31082 17672
rect 31553 17663 31611 17669
rect 31553 17660 31565 17663
rect 31076 17632 31565 17660
rect 31076 17620 31082 17632
rect 31553 17629 31565 17632
rect 31599 17629 31611 17663
rect 34790 17660 34796 17672
rect 34751 17632 34796 17660
rect 31553 17623 31611 17629
rect 34790 17620 34796 17632
rect 34848 17620 34854 17672
rect 34974 17660 34980 17672
rect 34935 17632 34980 17660
rect 34974 17620 34980 17632
rect 35032 17620 35038 17672
rect 36630 17669 36636 17672
rect 36624 17660 36636 17669
rect 36591 17632 36636 17660
rect 36624 17623 36636 17632
rect 36630 17620 36636 17623
rect 36688 17620 36694 17672
rect 38470 17660 38476 17672
rect 38431 17632 38476 17660
rect 38470 17620 38476 17632
rect 38528 17620 38534 17672
rect 38746 17660 38752 17672
rect 38707 17632 38752 17660
rect 38746 17620 38752 17632
rect 38804 17620 38810 17672
rect 39758 17620 39764 17672
rect 39816 17660 39822 17672
rect 41138 17660 41144 17672
rect 39816 17632 41144 17660
rect 39816 17620 39822 17632
rect 41138 17620 41144 17632
rect 41196 17660 41202 17672
rect 41325 17663 41383 17669
rect 41325 17660 41337 17663
rect 41196 17632 41337 17660
rect 41196 17620 41202 17632
rect 41325 17629 41337 17632
rect 41371 17629 41383 17663
rect 41325 17623 41383 17629
rect 19978 17592 19984 17604
rect 16776 17564 19984 17592
rect 16724 17555 16743 17561
rect 16724 17552 16730 17555
rect 19978 17552 19984 17564
rect 20036 17552 20042 17604
rect 20162 17552 20168 17604
rect 20220 17592 20226 17604
rect 20502 17595 20560 17601
rect 20502 17592 20514 17595
rect 20220 17564 20514 17592
rect 20220 17552 20226 17564
rect 20502 17561 20514 17564
rect 20548 17561 20560 17595
rect 22710 17595 22768 17601
rect 22710 17592 22722 17595
rect 20502 17555 20560 17561
rect 20916 17564 22722 17592
rect 2130 17484 2136 17536
rect 2188 17524 2194 17536
rect 2869 17527 2927 17533
rect 2869 17524 2881 17527
rect 2188 17496 2881 17524
rect 2188 17484 2194 17496
rect 2869 17493 2881 17496
rect 2915 17493 2927 17527
rect 2869 17487 2927 17493
rect 13357 17527 13415 17533
rect 13357 17493 13369 17527
rect 13403 17524 13415 17527
rect 15378 17524 15384 17536
rect 13403 17496 15384 17524
rect 13403 17493 13415 17496
rect 13357 17487 13415 17493
rect 15378 17484 15384 17496
rect 15436 17484 15442 17536
rect 17126 17484 17132 17536
rect 17184 17524 17190 17536
rect 17589 17527 17647 17533
rect 17589 17524 17601 17527
rect 17184 17496 17601 17524
rect 17184 17484 17190 17496
rect 17589 17493 17601 17496
rect 17635 17493 17647 17527
rect 17589 17487 17647 17493
rect 19705 17527 19763 17533
rect 19705 17493 19717 17527
rect 19751 17524 19763 17527
rect 20916 17524 20944 17564
rect 22710 17561 22722 17564
rect 22756 17561 22768 17595
rect 22710 17555 22768 17561
rect 26878 17552 26884 17604
rect 26936 17601 26942 17604
rect 26936 17592 26948 17601
rect 30006 17592 30012 17604
rect 26936 17564 26981 17592
rect 27540 17564 28764 17592
rect 29967 17564 30012 17592
rect 26936 17555 26948 17564
rect 26936 17552 26942 17555
rect 19751 17496 20944 17524
rect 21637 17527 21695 17533
rect 19751 17493 19763 17496
rect 19705 17487 19763 17493
rect 21637 17493 21649 17527
rect 21683 17524 21695 17527
rect 23658 17524 23664 17536
rect 21683 17496 23664 17524
rect 21683 17493 21695 17496
rect 21637 17487 21695 17493
rect 23658 17484 23664 17496
rect 23716 17484 23722 17536
rect 23842 17524 23848 17536
rect 23803 17496 23848 17524
rect 23842 17484 23848 17496
rect 23900 17484 23906 17536
rect 25777 17527 25835 17533
rect 25777 17493 25789 17527
rect 25823 17524 25835 17527
rect 27540 17524 27568 17564
rect 25823 17496 27568 17524
rect 27617 17527 27675 17533
rect 25823 17493 25835 17496
rect 25777 17487 25835 17493
rect 27617 17493 27629 17527
rect 27663 17524 27675 17527
rect 28626 17524 28632 17536
rect 27663 17496 28632 17524
rect 27663 17493 27675 17496
rect 27617 17487 27675 17493
rect 28626 17484 28632 17496
rect 28684 17484 28690 17536
rect 28736 17524 28764 17564
rect 30006 17552 30012 17564
rect 30064 17552 30070 17604
rect 28994 17524 29000 17536
rect 28736 17496 29000 17524
rect 28994 17484 29000 17496
rect 29052 17484 29058 17536
rect 30098 17524 30104 17536
rect 30059 17496 30104 17524
rect 30098 17484 30104 17496
rect 30156 17484 30162 17536
rect 32582 17484 32588 17536
rect 32640 17524 32646 17536
rect 32677 17527 32735 17533
rect 32677 17524 32689 17527
rect 32640 17496 32689 17524
rect 32640 17484 32646 17496
rect 32677 17493 32689 17496
rect 32723 17493 32735 17527
rect 32677 17487 32735 17493
rect 34790 17484 34796 17536
rect 34848 17524 34854 17536
rect 34885 17527 34943 17533
rect 34885 17524 34897 17527
rect 34848 17496 34897 17524
rect 34848 17484 34854 17496
rect 34885 17493 34897 17496
rect 34931 17493 34943 17527
rect 34885 17487 34943 17493
rect 37737 17527 37795 17533
rect 37737 17493 37749 17527
rect 37783 17524 37795 17527
rect 37918 17524 37924 17536
rect 37783 17496 37924 17524
rect 37783 17493 37795 17496
rect 37737 17487 37795 17493
rect 37918 17484 37924 17496
rect 37976 17484 37982 17536
rect 1104 17434 42872 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 42872 17434
rect 1104 17360 42872 17382
rect 13354 17280 13360 17332
rect 13412 17320 13418 17332
rect 13412 17292 14044 17320
rect 13412 17280 13418 17292
rect 2130 17252 2136 17264
rect 2091 17224 2136 17252
rect 2130 17212 2136 17224
rect 2188 17212 2194 17264
rect 13722 17252 13728 17264
rect 13683 17224 13728 17252
rect 13722 17212 13728 17224
rect 13780 17212 13786 17264
rect 14016 17252 14044 17292
rect 14090 17280 14096 17332
rect 14148 17320 14154 17332
rect 14553 17323 14611 17329
rect 14553 17320 14565 17323
rect 14148 17292 14565 17320
rect 14148 17280 14154 17292
rect 14553 17289 14565 17292
rect 14599 17289 14611 17323
rect 17954 17320 17960 17332
rect 14553 17283 14611 17289
rect 14660 17292 17960 17320
rect 14660 17252 14688 17292
rect 17954 17280 17960 17292
rect 18012 17280 18018 17332
rect 18966 17320 18972 17332
rect 18927 17292 18972 17320
rect 18966 17280 18972 17292
rect 19024 17280 19030 17332
rect 39758 17320 39764 17332
rect 22066 17292 39764 17320
rect 15194 17252 15200 17264
rect 14016 17224 14688 17252
rect 15155 17224 15200 17252
rect 1946 17184 1952 17196
rect 1907 17156 1952 17184
rect 1946 17144 1952 17156
rect 2004 17144 2010 17196
rect 11514 17184 11520 17196
rect 11475 17156 11520 17184
rect 11514 17144 11520 17156
rect 11572 17144 11578 17196
rect 11784 17187 11842 17193
rect 11784 17153 11796 17187
rect 11830 17184 11842 17187
rect 13357 17187 13415 17193
rect 13357 17184 13369 17187
rect 11830 17156 13369 17184
rect 11830 17153 11842 17156
rect 11784 17147 11842 17153
rect 13357 17153 13369 17156
rect 13403 17153 13415 17187
rect 13357 17147 13415 17153
rect 13446 17144 13452 17196
rect 13504 17184 13510 17196
rect 13541 17187 13599 17193
rect 13541 17184 13553 17187
rect 13504 17156 13553 17184
rect 13504 17144 13510 17156
rect 13541 17153 13553 17156
rect 13587 17153 13599 17187
rect 13541 17147 13599 17153
rect 13630 17144 13636 17196
rect 13688 17184 13694 17196
rect 14016 17193 14044 17224
rect 15194 17212 15200 17224
rect 15252 17212 15258 17264
rect 17862 17212 17868 17264
rect 17920 17252 17926 17264
rect 22066 17252 22094 17292
rect 39758 17280 39764 17292
rect 39816 17280 39822 17332
rect 17920 17224 19012 17252
rect 17920 17212 17926 17224
rect 13843 17187 13901 17193
rect 13688 17156 13733 17184
rect 13688 17144 13694 17156
rect 13843 17153 13855 17187
rect 13889 17153 13901 17187
rect 13843 17147 13901 17153
rect 14001 17187 14059 17193
rect 14001 17153 14013 17187
rect 14047 17153 14059 17187
rect 14001 17147 14059 17153
rect 2774 17116 2780 17128
rect 2735 17088 2780 17116
rect 2774 17076 2780 17088
rect 2832 17076 2838 17128
rect 13858 17116 13886 17147
rect 14366 17144 14372 17196
rect 14424 17184 14430 17196
rect 14461 17187 14519 17193
rect 14461 17184 14473 17187
rect 14424 17156 14473 17184
rect 14424 17144 14430 17156
rect 14461 17153 14473 17156
rect 14507 17153 14519 17187
rect 14461 17147 14519 17153
rect 14645 17187 14703 17193
rect 14645 17153 14657 17187
rect 14691 17184 14703 17187
rect 14918 17184 14924 17196
rect 14691 17156 14924 17184
rect 14691 17153 14703 17156
rect 14645 17147 14703 17153
rect 13858 17088 13952 17116
rect 12897 16983 12955 16989
rect 12897 16949 12909 16983
rect 12943 16980 12955 16983
rect 13814 16980 13820 16992
rect 12943 16952 13820 16980
rect 12943 16949 12955 16952
rect 12897 16943 12955 16949
rect 13814 16940 13820 16952
rect 13872 16940 13878 16992
rect 13924 16980 13952 17088
rect 14274 17076 14280 17128
rect 14332 17116 14338 17128
rect 14660 17116 14688 17147
rect 14918 17144 14924 17156
rect 14976 17144 14982 17196
rect 15470 17184 15476 17196
rect 15431 17156 15476 17184
rect 15470 17144 15476 17156
rect 15528 17144 15534 17196
rect 15746 17184 15752 17196
rect 15580 17156 15752 17184
rect 14332 17088 14688 17116
rect 14332 17076 14338 17088
rect 14734 17076 14740 17128
rect 14792 17116 14798 17128
rect 15381 17119 15439 17125
rect 15381 17116 15393 17119
rect 14792 17088 15393 17116
rect 14792 17076 14798 17088
rect 15381 17085 15393 17088
rect 15427 17116 15439 17119
rect 15580 17116 15608 17156
rect 15746 17144 15752 17156
rect 15804 17184 15810 17196
rect 17218 17184 17224 17196
rect 15804 17156 17080 17184
rect 17179 17156 17224 17184
rect 15804 17144 15810 17156
rect 16942 17116 16948 17128
rect 15427 17088 15608 17116
rect 16903 17088 16948 17116
rect 15427 17085 15439 17088
rect 15381 17079 15439 17085
rect 16942 17076 16948 17088
rect 17000 17076 17006 17128
rect 17052 17116 17080 17156
rect 17218 17144 17224 17156
rect 17276 17144 17282 17196
rect 18064 17193 18092 17224
rect 18984 17196 19012 17224
rect 19168 17224 22094 17252
rect 18049 17187 18107 17193
rect 18049 17153 18061 17187
rect 18095 17153 18107 17187
rect 18049 17147 18107 17153
rect 18230 17144 18236 17196
rect 18288 17184 18294 17196
rect 18877 17187 18935 17193
rect 18877 17184 18889 17187
rect 18288 17156 18889 17184
rect 18288 17144 18294 17156
rect 18877 17153 18889 17156
rect 18923 17153 18935 17187
rect 18877 17147 18935 17153
rect 18966 17144 18972 17196
rect 19024 17184 19030 17196
rect 19061 17187 19119 17193
rect 19061 17184 19073 17187
rect 19024 17156 19073 17184
rect 19024 17144 19030 17156
rect 19061 17153 19073 17156
rect 19107 17153 19119 17187
rect 19061 17147 19119 17153
rect 18141 17119 18199 17125
rect 18141 17116 18153 17119
rect 17052 17088 18153 17116
rect 18141 17085 18153 17088
rect 18187 17085 18199 17119
rect 18141 17079 18199 17085
rect 14366 17008 14372 17060
rect 14424 17048 14430 17060
rect 19168 17048 19196 17224
rect 29454 17212 29460 17264
rect 29512 17252 29518 17264
rect 29632 17255 29690 17261
rect 29632 17252 29644 17255
rect 29512 17224 29644 17252
rect 29512 17212 29518 17224
rect 29632 17221 29644 17224
rect 29678 17221 29690 17255
rect 34974 17252 34980 17264
rect 29632 17215 29690 17221
rect 34808 17224 34980 17252
rect 20070 17144 20076 17196
rect 20128 17184 20134 17196
rect 20349 17187 20407 17193
rect 20349 17184 20361 17187
rect 20128 17156 20361 17184
rect 20128 17144 20134 17156
rect 20349 17153 20361 17156
rect 20395 17153 20407 17187
rect 20349 17147 20407 17153
rect 21358 17144 21364 17196
rect 21416 17184 21422 17196
rect 21821 17187 21879 17193
rect 21821 17184 21833 17187
rect 21416 17156 21833 17184
rect 21416 17144 21422 17156
rect 21821 17153 21833 17156
rect 21867 17153 21879 17187
rect 22721 17187 22779 17193
rect 22721 17184 22733 17187
rect 21821 17147 21879 17153
rect 22020 17156 22733 17184
rect 19978 17076 19984 17128
rect 20036 17116 20042 17128
rect 20622 17116 20628 17128
rect 20036 17088 20628 17116
rect 20036 17076 20042 17088
rect 20622 17076 20628 17088
rect 20680 17076 20686 17128
rect 22020 17057 22048 17156
rect 22721 17153 22733 17156
rect 22767 17153 22779 17187
rect 22721 17147 22779 17153
rect 24762 17144 24768 17196
rect 24820 17184 24826 17196
rect 25409 17187 25467 17193
rect 25409 17184 25421 17187
rect 24820 17156 25421 17184
rect 24820 17144 24826 17156
rect 25409 17153 25421 17156
rect 25455 17153 25467 17187
rect 25590 17184 25596 17196
rect 25551 17156 25596 17184
rect 25409 17147 25467 17153
rect 25590 17144 25596 17156
rect 25648 17144 25654 17196
rect 29362 17184 29368 17196
rect 29323 17156 29368 17184
rect 29362 17144 29368 17156
rect 29420 17144 29426 17196
rect 34808 17193 34836 17224
rect 34974 17212 34980 17224
rect 35032 17212 35038 17264
rect 38746 17252 38752 17264
rect 37844 17224 38752 17252
rect 34793 17187 34851 17193
rect 34793 17184 34805 17187
rect 29472 17156 34805 17184
rect 22094 17076 22100 17128
rect 22152 17116 22158 17128
rect 22465 17119 22523 17125
rect 22465 17116 22477 17119
rect 22152 17088 22477 17116
rect 22152 17076 22158 17088
rect 22465 17085 22477 17088
rect 22511 17085 22523 17119
rect 22465 17079 22523 17085
rect 26421 17119 26479 17125
rect 26421 17085 26433 17119
rect 26467 17116 26479 17119
rect 26878 17116 26884 17128
rect 26467 17088 26884 17116
rect 26467 17085 26479 17088
rect 26421 17079 26479 17085
rect 26878 17076 26884 17088
rect 26936 17116 26942 17128
rect 29472 17116 29500 17156
rect 34793 17153 34805 17156
rect 34839 17153 34851 17187
rect 34793 17147 34851 17153
rect 34882 17144 34888 17196
rect 34940 17184 34946 17196
rect 37844 17193 37872 17224
rect 38746 17212 38752 17224
rect 38804 17212 38810 17264
rect 37829 17187 37887 17193
rect 34940 17156 34985 17184
rect 34940 17144 34946 17156
rect 37829 17153 37841 17187
rect 37875 17153 37887 17187
rect 37829 17147 37887 17153
rect 37918 17144 37924 17196
rect 37976 17184 37982 17196
rect 37976 17156 38021 17184
rect 37976 17144 37982 17156
rect 26936 17088 29500 17116
rect 26936 17076 26942 17088
rect 14424 17020 19196 17048
rect 22005 17051 22063 17057
rect 14424 17008 14430 17020
rect 22005 17017 22017 17051
rect 22051 17017 22063 17051
rect 22005 17011 22063 17017
rect 14550 16980 14556 16992
rect 13924 16952 14556 16980
rect 14550 16940 14556 16952
rect 14608 16940 14614 16992
rect 15102 16940 15108 16992
rect 15160 16980 15166 16992
rect 15197 16983 15255 16989
rect 15197 16980 15209 16983
rect 15160 16952 15209 16980
rect 15160 16940 15166 16952
rect 15197 16949 15209 16952
rect 15243 16949 15255 16983
rect 15197 16943 15255 16949
rect 15657 16983 15715 16989
rect 15657 16949 15669 16983
rect 15703 16980 15715 16983
rect 16574 16980 16580 16992
rect 15703 16952 16580 16980
rect 15703 16949 15715 16952
rect 15657 16943 15715 16949
rect 16574 16940 16580 16952
rect 16632 16940 16638 16992
rect 16666 16940 16672 16992
rect 16724 16980 16730 16992
rect 17126 16980 17132 16992
rect 16724 16952 16769 16980
rect 17087 16952 17132 16980
rect 16724 16940 16730 16952
rect 17126 16940 17132 16952
rect 17184 16940 17190 16992
rect 18046 16980 18052 16992
rect 18007 16952 18052 16980
rect 18046 16940 18052 16952
rect 18104 16940 18110 16992
rect 18414 16980 18420 16992
rect 18375 16952 18420 16980
rect 18414 16940 18420 16952
rect 18472 16940 18478 16992
rect 19242 16940 19248 16992
rect 19300 16980 19306 16992
rect 22186 16980 22192 16992
rect 19300 16952 22192 16980
rect 19300 16940 19306 16952
rect 22186 16940 22192 16952
rect 22244 16940 22250 16992
rect 23845 16983 23903 16989
rect 23845 16949 23857 16983
rect 23891 16980 23903 16983
rect 24486 16980 24492 16992
rect 23891 16952 24492 16980
rect 23891 16949 23903 16952
rect 23845 16943 23903 16949
rect 24486 16940 24492 16952
rect 24544 16940 24550 16992
rect 30742 16980 30748 16992
rect 30703 16952 30748 16980
rect 30742 16940 30748 16952
rect 30800 16940 30806 16992
rect 34606 16980 34612 16992
rect 34567 16952 34612 16980
rect 34606 16940 34612 16952
rect 34664 16940 34670 16992
rect 37642 16980 37648 16992
rect 37603 16952 37648 16980
rect 37642 16940 37648 16952
rect 37700 16940 37706 16992
rect 41785 16983 41843 16989
rect 41785 16949 41797 16983
rect 41831 16980 41843 16983
rect 42150 16980 42156 16992
rect 41831 16952 42156 16980
rect 41831 16949 41843 16952
rect 41785 16943 41843 16949
rect 42150 16940 42156 16952
rect 42208 16940 42214 16992
rect 1104 16890 42872 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 42872 16890
rect 1104 16816 42872 16838
rect 7650 16736 7656 16788
rect 7708 16776 7714 16788
rect 14366 16776 14372 16788
rect 7708 16748 14372 16776
rect 7708 16736 7714 16748
rect 14366 16736 14372 16748
rect 14424 16736 14430 16788
rect 14458 16736 14464 16788
rect 14516 16776 14522 16788
rect 14918 16776 14924 16788
rect 14516 16748 14924 16776
rect 14516 16736 14522 16748
rect 14918 16736 14924 16748
rect 14976 16776 14982 16788
rect 15102 16776 15108 16788
rect 14976 16748 15108 16776
rect 14976 16736 14982 16748
rect 15102 16736 15108 16748
rect 15160 16736 15166 16788
rect 16301 16779 16359 16785
rect 16301 16745 16313 16779
rect 16347 16776 16359 16779
rect 16482 16776 16488 16788
rect 16347 16748 16488 16776
rect 16347 16745 16359 16748
rect 16301 16739 16359 16745
rect 16482 16736 16488 16748
rect 16540 16736 16546 16788
rect 17865 16779 17923 16785
rect 17865 16776 17877 16779
rect 16929 16748 17877 16776
rect 13262 16668 13268 16720
rect 13320 16708 13326 16720
rect 15470 16708 15476 16720
rect 13320 16680 15476 16708
rect 13320 16668 13326 16680
rect 1854 16640 1860 16652
rect 1815 16612 1860 16640
rect 1854 16600 1860 16612
rect 1912 16600 1918 16652
rect 13541 16643 13599 16649
rect 13541 16609 13553 16643
rect 13587 16640 13599 16643
rect 13814 16640 13820 16652
rect 13587 16612 13820 16640
rect 13587 16609 13599 16612
rect 13541 16603 13599 16609
rect 13814 16600 13820 16612
rect 13872 16640 13878 16652
rect 14458 16640 14464 16652
rect 13872 16612 14464 16640
rect 13872 16600 13878 16612
rect 14458 16600 14464 16612
rect 14516 16600 14522 16652
rect 15212 16649 15240 16680
rect 15470 16668 15476 16680
rect 15528 16668 15534 16720
rect 16929 16708 16957 16748
rect 17865 16745 17877 16748
rect 17911 16776 17923 16779
rect 17911 16748 18083 16776
rect 17911 16745 17923 16748
rect 17865 16739 17923 16745
rect 15856 16680 16957 16708
rect 17773 16711 17831 16717
rect 15197 16643 15255 16649
rect 15197 16609 15209 16643
rect 15243 16609 15255 16643
rect 15197 16603 15255 16609
rect 1394 16572 1400 16584
rect 1355 16544 1400 16572
rect 1394 16532 1400 16544
rect 1452 16532 1458 16584
rect 13265 16575 13323 16581
rect 13265 16541 13277 16575
rect 13311 16572 13323 16575
rect 13354 16572 13360 16584
rect 13311 16544 13360 16572
rect 13311 16541 13323 16544
rect 13265 16535 13323 16541
rect 13354 16532 13360 16544
rect 13412 16532 13418 16584
rect 14274 16572 14280 16584
rect 14235 16544 14280 16572
rect 14274 16532 14280 16544
rect 14332 16532 14338 16584
rect 15102 16572 15108 16584
rect 15063 16544 15108 16572
rect 15102 16532 15108 16544
rect 15160 16572 15166 16584
rect 15856 16572 15884 16680
rect 17773 16677 17785 16711
rect 17819 16708 17831 16711
rect 17954 16708 17960 16720
rect 17819 16680 17960 16708
rect 17819 16677 17831 16680
rect 17773 16671 17831 16677
rect 17954 16668 17960 16680
rect 18012 16668 18018 16720
rect 18055 16708 18083 16748
rect 18414 16736 18420 16788
rect 18472 16776 18478 16788
rect 21177 16779 21235 16785
rect 21177 16776 21189 16779
rect 18472 16748 21189 16776
rect 18472 16736 18478 16748
rect 21177 16745 21189 16748
rect 21223 16745 21235 16779
rect 21358 16776 21364 16788
rect 21319 16748 21364 16776
rect 21177 16739 21235 16745
rect 21358 16736 21364 16748
rect 21416 16736 21422 16788
rect 23842 16736 23848 16788
rect 23900 16776 23906 16788
rect 24397 16779 24455 16785
rect 24397 16776 24409 16779
rect 23900 16748 24409 16776
rect 23900 16736 23906 16748
rect 24397 16745 24409 16748
rect 24443 16776 24455 16779
rect 24762 16776 24768 16788
rect 24443 16748 24768 16776
rect 24443 16745 24455 16748
rect 24397 16739 24455 16745
rect 24762 16736 24768 16748
rect 24820 16736 24826 16788
rect 27433 16779 27491 16785
rect 27433 16745 27445 16779
rect 27479 16776 27491 16779
rect 27706 16776 27712 16788
rect 27479 16748 27712 16776
rect 27479 16745 27491 16748
rect 27433 16739 27491 16745
rect 27706 16736 27712 16748
rect 27764 16736 27770 16788
rect 27798 16736 27804 16788
rect 27856 16776 27862 16788
rect 28077 16779 28135 16785
rect 28077 16776 28089 16779
rect 27856 16748 28089 16776
rect 27856 16736 27862 16748
rect 28077 16745 28089 16748
rect 28123 16776 28135 16779
rect 29362 16776 29368 16788
rect 28123 16748 29368 16776
rect 28123 16745 28135 16748
rect 28077 16739 28135 16745
rect 29362 16736 29368 16748
rect 29420 16736 29426 16788
rect 20809 16711 20867 16717
rect 20809 16708 20821 16711
rect 18055 16680 20821 16708
rect 16393 16643 16451 16649
rect 16393 16609 16405 16643
rect 16439 16640 16451 16643
rect 16942 16640 16948 16652
rect 16439 16612 16948 16640
rect 16439 16609 16451 16612
rect 16393 16603 16451 16609
rect 16942 16600 16948 16612
rect 17000 16640 17006 16652
rect 17221 16643 17279 16649
rect 17221 16640 17233 16643
rect 17000 16612 17233 16640
rect 17000 16600 17006 16612
rect 17221 16609 17233 16612
rect 17267 16609 17279 16643
rect 17678 16640 17684 16652
rect 17639 16612 17684 16640
rect 17221 16603 17279 16609
rect 17678 16600 17684 16612
rect 17736 16600 17742 16652
rect 15160 16544 15884 16572
rect 15160 16532 15166 16544
rect 15930 16532 15936 16584
rect 15988 16572 15994 16584
rect 16117 16575 16175 16581
rect 16117 16572 16129 16575
rect 15988 16544 16129 16572
rect 15988 16532 15994 16544
rect 16117 16541 16129 16544
rect 16163 16541 16175 16575
rect 16117 16535 16175 16541
rect 16574 16532 16580 16584
rect 16632 16572 16638 16584
rect 16853 16575 16911 16581
rect 16853 16572 16865 16575
rect 16632 16544 16865 16572
rect 16632 16532 16638 16544
rect 16853 16541 16865 16544
rect 16899 16541 16911 16575
rect 16853 16535 16911 16541
rect 17957 16575 18015 16581
rect 17957 16541 17969 16575
rect 18003 16572 18015 16575
rect 18046 16572 18052 16584
rect 18003 16544 18052 16572
rect 18003 16541 18015 16544
rect 17957 16535 18015 16541
rect 18046 16532 18052 16544
rect 18104 16572 18110 16584
rect 19242 16574 19248 16584
rect 19168 16572 19248 16574
rect 18104 16546 19248 16572
rect 18104 16544 19196 16546
rect 18104 16532 18110 16544
rect 19242 16532 19248 16546
rect 19300 16572 19306 16584
rect 19444 16581 19472 16680
rect 20809 16677 20821 16680
rect 20855 16708 20867 16711
rect 25777 16711 25835 16717
rect 20855 16680 22048 16708
rect 20855 16677 20867 16680
rect 20809 16671 20867 16677
rect 19889 16643 19947 16649
rect 19889 16640 19901 16643
rect 19536 16612 19901 16640
rect 19429 16575 19487 16581
rect 19300 16544 19345 16572
rect 19300 16532 19306 16544
rect 19429 16541 19441 16575
rect 19475 16541 19487 16575
rect 19429 16535 19487 16541
rect 1581 16507 1639 16513
rect 1581 16473 1593 16507
rect 1627 16504 1639 16507
rect 2130 16504 2136 16516
rect 1627 16476 2136 16504
rect 1627 16473 1639 16476
rect 1581 16467 1639 16473
rect 2130 16464 2136 16476
rect 2188 16464 2194 16516
rect 17034 16504 17040 16516
rect 16995 16476 17040 16504
rect 17034 16464 17040 16476
rect 17092 16464 17098 16516
rect 19337 16507 19395 16513
rect 19337 16473 19349 16507
rect 19383 16504 19395 16507
rect 19536 16504 19564 16612
rect 19889 16609 19901 16612
rect 19935 16609 19947 16643
rect 19889 16603 19947 16609
rect 20349 16643 20407 16649
rect 20349 16609 20361 16643
rect 20395 16640 20407 16643
rect 21174 16640 21180 16652
rect 20395 16612 21180 16640
rect 20395 16609 20407 16612
rect 20349 16603 20407 16609
rect 21174 16600 21180 16612
rect 21232 16600 21238 16652
rect 19981 16575 20039 16581
rect 19981 16541 19993 16575
rect 20027 16541 20039 16575
rect 19981 16535 20039 16541
rect 19383 16476 19564 16504
rect 19996 16504 20024 16535
rect 20070 16532 20076 16584
rect 20128 16572 20134 16584
rect 22020 16581 22048 16680
rect 25777 16677 25789 16711
rect 25823 16708 25835 16711
rect 26234 16708 26240 16720
rect 25823 16680 26240 16708
rect 25823 16677 25835 16680
rect 25777 16671 25835 16677
rect 26234 16668 26240 16680
rect 26292 16708 26298 16720
rect 31205 16711 31263 16717
rect 26292 16680 27568 16708
rect 26292 16668 26298 16680
rect 22186 16640 22192 16652
rect 22147 16612 22192 16640
rect 22186 16600 22192 16612
rect 22244 16600 22250 16652
rect 24486 16640 24492 16652
rect 24447 16612 24492 16640
rect 24486 16600 24492 16612
rect 24544 16640 24550 16652
rect 24544 16612 24808 16640
rect 24544 16600 24550 16612
rect 20165 16575 20223 16581
rect 20165 16572 20177 16575
rect 20128 16544 20177 16572
rect 20128 16532 20134 16544
rect 20165 16541 20177 16544
rect 20211 16541 20223 16575
rect 20165 16535 20223 16541
rect 22005 16575 22063 16581
rect 22005 16541 22017 16575
rect 22051 16541 22063 16575
rect 22005 16535 22063 16541
rect 23658 16532 23664 16584
rect 23716 16572 23722 16584
rect 24673 16575 24731 16581
rect 24673 16572 24685 16575
rect 23716 16544 24685 16572
rect 23716 16532 23722 16544
rect 24673 16541 24685 16544
rect 24719 16541 24731 16575
rect 24780 16572 24808 16612
rect 24854 16600 24860 16652
rect 24912 16640 24918 16652
rect 26421 16643 26479 16649
rect 26421 16640 26433 16643
rect 24912 16612 26433 16640
rect 24912 16600 24918 16612
rect 26421 16609 26433 16612
rect 26467 16609 26479 16643
rect 26421 16603 26479 16609
rect 25409 16575 25467 16581
rect 25409 16572 25421 16575
rect 24780 16544 25421 16572
rect 24673 16535 24731 16541
rect 25409 16541 25421 16544
rect 25455 16541 25467 16575
rect 25590 16572 25596 16584
rect 25551 16544 25596 16572
rect 25409 16535 25467 16541
rect 25590 16532 25596 16544
rect 25648 16532 25654 16584
rect 25777 16575 25835 16581
rect 25777 16541 25789 16575
rect 25823 16541 25835 16575
rect 25777 16535 25835 16541
rect 26605 16575 26663 16581
rect 26605 16541 26617 16575
rect 26651 16541 26663 16575
rect 26605 16535 26663 16541
rect 21821 16507 21879 16513
rect 21821 16504 21833 16507
rect 19996 16476 21833 16504
rect 19383 16473 19395 16476
rect 19337 16467 19395 16473
rect 21821 16473 21833 16476
rect 21867 16473 21879 16507
rect 21821 16467 21879 16473
rect 23750 16464 23756 16516
rect 23808 16504 23814 16516
rect 24397 16507 24455 16513
rect 24397 16504 24409 16507
rect 23808 16476 24409 16504
rect 23808 16464 23814 16476
rect 24397 16473 24409 16476
rect 24443 16504 24455 16507
rect 24443 16476 24716 16504
rect 24443 16473 24455 16476
rect 24397 16467 24455 16473
rect 24688 16448 24716 16476
rect 24762 16464 24768 16516
rect 24820 16504 24826 16516
rect 25792 16504 25820 16535
rect 26620 16504 26648 16535
rect 24820 16476 25820 16504
rect 25884 16476 26648 16504
rect 26789 16507 26847 16513
rect 24820 16464 24826 16476
rect 13538 16396 13544 16448
rect 13596 16436 13602 16448
rect 14093 16439 14151 16445
rect 14093 16436 14105 16439
rect 13596 16408 14105 16436
rect 13596 16396 13602 16408
rect 14093 16405 14105 16408
rect 14139 16405 14151 16439
rect 15470 16436 15476 16448
rect 15431 16408 15476 16436
rect 14093 16399 14151 16405
rect 15470 16396 15476 16408
rect 15528 16396 15534 16448
rect 15746 16396 15752 16448
rect 15804 16436 15810 16448
rect 15933 16439 15991 16445
rect 15933 16436 15945 16439
rect 15804 16408 15945 16436
rect 15804 16396 15810 16408
rect 15933 16405 15945 16408
rect 15979 16405 15991 16439
rect 15933 16399 15991 16405
rect 21177 16439 21235 16445
rect 21177 16405 21189 16439
rect 21223 16436 21235 16439
rect 21726 16436 21732 16448
rect 21223 16408 21732 16436
rect 21223 16405 21235 16408
rect 21177 16399 21235 16405
rect 21726 16396 21732 16408
rect 21784 16396 21790 16448
rect 24670 16396 24676 16448
rect 24728 16396 24734 16448
rect 24857 16439 24915 16445
rect 24857 16405 24869 16439
rect 24903 16436 24915 16439
rect 25130 16436 25136 16448
rect 24903 16408 25136 16436
rect 24903 16405 24915 16408
rect 24857 16399 24915 16405
rect 25130 16396 25136 16408
rect 25188 16436 25194 16448
rect 25884 16436 25912 16476
rect 26789 16473 26801 16507
rect 26835 16504 26847 16507
rect 27341 16507 27399 16513
rect 27341 16504 27353 16507
rect 26835 16476 27353 16504
rect 26835 16473 26847 16476
rect 26789 16467 26847 16473
rect 27341 16473 27353 16476
rect 27387 16473 27399 16507
rect 27540 16504 27568 16680
rect 31205 16677 31217 16711
rect 31251 16708 31263 16711
rect 32766 16708 32772 16720
rect 31251 16680 32772 16708
rect 31251 16677 31263 16680
rect 31205 16671 31263 16677
rect 32766 16668 32772 16680
rect 32824 16708 32830 16720
rect 33318 16708 33324 16720
rect 32824 16680 33324 16708
rect 32824 16668 32830 16680
rect 33318 16668 33324 16680
rect 33376 16708 33382 16720
rect 33873 16711 33931 16717
rect 33873 16708 33885 16711
rect 33376 16680 33885 16708
rect 33376 16668 33382 16680
rect 33873 16677 33885 16680
rect 33919 16677 33931 16711
rect 33873 16671 33931 16677
rect 34790 16600 34796 16652
rect 34848 16640 34854 16652
rect 41690 16640 41696 16652
rect 34848 16612 35020 16640
rect 41651 16612 41696 16640
rect 34848 16600 34854 16612
rect 28169 16575 28227 16581
rect 28169 16541 28181 16575
rect 28215 16572 28227 16575
rect 30098 16572 30104 16584
rect 28215 16544 30104 16572
rect 28215 16541 28227 16544
rect 28169 16535 28227 16541
rect 30098 16532 30104 16544
rect 30156 16532 30162 16584
rect 30742 16532 30748 16584
rect 30800 16572 30806 16584
rect 30837 16575 30895 16581
rect 30837 16572 30849 16575
rect 30800 16544 30849 16572
rect 30800 16532 30806 16544
rect 30837 16541 30849 16544
rect 30883 16541 30895 16575
rect 30837 16535 30895 16541
rect 30929 16575 30987 16581
rect 30929 16541 30941 16575
rect 30975 16541 30987 16575
rect 30929 16535 30987 16541
rect 30944 16504 30972 16535
rect 31018 16532 31024 16584
rect 31076 16572 31082 16584
rect 32488 16575 32546 16581
rect 31076 16544 31121 16572
rect 31076 16532 31082 16544
rect 32488 16541 32500 16575
rect 32534 16541 32546 16575
rect 32488 16535 32546 16541
rect 31110 16504 31116 16516
rect 27540 16476 31116 16504
rect 27341 16467 27399 16473
rect 31110 16464 31116 16476
rect 31168 16464 31174 16516
rect 32508 16504 32536 16535
rect 32582 16532 32588 16584
rect 32640 16572 32646 16584
rect 32858 16572 32864 16584
rect 32640 16544 32685 16572
rect 32819 16544 32864 16572
rect 32640 16532 32646 16544
rect 32858 16532 32864 16544
rect 32916 16532 32922 16584
rect 32950 16532 32956 16584
rect 33008 16572 33014 16584
rect 34992 16581 35020 16612
rect 41690 16600 41696 16612
rect 41748 16600 41754 16652
rect 42150 16640 42156 16652
rect 42111 16612 42156 16640
rect 42150 16600 42156 16612
rect 42208 16600 42214 16652
rect 33597 16575 33655 16581
rect 33597 16572 33609 16575
rect 33008 16544 33609 16572
rect 33008 16532 33014 16544
rect 33597 16541 33609 16544
rect 33643 16541 33655 16575
rect 33597 16535 33655 16541
rect 34977 16575 35035 16581
rect 34977 16541 34989 16575
rect 35023 16541 35035 16575
rect 34977 16535 35035 16541
rect 35161 16575 35219 16581
rect 35161 16541 35173 16575
rect 35207 16541 35219 16575
rect 37642 16572 37648 16584
rect 37603 16544 37648 16572
rect 35161 16535 35219 16541
rect 32677 16507 32735 16513
rect 32508 16476 32628 16504
rect 32600 16448 32628 16476
rect 32677 16473 32689 16507
rect 32723 16504 32735 16507
rect 32766 16504 32772 16516
rect 32723 16476 32772 16504
rect 32723 16473 32735 16476
rect 32677 16467 32735 16473
rect 32766 16464 32772 16476
rect 32824 16464 32830 16516
rect 32876 16504 32904 16532
rect 34606 16504 34612 16516
rect 32876 16476 34612 16504
rect 34606 16464 34612 16476
rect 34664 16504 34670 16516
rect 35176 16504 35204 16535
rect 37642 16532 37648 16544
rect 37700 16532 37706 16584
rect 35342 16504 35348 16516
rect 34664 16476 35348 16504
rect 34664 16464 34670 16476
rect 35342 16464 35348 16476
rect 35400 16464 35406 16516
rect 41414 16464 41420 16516
rect 41472 16504 41478 16516
rect 41969 16507 42027 16513
rect 41969 16504 41981 16507
rect 41472 16476 41981 16504
rect 41472 16464 41478 16476
rect 41969 16473 41981 16476
rect 42015 16473 42027 16507
rect 41969 16467 42027 16473
rect 25188 16408 25912 16436
rect 25188 16396 25194 16408
rect 26142 16396 26148 16448
rect 26200 16436 26206 16448
rect 31018 16436 31024 16448
rect 26200 16408 31024 16436
rect 26200 16396 26206 16408
rect 31018 16396 31024 16408
rect 31076 16396 31082 16448
rect 32306 16436 32312 16448
rect 32267 16408 32312 16436
rect 32306 16396 32312 16408
rect 32364 16396 32370 16448
rect 32582 16396 32588 16448
rect 32640 16396 32646 16448
rect 34057 16439 34115 16445
rect 34057 16405 34069 16439
rect 34103 16436 34115 16439
rect 34698 16436 34704 16448
rect 34103 16408 34704 16436
rect 34103 16405 34115 16408
rect 34057 16399 34115 16405
rect 34698 16396 34704 16408
rect 34756 16396 34762 16448
rect 34790 16396 34796 16448
rect 34848 16436 34854 16448
rect 35069 16439 35127 16445
rect 35069 16436 35081 16439
rect 34848 16408 35081 16436
rect 34848 16396 34854 16408
rect 35069 16405 35081 16408
rect 35115 16405 35127 16439
rect 35069 16399 35127 16405
rect 37274 16396 37280 16448
rect 37332 16436 37338 16448
rect 37461 16439 37519 16445
rect 37461 16436 37473 16439
rect 37332 16408 37473 16436
rect 37332 16396 37338 16408
rect 37461 16405 37473 16408
rect 37507 16405 37519 16439
rect 37461 16399 37519 16405
rect 1104 16346 42872 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 42872 16346
rect 1104 16272 42872 16294
rect 2130 16232 2136 16244
rect 2091 16204 2136 16232
rect 2130 16192 2136 16204
rect 2188 16192 2194 16244
rect 14752 16204 15148 16232
rect 13354 16164 13360 16176
rect 12820 16136 13360 16164
rect 1394 16096 1400 16108
rect 1355 16068 1400 16096
rect 1394 16056 1400 16068
rect 1452 16056 1458 16108
rect 2225 16099 2283 16105
rect 2225 16065 2237 16099
rect 2271 16096 2283 16099
rect 7098 16096 7104 16108
rect 2271 16068 7104 16096
rect 2271 16065 2283 16068
rect 2225 16059 2283 16065
rect 7098 16056 7104 16068
rect 7156 16056 7162 16108
rect 12820 16105 12848 16136
rect 13354 16124 13360 16136
rect 13412 16124 13418 16176
rect 14366 16124 14372 16176
rect 14424 16164 14430 16176
rect 14752 16173 14780 16204
rect 14737 16167 14795 16173
rect 14737 16164 14749 16167
rect 14424 16136 14749 16164
rect 14424 16124 14430 16136
rect 14737 16133 14749 16136
rect 14783 16133 14795 16167
rect 14737 16127 14795 16133
rect 14967 16133 15025 16139
rect 14967 16130 14979 16133
rect 12805 16099 12863 16105
rect 12805 16065 12817 16099
rect 12851 16065 12863 16099
rect 12805 16059 12863 16065
rect 12989 16099 13047 16105
rect 12989 16065 13001 16099
rect 13035 16096 13047 16099
rect 14274 16096 14280 16108
rect 13035 16068 14280 16096
rect 13035 16065 13047 16068
rect 12989 16059 13047 16065
rect 14274 16056 14280 16068
rect 14332 16096 14338 16108
rect 14952 16099 14979 16130
rect 15013 16099 15025 16133
rect 14952 16096 15025 16099
rect 14332 16093 15025 16096
rect 14332 16068 14980 16093
rect 14332 16056 14338 16068
rect 13262 15988 13268 16040
rect 13320 16028 13326 16040
rect 13449 16031 13507 16037
rect 13449 16028 13461 16031
rect 13320 16000 13461 16028
rect 13320 15988 13326 16000
rect 13449 15997 13461 16000
rect 13495 15997 13507 16031
rect 13449 15991 13507 15997
rect 13725 16031 13783 16037
rect 13725 15997 13737 16031
rect 13771 16028 13783 16031
rect 14366 16028 14372 16040
rect 13771 16000 14372 16028
rect 13771 15997 13783 16000
rect 13725 15991 13783 15997
rect 14366 15988 14372 16000
rect 14424 15988 14430 16040
rect 15120 16028 15148 16204
rect 15470 16192 15476 16244
rect 15528 16232 15534 16244
rect 18049 16235 18107 16241
rect 18049 16232 18061 16235
rect 15528 16204 18061 16232
rect 15528 16192 15534 16204
rect 18049 16201 18061 16204
rect 18095 16232 18107 16235
rect 18138 16232 18144 16244
rect 18095 16204 18144 16232
rect 18095 16201 18107 16204
rect 18049 16195 18107 16201
rect 18138 16192 18144 16204
rect 18196 16192 18202 16244
rect 20714 16232 20720 16244
rect 20675 16204 20720 16232
rect 20714 16192 20720 16204
rect 20772 16192 20778 16244
rect 41414 16232 41420 16244
rect 20824 16204 40908 16232
rect 41375 16204 41420 16232
rect 20824 16164 20852 16204
rect 17788 16136 20852 16164
rect 15746 16096 15752 16108
rect 15707 16068 15752 16096
rect 15746 16056 15752 16068
rect 15804 16056 15810 16108
rect 17678 16028 17684 16040
rect 15120 16000 17684 16028
rect 17678 15988 17684 16000
rect 17736 15988 17742 16040
rect 14458 15920 14464 15972
rect 14516 15960 14522 15972
rect 17788 15960 17816 16136
rect 21174 16124 21180 16176
rect 21232 16164 21238 16176
rect 22250 16167 22308 16173
rect 22250 16164 22262 16167
rect 21232 16136 22262 16164
rect 21232 16124 21238 16136
rect 22250 16133 22262 16136
rect 22296 16133 22308 16167
rect 22250 16127 22308 16133
rect 24596 16136 25268 16164
rect 17954 16096 17960 16108
rect 17915 16068 17960 16096
rect 17954 16056 17960 16068
rect 18012 16056 18018 16108
rect 18233 16099 18291 16105
rect 18233 16065 18245 16099
rect 18279 16096 18291 16099
rect 19593 16099 19651 16105
rect 19593 16096 19605 16099
rect 18279 16068 19605 16096
rect 18279 16065 18291 16068
rect 18233 16059 18291 16065
rect 19593 16065 19605 16068
rect 19639 16065 19651 16099
rect 19593 16059 19651 16065
rect 22005 16099 22063 16105
rect 22005 16065 22017 16099
rect 22051 16096 22063 16099
rect 22094 16096 22100 16108
rect 22051 16068 22100 16096
rect 22051 16065 22063 16068
rect 22005 16059 22063 16065
rect 22094 16056 22100 16068
rect 22152 16056 22158 16108
rect 23658 16056 23664 16108
rect 23716 16096 23722 16108
rect 24305 16099 24363 16105
rect 24305 16096 24317 16099
rect 23716 16068 24317 16096
rect 23716 16056 23722 16068
rect 24305 16065 24317 16068
rect 24351 16065 24363 16099
rect 24305 16059 24363 16065
rect 18417 16031 18475 16037
rect 18417 15997 18429 16031
rect 18463 15997 18475 16031
rect 19334 16028 19340 16040
rect 19295 16000 19340 16028
rect 18417 15991 18475 15997
rect 14516 15932 17816 15960
rect 14516 15920 14522 15932
rect 12989 15895 13047 15901
rect 12989 15861 13001 15895
rect 13035 15892 13047 15895
rect 13354 15892 13360 15904
rect 13035 15864 13360 15892
rect 13035 15861 13047 15864
rect 12989 15855 13047 15861
rect 13354 15852 13360 15864
rect 13412 15852 13418 15904
rect 14918 15892 14924 15904
rect 14879 15864 14924 15892
rect 14918 15852 14924 15864
rect 14976 15852 14982 15904
rect 15102 15892 15108 15904
rect 15063 15864 15108 15892
rect 15102 15852 15108 15864
rect 15160 15852 15166 15904
rect 15562 15852 15568 15904
rect 15620 15892 15626 15904
rect 15657 15895 15715 15901
rect 15657 15892 15669 15895
rect 15620 15864 15669 15892
rect 15620 15852 15626 15864
rect 15657 15861 15669 15864
rect 15703 15861 15715 15895
rect 18432 15892 18460 15991
rect 19334 15988 19340 16000
rect 19392 15988 19398 16040
rect 24320 16028 24348 16059
rect 24486 16056 24492 16108
rect 24544 16096 24550 16108
rect 24596 16105 24624 16136
rect 24581 16099 24639 16105
rect 24581 16096 24593 16099
rect 24544 16068 24593 16096
rect 24544 16056 24550 16068
rect 24581 16065 24593 16068
rect 24627 16065 24639 16099
rect 24581 16059 24639 16065
rect 24670 16056 24676 16108
rect 24728 16096 24734 16108
rect 25240 16105 25268 16136
rect 26142 16124 26148 16176
rect 26200 16164 26206 16176
rect 31018 16164 31024 16176
rect 26200 16136 26464 16164
rect 30979 16136 31024 16164
rect 26200 16124 26206 16136
rect 24765 16099 24823 16105
rect 24765 16096 24777 16099
rect 24728 16068 24777 16096
rect 24728 16056 24734 16068
rect 24765 16065 24777 16068
rect 24811 16065 24823 16099
rect 24765 16059 24823 16065
rect 25225 16099 25283 16105
rect 25225 16065 25237 16099
rect 25271 16065 25283 16099
rect 26234 16096 26240 16108
rect 26195 16068 26240 16096
rect 25225 16059 25283 16065
rect 26234 16056 26240 16068
rect 26292 16056 26298 16108
rect 26436 16105 26464 16136
rect 31018 16124 31024 16136
rect 31076 16124 31082 16176
rect 32217 16167 32275 16173
rect 32217 16133 32229 16167
rect 32263 16164 32275 16167
rect 32306 16164 32312 16176
rect 32263 16136 32312 16164
rect 32263 16133 32275 16136
rect 32217 16127 32275 16133
rect 32306 16124 32312 16136
rect 32364 16124 32370 16176
rect 32950 16164 32956 16176
rect 32416 16136 32956 16164
rect 26421 16099 26479 16105
rect 26421 16065 26433 16099
rect 26467 16065 26479 16099
rect 26421 16059 26479 16065
rect 26694 16056 26700 16108
rect 26752 16096 26758 16108
rect 26973 16099 27031 16105
rect 26973 16096 26985 16099
rect 26752 16068 26985 16096
rect 26752 16056 26758 16068
rect 26973 16065 26985 16068
rect 27019 16065 27031 16099
rect 27229 16099 27287 16105
rect 27229 16096 27241 16099
rect 26973 16059 27031 16065
rect 27080 16068 27241 16096
rect 25317 16031 25375 16037
rect 25317 16028 25329 16031
rect 24320 16000 25329 16028
rect 25317 15997 25329 16000
rect 25363 16028 25375 16031
rect 25590 16028 25596 16040
rect 25363 16000 25596 16028
rect 25363 15997 25375 16000
rect 25317 15991 25375 15997
rect 25590 15988 25596 16000
rect 25648 15988 25654 16040
rect 26329 16031 26387 16037
rect 26329 15997 26341 16031
rect 26375 16028 26387 16031
rect 27080 16028 27108 16068
rect 27229 16065 27241 16068
rect 27275 16065 27287 16099
rect 29089 16099 29147 16105
rect 29089 16096 29101 16099
rect 27229 16059 27287 16065
rect 28368 16068 29101 16096
rect 26375 16000 27108 16028
rect 26375 15997 26387 16000
rect 26329 15991 26387 15997
rect 23385 15963 23443 15969
rect 23385 15929 23397 15963
rect 23431 15960 23443 15963
rect 23750 15960 23756 15972
rect 23431 15932 23756 15960
rect 23431 15929 23443 15932
rect 23385 15923 23443 15929
rect 23750 15920 23756 15932
rect 23808 15920 23814 15972
rect 24762 15920 24768 15972
rect 24820 15960 24826 15972
rect 28368 15969 28396 16068
rect 29089 16065 29101 16068
rect 29135 16065 29147 16099
rect 29089 16059 29147 16065
rect 30653 16099 30711 16105
rect 30653 16065 30665 16099
rect 30699 16096 30711 16099
rect 30742 16096 30748 16108
rect 30699 16068 30748 16096
rect 30699 16065 30711 16068
rect 30653 16059 30711 16065
rect 30742 16056 30748 16068
rect 30800 16056 30806 16108
rect 31110 16056 31116 16108
rect 31168 16096 31174 16108
rect 32416 16096 32444 16136
rect 32950 16124 32956 16136
rect 33008 16124 33014 16176
rect 32582 16096 32588 16108
rect 31168 16068 31213 16096
rect 31726 16068 32444 16096
rect 32543 16068 32588 16096
rect 31168 16056 31174 16068
rect 28810 16028 28816 16040
rect 28771 16000 28816 16028
rect 28810 15988 28816 16000
rect 28868 15988 28874 16040
rect 28994 16028 29000 16040
rect 28955 16000 29000 16028
rect 28994 15988 29000 16000
rect 29052 15988 29058 16040
rect 30837 16031 30895 16037
rect 30837 15997 30849 16031
rect 30883 16028 30895 16031
rect 31726 16028 31754 16068
rect 32582 16056 32588 16068
rect 32640 16056 32646 16108
rect 33413 16099 33471 16105
rect 33413 16096 33425 16099
rect 32692 16068 33425 16096
rect 32692 16040 32720 16068
rect 33413 16065 33425 16068
rect 33459 16065 33471 16099
rect 33413 16059 33471 16065
rect 33686 16056 33692 16108
rect 33744 16096 33750 16108
rect 34425 16099 34483 16105
rect 34425 16096 34437 16099
rect 33744 16068 34437 16096
rect 33744 16056 33750 16068
rect 34425 16065 34437 16068
rect 34471 16065 34483 16099
rect 34425 16059 34483 16065
rect 34698 16056 34704 16108
rect 34756 16096 34762 16108
rect 35437 16099 35495 16105
rect 35437 16096 35449 16099
rect 34756 16068 35449 16096
rect 34756 16056 34762 16068
rect 35437 16065 35449 16068
rect 35483 16065 35495 16099
rect 37274 16096 37280 16108
rect 37235 16068 37280 16096
rect 35437 16059 35495 16065
rect 37274 16056 37280 16068
rect 37332 16056 37338 16108
rect 40880 16105 40908 16204
rect 41414 16192 41420 16204
rect 41472 16192 41478 16244
rect 40865 16099 40923 16105
rect 40865 16065 40877 16099
rect 40911 16065 40923 16099
rect 40865 16059 40923 16065
rect 32674 16028 32680 16040
rect 30883 16000 31754 16028
rect 32635 16000 32680 16028
rect 30883 15997 30895 16000
rect 30837 15991 30895 15997
rect 32674 15988 32680 16000
rect 32732 15988 32738 16040
rect 33321 16031 33379 16037
rect 33321 15997 33333 16031
rect 33367 15997 33379 16031
rect 33321 15991 33379 15997
rect 33781 16031 33839 16037
rect 33781 15997 33793 16031
rect 33827 16028 33839 16031
rect 34333 16031 34391 16037
rect 34333 16028 34345 16031
rect 33827 16000 34345 16028
rect 33827 15997 33839 16000
rect 33781 15991 33839 15997
rect 34333 15997 34345 16000
rect 34379 15997 34391 16031
rect 35342 16028 35348 16040
rect 35303 16000 35348 16028
rect 34333 15991 34391 15997
rect 28353 15963 28411 15969
rect 24820 15932 25268 15960
rect 24820 15920 24826 15932
rect 21818 15892 21824 15904
rect 18432 15864 21824 15892
rect 15657 15855 15715 15861
rect 21818 15852 21824 15864
rect 21876 15852 21882 15904
rect 24443 15895 24501 15901
rect 24443 15861 24455 15895
rect 24489 15892 24501 15895
rect 24578 15892 24584 15904
rect 24489 15864 24584 15892
rect 24489 15861 24501 15864
rect 24443 15855 24501 15861
rect 24578 15852 24584 15864
rect 24636 15852 24642 15904
rect 24673 15895 24731 15901
rect 24673 15861 24685 15895
rect 24719 15892 24731 15895
rect 24854 15892 24860 15904
rect 24719 15864 24860 15892
rect 24719 15861 24731 15864
rect 24673 15855 24731 15861
rect 24854 15852 24860 15864
rect 24912 15852 24918 15904
rect 25240 15901 25268 15932
rect 28353 15929 28365 15963
rect 28399 15929 28411 15963
rect 28353 15923 28411 15929
rect 32582 15920 32588 15972
rect 32640 15960 32646 15972
rect 33336 15960 33364 15991
rect 35342 15988 35348 16000
rect 35400 15988 35406 16040
rect 37458 16028 37464 16040
rect 37419 16000 37464 16028
rect 37458 15988 37464 16000
rect 37516 15988 37522 16040
rect 38930 16028 38936 16040
rect 38891 16000 38936 16028
rect 38930 15988 38936 16000
rect 38988 15988 38994 16040
rect 40880 16028 40908 16059
rect 40954 16056 40960 16108
rect 41012 16096 41018 16108
rect 41325 16099 41383 16105
rect 41325 16096 41337 16099
rect 41012 16068 41337 16096
rect 41012 16056 41018 16068
rect 41325 16065 41337 16068
rect 41371 16096 41383 16099
rect 42334 16096 42340 16108
rect 41371 16068 42340 16096
rect 41371 16065 41383 16068
rect 41325 16059 41383 16065
rect 42334 16056 42340 16068
rect 42392 16056 42398 16108
rect 41874 16028 41880 16040
rect 40880 16000 41880 16028
rect 41874 15988 41880 16000
rect 41932 15988 41938 16040
rect 32640 15932 33364 15960
rect 32640 15920 32646 15932
rect 25225 15895 25283 15901
rect 25225 15861 25237 15895
rect 25271 15861 25283 15895
rect 25590 15892 25596 15904
rect 25503 15864 25596 15892
rect 25225 15855 25283 15861
rect 25590 15852 25596 15864
rect 25648 15892 25654 15904
rect 26142 15892 26148 15904
rect 25648 15864 26148 15892
rect 25648 15852 25654 15864
rect 26142 15852 26148 15864
rect 26200 15852 26206 15904
rect 28902 15892 28908 15904
rect 28863 15864 28908 15892
rect 28902 15852 28908 15864
rect 28960 15852 28966 15904
rect 32030 15852 32036 15904
rect 32088 15892 32094 15904
rect 32309 15895 32367 15901
rect 32309 15892 32321 15895
rect 32088 15864 32321 15892
rect 32088 15852 32094 15864
rect 32309 15861 32321 15864
rect 32355 15861 32367 15895
rect 32309 15855 32367 15861
rect 34606 15852 34612 15904
rect 34664 15892 34670 15904
rect 34701 15895 34759 15901
rect 34701 15892 34713 15895
rect 34664 15864 34713 15892
rect 34664 15852 34670 15864
rect 34701 15861 34713 15864
rect 34747 15861 34759 15895
rect 34701 15855 34759 15861
rect 35805 15895 35863 15901
rect 35805 15861 35817 15895
rect 35851 15892 35863 15895
rect 36078 15892 36084 15904
rect 35851 15864 36084 15892
rect 35851 15861 35863 15864
rect 35805 15855 35863 15861
rect 36078 15852 36084 15864
rect 36136 15852 36142 15904
rect 40221 15895 40279 15901
rect 40221 15861 40233 15895
rect 40267 15892 40279 15895
rect 40310 15892 40316 15904
rect 40267 15864 40316 15892
rect 40267 15861 40279 15864
rect 40221 15855 40279 15861
rect 40310 15852 40316 15864
rect 40368 15852 40374 15904
rect 40494 15852 40500 15904
rect 40552 15892 40558 15904
rect 40773 15895 40831 15901
rect 40773 15892 40785 15895
rect 40552 15864 40785 15892
rect 40552 15852 40558 15864
rect 40773 15861 40785 15864
rect 40819 15861 40831 15895
rect 40773 15855 40831 15861
rect 1104 15802 42872 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 42872 15802
rect 1104 15728 42872 15750
rect 11517 15691 11575 15697
rect 11517 15657 11529 15691
rect 11563 15688 11575 15691
rect 13262 15688 13268 15700
rect 11563 15660 13268 15688
rect 11563 15657 11575 15660
rect 11517 15651 11575 15657
rect 13262 15648 13268 15660
rect 13320 15648 13326 15700
rect 13446 15648 13452 15700
rect 13504 15688 13510 15700
rect 13541 15691 13599 15697
rect 13541 15688 13553 15691
rect 13504 15660 13553 15688
rect 13504 15648 13510 15660
rect 13541 15657 13553 15660
rect 13587 15657 13599 15691
rect 13541 15651 13599 15657
rect 15102 15648 15108 15700
rect 15160 15688 15166 15700
rect 18138 15688 18144 15700
rect 15160 15660 15516 15688
rect 18099 15660 18144 15688
rect 15160 15648 15166 15660
rect 13630 15580 13636 15632
rect 13688 15620 13694 15632
rect 14274 15620 14280 15632
rect 13688 15592 14280 15620
rect 13688 15580 13694 15592
rect 14274 15580 14280 15592
rect 14332 15580 14338 15632
rect 12897 15555 12955 15561
rect 12897 15521 12909 15555
rect 12943 15552 12955 15555
rect 13998 15552 14004 15564
rect 12943 15524 14004 15552
rect 12943 15521 12955 15524
rect 12897 15515 12955 15521
rect 13998 15512 14004 15524
rect 14056 15512 14062 15564
rect 15378 15552 15384 15564
rect 15339 15524 15384 15552
rect 15378 15512 15384 15524
rect 15436 15512 15442 15564
rect 15488 15561 15516 15660
rect 18138 15648 18144 15660
rect 18196 15648 18202 15700
rect 21637 15691 21695 15697
rect 21637 15657 21649 15691
rect 21683 15688 21695 15691
rect 22462 15688 22468 15700
rect 21683 15660 22468 15688
rect 21683 15657 21695 15660
rect 21637 15651 21695 15657
rect 22462 15648 22468 15660
rect 22520 15648 22526 15700
rect 28442 15688 28448 15700
rect 27448 15660 28448 15688
rect 15473 15555 15531 15561
rect 15473 15521 15485 15555
rect 15519 15521 15531 15555
rect 16114 15552 16120 15564
rect 16075 15524 16120 15552
rect 15473 15515 15531 15521
rect 16114 15512 16120 15524
rect 16172 15512 16178 15564
rect 18156 15552 18184 15648
rect 21726 15580 21732 15632
rect 21784 15620 21790 15632
rect 27448 15620 27476 15660
rect 28442 15648 28448 15660
rect 28500 15648 28506 15700
rect 28810 15688 28816 15700
rect 28771 15660 28816 15688
rect 28810 15648 28816 15660
rect 28868 15648 28874 15700
rect 32582 15688 32588 15700
rect 28920 15660 32588 15688
rect 21784 15592 27476 15620
rect 21784 15580 21790 15592
rect 19426 15552 19432 15564
rect 17604 15524 19432 15552
rect 1762 15484 1768 15496
rect 1723 15456 1768 15484
rect 1762 15444 1768 15456
rect 1820 15444 1826 15496
rect 13354 15484 13360 15496
rect 13315 15456 13360 15484
rect 13354 15444 13360 15456
rect 13412 15444 13418 15496
rect 13538 15484 13544 15496
rect 13499 15456 13544 15484
rect 13538 15444 13544 15456
rect 13596 15444 13602 15496
rect 13814 15444 13820 15496
rect 13872 15484 13878 15496
rect 14093 15487 14151 15493
rect 14093 15484 14105 15487
rect 13872 15456 14105 15484
rect 13872 15444 13878 15456
rect 14093 15453 14105 15456
rect 14139 15453 14151 15487
rect 14366 15484 14372 15496
rect 14093 15447 14151 15453
rect 14200 15456 14372 15484
rect 12652 15419 12710 15425
rect 12652 15385 12664 15419
rect 12698 15416 12710 15419
rect 13170 15416 13176 15428
rect 12698 15388 13176 15416
rect 12698 15385 12710 15388
rect 12652 15379 12710 15385
rect 13170 15376 13176 15388
rect 13228 15376 13234 15428
rect 13446 15376 13452 15428
rect 13504 15416 13510 15428
rect 14200 15416 14228 15456
rect 14366 15444 14372 15456
rect 14424 15444 14430 15496
rect 14461 15487 14519 15493
rect 14461 15453 14473 15487
rect 14507 15484 14519 15487
rect 15194 15484 15200 15496
rect 14507 15456 15056 15484
rect 15155 15456 15200 15484
rect 14507 15453 14519 15456
rect 14461 15447 14519 15453
rect 13504 15388 14228 15416
rect 13504 15376 13510 15388
rect 14274 15376 14280 15428
rect 14332 15416 14338 15428
rect 14332 15388 14377 15416
rect 14332 15376 14338 15388
rect 7098 15308 7104 15360
rect 7156 15348 7162 15360
rect 7558 15348 7564 15360
rect 7156 15320 7564 15348
rect 7156 15308 7162 15320
rect 7558 15308 7564 15320
rect 7616 15308 7622 15360
rect 11146 15308 11152 15360
rect 11204 15348 11210 15360
rect 12066 15348 12072 15360
rect 11204 15320 12072 15348
rect 11204 15308 11210 15320
rect 12066 15308 12072 15320
rect 12124 15348 12130 15360
rect 14458 15348 14464 15360
rect 12124 15320 14464 15348
rect 12124 15308 12130 15320
rect 14458 15308 14464 15320
rect 14516 15308 14522 15360
rect 14642 15348 14648 15360
rect 14603 15320 14648 15348
rect 14642 15308 14648 15320
rect 14700 15308 14706 15360
rect 15028 15348 15056 15456
rect 15194 15444 15200 15456
rect 15252 15444 15258 15496
rect 15289 15487 15347 15493
rect 15289 15453 15301 15487
rect 15335 15484 15347 15487
rect 15654 15484 15660 15496
rect 15335 15456 15660 15484
rect 15335 15453 15347 15456
rect 15289 15447 15347 15453
rect 15654 15444 15660 15456
rect 15712 15444 15718 15496
rect 15746 15444 15752 15496
rect 15804 15484 15810 15496
rect 16209 15487 16267 15493
rect 16209 15484 16221 15487
rect 15804 15456 16221 15484
rect 15804 15444 15810 15456
rect 16209 15453 16221 15456
rect 16255 15453 16267 15487
rect 16390 15484 16396 15496
rect 16351 15456 16396 15484
rect 16209 15447 16267 15453
rect 16390 15444 16396 15456
rect 16448 15444 16454 15496
rect 17034 15444 17040 15496
rect 17092 15484 17098 15496
rect 17402 15484 17408 15496
rect 17092 15456 17408 15484
rect 17092 15444 17098 15456
rect 17402 15444 17408 15456
rect 17460 15444 17466 15496
rect 17604 15493 17632 15524
rect 19426 15512 19432 15524
rect 19484 15512 19490 15564
rect 20714 15512 20720 15564
rect 20772 15552 20778 15564
rect 20772 15524 22094 15552
rect 20772 15512 20778 15524
rect 17589 15487 17647 15493
rect 17589 15453 17601 15487
rect 17635 15453 17647 15487
rect 18046 15484 18052 15496
rect 18007 15456 18052 15484
rect 17589 15447 17647 15453
rect 18046 15444 18052 15456
rect 18104 15444 18110 15496
rect 18322 15484 18328 15496
rect 18283 15456 18328 15484
rect 18322 15444 18328 15456
rect 18380 15444 18386 15496
rect 20806 15484 20812 15496
rect 20767 15456 20812 15484
rect 20806 15444 20812 15456
rect 20864 15444 20870 15496
rect 21358 15484 21364 15496
rect 21319 15456 21364 15484
rect 21358 15444 21364 15456
rect 21416 15444 21422 15496
rect 21818 15484 21824 15496
rect 21779 15456 21824 15484
rect 21818 15444 21824 15456
rect 21876 15444 21882 15496
rect 22066 15484 22094 15524
rect 24854 15512 24860 15564
rect 24912 15552 24918 15564
rect 24949 15555 25007 15561
rect 24949 15552 24961 15555
rect 24912 15524 24961 15552
rect 24912 15512 24918 15524
rect 24949 15521 24961 15524
rect 24995 15521 25007 15555
rect 24949 15515 25007 15521
rect 24762 15484 24768 15496
rect 22066 15456 24768 15484
rect 24762 15444 24768 15456
rect 24820 15484 24826 15496
rect 25041 15487 25099 15493
rect 25041 15484 25053 15487
rect 24820 15456 25053 15484
rect 24820 15444 24826 15456
rect 25041 15453 25053 15456
rect 25087 15453 25099 15487
rect 25041 15447 25099 15453
rect 26694 15444 26700 15496
rect 26752 15484 26758 15496
rect 27706 15493 27712 15496
rect 27433 15487 27491 15493
rect 27433 15484 27445 15487
rect 26752 15456 27445 15484
rect 26752 15444 26758 15456
rect 27433 15453 27445 15456
rect 27479 15453 27491 15487
rect 27700 15484 27712 15493
rect 27619 15456 27712 15484
rect 27433 15447 27491 15453
rect 27700 15447 27712 15456
rect 27764 15484 27770 15496
rect 28920 15484 28948 15660
rect 32582 15648 32588 15660
rect 32640 15648 32646 15700
rect 33686 15688 33692 15700
rect 33647 15660 33692 15688
rect 33686 15648 33692 15660
rect 33744 15648 33750 15700
rect 37277 15691 37335 15697
rect 37277 15657 37289 15691
rect 37323 15688 37335 15691
rect 37458 15688 37464 15700
rect 37323 15660 37464 15688
rect 37323 15657 37335 15660
rect 37277 15651 37335 15657
rect 37458 15648 37464 15660
rect 37516 15648 37522 15700
rect 34790 15580 34796 15632
rect 34848 15620 34854 15632
rect 34977 15623 35035 15629
rect 34977 15620 34989 15623
rect 34848 15592 34989 15620
rect 34848 15580 34854 15592
rect 34977 15589 34989 15592
rect 35023 15620 35035 15623
rect 35526 15620 35532 15632
rect 35023 15592 35532 15620
rect 35023 15589 35035 15592
rect 34977 15583 35035 15589
rect 35526 15580 35532 15592
rect 35584 15620 35590 15632
rect 41506 15620 41512 15632
rect 35584 15592 35664 15620
rect 35584 15580 35590 15592
rect 29362 15512 29368 15564
rect 29420 15552 29426 15564
rect 29549 15555 29607 15561
rect 29549 15552 29561 15555
rect 29420 15524 29561 15552
rect 29420 15512 29426 15524
rect 29549 15521 29561 15524
rect 29595 15521 29607 15555
rect 29549 15515 29607 15521
rect 32950 15512 32956 15564
rect 33008 15552 33014 15564
rect 34698 15552 34704 15564
rect 33008 15524 33548 15552
rect 34659 15524 34704 15552
rect 33008 15512 33014 15524
rect 27764 15456 28948 15484
rect 27706 15444 27712 15447
rect 27764 15444 27770 15456
rect 29638 15444 29644 15496
rect 29696 15484 29702 15496
rect 29805 15487 29863 15493
rect 29805 15484 29817 15487
rect 29696 15456 29817 15484
rect 29696 15444 29702 15456
rect 29805 15453 29817 15456
rect 29851 15453 29863 15487
rect 29805 15447 29863 15453
rect 32858 15444 32864 15496
rect 32916 15484 32922 15496
rect 33229 15487 33287 15493
rect 33229 15484 33241 15487
rect 32916 15456 33241 15484
rect 32916 15444 32922 15456
rect 33229 15453 33241 15456
rect 33275 15453 33287 15487
rect 33229 15447 33287 15453
rect 33318 15444 33324 15496
rect 33376 15484 33382 15496
rect 33520 15493 33548 15524
rect 34698 15512 34704 15524
rect 34756 15512 34762 15564
rect 35636 15561 35664 15592
rect 37200 15592 41512 15620
rect 35621 15555 35679 15561
rect 35621 15521 35633 15555
rect 35667 15521 35679 15555
rect 35621 15515 35679 15521
rect 33505 15487 33563 15493
rect 33376 15456 33421 15484
rect 33376 15444 33382 15456
rect 33505 15453 33517 15487
rect 33551 15453 33563 15487
rect 35894 15484 35900 15496
rect 35855 15456 35900 15484
rect 33505 15447 33563 15453
rect 35894 15444 35900 15456
rect 35952 15444 35958 15496
rect 36538 15444 36544 15496
rect 36596 15484 36602 15496
rect 37200 15493 37228 15592
rect 41506 15580 41512 15592
rect 41564 15580 41570 15632
rect 40310 15552 40316 15564
rect 40271 15524 40316 15552
rect 40310 15512 40316 15524
rect 40368 15512 40374 15564
rect 40494 15552 40500 15564
rect 40455 15524 40500 15552
rect 40494 15512 40500 15524
rect 40552 15512 40558 15564
rect 42150 15552 42156 15564
rect 42111 15524 42156 15552
rect 42150 15512 42156 15524
rect 42208 15512 42214 15564
rect 37185 15487 37243 15493
rect 37185 15484 37197 15487
rect 36596 15456 37197 15484
rect 36596 15444 36602 15456
rect 37185 15453 37197 15456
rect 37231 15453 37243 15487
rect 37185 15447 37243 15453
rect 16408 15416 16436 15444
rect 15304 15388 16436 15416
rect 15304 15348 15332 15388
rect 19334 15376 19340 15428
rect 19392 15416 19398 15428
rect 19613 15419 19671 15425
rect 19613 15416 19625 15419
rect 19392 15388 19625 15416
rect 19392 15376 19398 15388
rect 19613 15385 19625 15388
rect 19659 15385 19671 15419
rect 19613 15379 19671 15385
rect 19797 15419 19855 15425
rect 19797 15385 19809 15419
rect 19843 15416 19855 15419
rect 20625 15419 20683 15425
rect 20625 15416 20637 15419
rect 19843 15388 20637 15416
rect 19843 15385 19855 15388
rect 19797 15379 19855 15385
rect 20625 15385 20637 15388
rect 20671 15416 20683 15419
rect 20714 15416 20720 15428
rect 20671 15388 20720 15416
rect 20671 15385 20683 15388
rect 20625 15379 20683 15385
rect 20714 15376 20720 15388
rect 20772 15376 20778 15428
rect 21453 15419 21511 15425
rect 21453 15385 21465 15419
rect 21499 15416 21511 15419
rect 22646 15416 22652 15428
rect 21499 15388 22652 15416
rect 21499 15385 21511 15388
rect 21453 15379 21511 15385
rect 22646 15376 22652 15388
rect 22704 15376 22710 15428
rect 15028 15320 15332 15348
rect 15470 15308 15476 15360
rect 15528 15348 15534 15360
rect 15657 15351 15715 15357
rect 15657 15348 15669 15351
rect 15528 15320 15669 15348
rect 15528 15308 15534 15320
rect 15657 15317 15669 15320
rect 15703 15317 15715 15351
rect 15657 15311 15715 15317
rect 17497 15351 17555 15357
rect 17497 15317 17509 15351
rect 17543 15348 17555 15351
rect 18414 15348 18420 15360
rect 17543 15320 18420 15348
rect 17543 15317 17555 15320
rect 17497 15311 17555 15317
rect 18414 15308 18420 15320
rect 18472 15308 18478 15360
rect 18509 15351 18567 15357
rect 18509 15317 18521 15351
rect 18555 15348 18567 15351
rect 20530 15348 20536 15360
rect 18555 15320 20536 15348
rect 18555 15317 18567 15320
rect 18509 15311 18567 15317
rect 20530 15308 20536 15320
rect 20588 15308 20594 15360
rect 25409 15351 25467 15357
rect 25409 15317 25421 15351
rect 25455 15348 25467 15351
rect 26878 15348 26884 15360
rect 25455 15320 26884 15348
rect 25455 15317 25467 15320
rect 25409 15311 25467 15317
rect 26878 15308 26884 15320
rect 26936 15308 26942 15360
rect 30926 15348 30932 15360
rect 30887 15320 30932 15348
rect 30926 15308 30932 15320
rect 30984 15308 30990 15360
rect 35161 15351 35219 15357
rect 35161 15317 35173 15351
rect 35207 15348 35219 15351
rect 35342 15348 35348 15360
rect 35207 15320 35348 15348
rect 35207 15317 35219 15320
rect 35161 15311 35219 15317
rect 35342 15308 35348 15320
rect 35400 15308 35406 15360
rect 1104 15258 42872 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 42872 15258
rect 1104 15184 42872 15206
rect 13170 15144 13176 15156
rect 13131 15116 13176 15144
rect 13170 15104 13176 15116
rect 13228 15104 13234 15156
rect 13538 15104 13544 15156
rect 13596 15104 13602 15156
rect 15010 15104 15016 15156
rect 15068 15144 15074 15156
rect 15068 15116 17080 15144
rect 15068 15104 15074 15116
rect 13556 15023 13584 15104
rect 14642 15076 14648 15088
rect 13648 15048 14648 15076
rect 1762 15008 1768 15020
rect 1723 14980 1768 15008
rect 1762 14968 1768 14980
rect 1820 14968 1826 15020
rect 13446 15008 13452 15020
rect 13407 14980 13452 15008
rect 13446 14968 13452 14980
rect 13504 14968 13510 15020
rect 13538 15017 13596 15023
rect 13648 15017 13676 15048
rect 14642 15036 14648 15048
rect 14700 15036 14706 15088
rect 14737 15079 14795 15085
rect 14737 15045 14749 15079
rect 14783 15076 14795 15079
rect 15194 15076 15200 15088
rect 14783 15048 15200 15076
rect 14783 15045 14795 15048
rect 14737 15039 14795 15045
rect 15194 15036 15200 15048
rect 15252 15036 15258 15088
rect 13538 14983 13550 15017
rect 13584 14983 13596 15017
rect 13538 14977 13596 14983
rect 13633 15011 13691 15017
rect 13633 14977 13645 15011
rect 13679 14977 13691 15011
rect 13633 14971 13691 14977
rect 13817 15011 13875 15017
rect 13817 14977 13829 15011
rect 13863 15008 13875 15011
rect 14182 15008 14188 15020
rect 13863 14980 14188 15008
rect 13863 14977 13875 14980
rect 13817 14971 13875 14977
rect 14182 14968 14188 14980
rect 14240 14968 14246 15020
rect 14274 14968 14280 15020
rect 14332 15008 14338 15020
rect 14369 15011 14427 15017
rect 14369 15008 14381 15011
rect 14332 14980 14381 15008
rect 14332 14968 14338 14980
rect 14369 14977 14381 14980
rect 14415 14977 14427 15011
rect 14369 14971 14427 14977
rect 14829 15011 14887 15017
rect 14829 14977 14841 15011
rect 14875 15008 14887 15011
rect 15102 15008 15108 15020
rect 14875 14980 15108 15008
rect 14875 14977 14887 14980
rect 14829 14971 14887 14977
rect 15102 14968 15108 14980
rect 15160 14968 15166 15020
rect 15304 15017 15332 15116
rect 15933 15079 15991 15085
rect 15933 15045 15945 15079
rect 15979 15076 15991 15079
rect 16914 15079 16972 15085
rect 16914 15076 16926 15079
rect 15979 15048 16926 15076
rect 15979 15045 15991 15048
rect 15933 15039 15991 15045
rect 16914 15045 16926 15048
rect 16960 15045 16972 15079
rect 17052 15076 17080 15116
rect 17402 15104 17408 15156
rect 17460 15144 17466 15156
rect 18049 15147 18107 15153
rect 18049 15144 18061 15147
rect 17460 15116 18061 15144
rect 17460 15104 17466 15116
rect 18049 15113 18061 15116
rect 18095 15113 18107 15147
rect 18049 15107 18107 15113
rect 24975 15147 25033 15153
rect 24975 15113 24987 15147
rect 25021 15144 25033 15147
rect 25590 15144 25596 15156
rect 25021 15116 25596 15144
rect 25021 15113 25033 15116
rect 24975 15107 25033 15113
rect 25590 15104 25596 15116
rect 25648 15104 25654 15156
rect 19058 15076 19064 15088
rect 17052 15048 19064 15076
rect 16914 15039 16972 15045
rect 19058 15036 19064 15048
rect 19116 15036 19122 15088
rect 20438 15076 20444 15088
rect 20088 15048 20444 15076
rect 20088 15020 20116 15048
rect 20438 15036 20444 15048
rect 20496 15076 20502 15088
rect 22738 15076 22744 15088
rect 20496 15048 20944 15076
rect 22699 15048 22744 15076
rect 20496 15036 20502 15048
rect 15289 15011 15347 15017
rect 15289 14977 15301 15011
rect 15335 14977 15347 15011
rect 15470 15008 15476 15020
rect 15431 14980 15476 15008
rect 15289 14971 15347 14977
rect 15470 14968 15476 14980
rect 15528 14968 15534 15020
rect 15565 15011 15623 15017
rect 15565 14977 15577 15011
rect 15611 14977 15623 15011
rect 15565 14971 15623 14977
rect 15657 15011 15715 15017
rect 15657 14977 15669 15011
rect 15703 15008 15715 15011
rect 16390 15008 16396 15020
rect 15703 14980 16396 15008
rect 15703 14977 15715 14980
rect 15657 14971 15715 14977
rect 1949 14943 2007 14949
rect 1949 14909 1961 14943
rect 1995 14940 2007 14943
rect 2222 14940 2228 14952
rect 1995 14912 2228 14940
rect 1995 14909 2007 14912
rect 1949 14903 2007 14909
rect 2222 14900 2228 14912
rect 2280 14900 2286 14952
rect 2774 14940 2780 14952
rect 2735 14912 2780 14940
rect 2774 14900 2780 14912
rect 2832 14900 2838 14952
rect 14553 14943 14611 14949
rect 14553 14909 14565 14943
rect 14599 14940 14611 14943
rect 15580 14940 15608 14971
rect 16390 14968 16396 14980
rect 16448 14968 16454 15020
rect 18322 15008 18328 15020
rect 16592 14980 18328 15008
rect 14599 14912 15608 14940
rect 14599 14909 14611 14912
rect 14553 14903 14611 14909
rect 15930 14900 15936 14952
rect 15988 14940 15994 14952
rect 16592 14940 16620 14980
rect 18322 14968 18328 14980
rect 18380 15008 18386 15020
rect 18785 15011 18843 15017
rect 18785 15008 18797 15011
rect 18380 14980 18797 15008
rect 18380 14968 18386 14980
rect 18785 14977 18797 14980
rect 18831 14977 18843 15011
rect 18785 14971 18843 14977
rect 19981 15011 20039 15017
rect 19981 14977 19993 15011
rect 20027 15008 20039 15011
rect 20070 15008 20076 15020
rect 20027 14980 20076 15008
rect 20027 14977 20039 14980
rect 19981 14971 20039 14977
rect 20070 14968 20076 14980
rect 20128 14968 20134 15020
rect 20530 14968 20536 15020
rect 20588 15008 20594 15020
rect 20916 15017 20944 15048
rect 22738 15036 22744 15048
rect 22796 15036 22802 15088
rect 23661 15079 23719 15085
rect 23661 15045 23673 15079
rect 23707 15076 23719 15079
rect 24394 15076 24400 15088
rect 23707 15048 24400 15076
rect 23707 15045 23719 15048
rect 23661 15039 23719 15045
rect 24394 15036 24400 15048
rect 24452 15036 24458 15088
rect 24762 15076 24768 15088
rect 24723 15048 24768 15076
rect 24762 15036 24768 15048
rect 24820 15036 24826 15088
rect 30926 15076 30932 15088
rect 30300 15048 30932 15076
rect 20717 15011 20775 15017
rect 20717 15008 20729 15011
rect 20588 14980 20729 15008
rect 20588 14968 20594 14980
rect 20717 14977 20729 14980
rect 20763 14977 20775 15011
rect 20717 14971 20775 14977
rect 20901 15011 20959 15017
rect 20901 14977 20913 15011
rect 20947 14977 20959 15011
rect 20901 14971 20959 14977
rect 26878 14968 26884 15020
rect 26936 15008 26942 15020
rect 30300 15017 30328 15048
rect 30926 15036 30932 15048
rect 30984 15036 30990 15088
rect 30101 15011 30159 15017
rect 30101 15008 30113 15011
rect 26936 14980 30113 15008
rect 26936 14968 26942 14980
rect 30101 14977 30113 14980
rect 30147 14977 30159 15011
rect 30101 14971 30159 14977
rect 30285 15011 30343 15017
rect 30285 14977 30297 15011
rect 30331 14977 30343 15011
rect 30285 14971 30343 14977
rect 30745 15011 30803 15017
rect 30745 14977 30757 15011
rect 30791 14977 30803 15011
rect 30745 14971 30803 14977
rect 15988 14912 16620 14940
rect 16669 14943 16727 14949
rect 15988 14900 15994 14912
rect 16669 14909 16681 14943
rect 16715 14909 16727 14943
rect 19705 14943 19763 14949
rect 19705 14940 19717 14943
rect 16669 14903 16727 14909
rect 19076 14912 19717 14940
rect 14090 14832 14096 14884
rect 14148 14872 14154 14884
rect 16684 14872 16712 14903
rect 14148 14844 16712 14872
rect 14148 14832 14154 14844
rect 16684 14804 16712 14844
rect 18414 14832 18420 14884
rect 18472 14872 18478 14884
rect 19076 14881 19104 14912
rect 19705 14909 19717 14912
rect 19751 14909 19763 14943
rect 20625 14943 20683 14949
rect 20625 14940 20637 14943
rect 19705 14903 19763 14909
rect 20088 14912 20637 14940
rect 19061 14875 19119 14881
rect 19061 14872 19073 14875
rect 18472 14844 19073 14872
rect 18472 14832 18478 14844
rect 19061 14841 19073 14844
rect 19107 14841 19119 14875
rect 19061 14835 19119 14841
rect 19245 14875 19303 14881
rect 19245 14841 19257 14875
rect 19291 14872 19303 14875
rect 20088 14872 20116 14912
rect 20625 14909 20637 14912
rect 20671 14940 20683 14943
rect 22373 14943 22431 14949
rect 22373 14940 22385 14943
rect 20671 14912 22385 14940
rect 20671 14909 20683 14912
rect 20625 14903 20683 14909
rect 22373 14909 22385 14912
rect 22419 14909 22431 14943
rect 30116 14940 30144 14971
rect 30760 14940 30788 14971
rect 34698 14968 34704 15020
rect 34756 15008 34762 15020
rect 35345 15011 35403 15017
rect 35345 15008 35357 15011
rect 34756 14980 35357 15008
rect 34756 14968 34762 14980
rect 35345 14977 35357 14980
rect 35391 14977 35403 15011
rect 35526 15008 35532 15020
rect 35487 14980 35532 15008
rect 35345 14971 35403 14977
rect 35526 14968 35532 14980
rect 35584 14968 35590 15020
rect 41322 14940 41328 14952
rect 30116 14912 30788 14940
rect 41283 14912 41328 14940
rect 22373 14903 22431 14909
rect 41322 14900 41328 14912
rect 41380 14900 41386 14952
rect 41414 14900 41420 14952
rect 41472 14940 41478 14952
rect 41693 14943 41751 14949
rect 41693 14940 41705 14943
rect 41472 14912 41705 14940
rect 41472 14900 41478 14912
rect 41693 14909 41705 14912
rect 41739 14909 41751 14943
rect 41693 14903 41751 14909
rect 41877 14943 41935 14949
rect 41877 14909 41889 14943
rect 41923 14940 41935 14943
rect 41966 14940 41972 14952
rect 41923 14912 41972 14940
rect 41923 14909 41935 14912
rect 41877 14903 41935 14909
rect 41966 14900 41972 14912
rect 42024 14900 42030 14952
rect 19291 14844 20116 14872
rect 20165 14875 20223 14881
rect 19291 14841 19303 14844
rect 19245 14835 19303 14841
rect 20165 14841 20177 14875
rect 20211 14872 20223 14875
rect 22278 14872 22284 14884
rect 20211 14844 22284 14872
rect 20211 14841 20223 14844
rect 20165 14835 20223 14841
rect 22278 14832 22284 14844
rect 22336 14832 22342 14884
rect 22925 14875 22983 14881
rect 22925 14841 22937 14875
rect 22971 14872 22983 14875
rect 38470 14872 38476 14884
rect 22971 14844 38476 14872
rect 22971 14841 22983 14844
rect 22925 14835 22983 14841
rect 38470 14832 38476 14844
rect 38528 14832 38534 14884
rect 17954 14804 17960 14816
rect 16684 14776 17960 14804
rect 17954 14764 17960 14776
rect 18012 14764 18018 14816
rect 19610 14764 19616 14816
rect 19668 14804 19674 14816
rect 19797 14807 19855 14813
rect 19797 14804 19809 14807
rect 19668 14776 19809 14804
rect 19668 14764 19674 14776
rect 19797 14773 19809 14776
rect 19843 14773 19855 14807
rect 19797 14767 19855 14773
rect 21085 14807 21143 14813
rect 21085 14773 21097 14807
rect 21131 14804 21143 14807
rect 22370 14804 22376 14816
rect 21131 14776 22376 14804
rect 21131 14773 21143 14776
rect 21085 14767 21143 14773
rect 22370 14764 22376 14776
rect 22428 14764 22434 14816
rect 22646 14764 22652 14816
rect 22704 14804 22710 14816
rect 22741 14807 22799 14813
rect 22741 14804 22753 14807
rect 22704 14776 22753 14804
rect 22704 14764 22710 14776
rect 22741 14773 22753 14776
rect 22787 14773 22799 14807
rect 22741 14767 22799 14773
rect 23474 14764 23480 14816
rect 23532 14804 23538 14816
rect 23569 14807 23627 14813
rect 23569 14804 23581 14807
rect 23532 14776 23581 14804
rect 23532 14764 23538 14776
rect 23569 14773 23581 14776
rect 23615 14773 23627 14807
rect 23569 14767 23627 14773
rect 24670 14764 24676 14816
rect 24728 14804 24734 14816
rect 24949 14807 25007 14813
rect 24949 14804 24961 14807
rect 24728 14776 24961 14804
rect 24728 14764 24734 14776
rect 24949 14773 24961 14776
rect 24995 14773 25007 14807
rect 24949 14767 25007 14773
rect 25133 14807 25191 14813
rect 25133 14773 25145 14807
rect 25179 14804 25191 14807
rect 25222 14804 25228 14816
rect 25179 14776 25228 14804
rect 25179 14773 25191 14776
rect 25133 14767 25191 14773
rect 25222 14764 25228 14776
rect 25280 14764 25286 14816
rect 30190 14804 30196 14816
rect 30151 14776 30196 14804
rect 30190 14764 30196 14776
rect 30248 14764 30254 14816
rect 31113 14807 31171 14813
rect 31113 14773 31125 14807
rect 31159 14804 31171 14807
rect 31662 14804 31668 14816
rect 31159 14776 31668 14804
rect 31159 14773 31171 14776
rect 31113 14767 31171 14773
rect 31662 14764 31668 14776
rect 31720 14764 31726 14816
rect 35713 14807 35771 14813
rect 35713 14773 35725 14807
rect 35759 14804 35771 14807
rect 35802 14804 35808 14816
rect 35759 14776 35808 14804
rect 35759 14773 35771 14776
rect 35713 14767 35771 14773
rect 35802 14764 35808 14776
rect 35860 14764 35866 14816
rect 1104 14714 42872 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 42872 14714
rect 1104 14640 42872 14662
rect 2222 14600 2228 14612
rect 2183 14572 2228 14600
rect 2222 14560 2228 14572
rect 2280 14560 2286 14612
rect 13357 14603 13415 14609
rect 13357 14569 13369 14603
rect 13403 14600 13415 14603
rect 13814 14600 13820 14612
rect 13403 14572 13820 14600
rect 13403 14569 13415 14572
rect 13357 14563 13415 14569
rect 13814 14560 13820 14572
rect 13872 14560 13878 14612
rect 15194 14560 15200 14612
rect 15252 14600 15258 14612
rect 19610 14600 19616 14612
rect 15252 14572 15884 14600
rect 19571 14572 19616 14600
rect 15252 14560 15258 14572
rect 15562 14532 15568 14544
rect 12360 14504 14587 14532
rect 2317 14399 2375 14405
rect 2317 14365 2329 14399
rect 2363 14396 2375 14399
rect 2958 14396 2964 14408
rect 2363 14368 2964 14396
rect 2363 14365 2375 14368
rect 2317 14359 2375 14365
rect 2958 14356 2964 14368
rect 3016 14396 3022 14408
rect 11606 14396 11612 14408
rect 3016 14368 11612 14396
rect 3016 14356 3022 14368
rect 11606 14356 11612 14368
rect 11664 14356 11670 14408
rect 12360 14405 12388 14504
rect 13538 14464 13544 14476
rect 13280 14436 13544 14464
rect 13280 14405 13308 14436
rect 13538 14424 13544 14436
rect 13596 14424 13602 14476
rect 12345 14399 12403 14405
rect 12345 14365 12357 14399
rect 12391 14365 12403 14399
rect 12345 14359 12403 14365
rect 13265 14399 13323 14405
rect 13265 14365 13277 14399
rect 13311 14365 13323 14399
rect 13446 14396 13452 14408
rect 13407 14368 13452 14396
rect 13265 14359 13323 14365
rect 13446 14356 13452 14368
rect 13504 14356 13510 14408
rect 11790 14220 11796 14272
rect 11848 14260 11854 14272
rect 12161 14263 12219 14269
rect 12161 14260 12173 14263
rect 11848 14232 12173 14260
rect 11848 14220 11854 14232
rect 12161 14229 12173 14232
rect 12207 14229 12219 14263
rect 14366 14260 14372 14272
rect 14327 14232 14372 14260
rect 12161 14223 12219 14229
rect 14366 14220 14372 14232
rect 14424 14220 14430 14272
rect 14559 14260 14587 14504
rect 14752 14504 15568 14532
rect 14752 14405 14780 14504
rect 15562 14492 15568 14504
rect 15620 14492 15626 14544
rect 15654 14492 15660 14544
rect 15712 14492 15718 14544
rect 15856 14532 15884 14572
rect 19610 14560 19616 14572
rect 19668 14560 19674 14612
rect 20717 14603 20775 14609
rect 20717 14569 20729 14603
rect 20763 14600 20775 14603
rect 20990 14600 20996 14612
rect 20763 14572 20996 14600
rect 20763 14569 20775 14572
rect 20717 14563 20775 14569
rect 20990 14560 20996 14572
rect 21048 14560 21054 14612
rect 21729 14603 21787 14609
rect 21729 14569 21741 14603
rect 21775 14600 21787 14603
rect 22186 14600 22192 14612
rect 21775 14572 22192 14600
rect 21775 14569 21787 14572
rect 21729 14563 21787 14569
rect 22186 14560 22192 14572
rect 22244 14560 22250 14612
rect 22738 14560 22744 14612
rect 22796 14600 22802 14612
rect 24857 14603 24915 14609
rect 24857 14600 24869 14603
rect 22796 14572 24869 14600
rect 22796 14560 22802 14572
rect 24857 14569 24869 14572
rect 24903 14569 24915 14603
rect 24857 14563 24915 14569
rect 34514 14560 34520 14612
rect 34572 14600 34578 14612
rect 35526 14600 35532 14612
rect 34572 14572 35532 14600
rect 34572 14560 34578 14572
rect 35526 14560 35532 14572
rect 35584 14560 35590 14612
rect 35805 14603 35863 14609
rect 35805 14569 35817 14603
rect 35851 14600 35863 14603
rect 35894 14600 35900 14612
rect 35851 14572 35900 14600
rect 35851 14569 35863 14572
rect 35805 14563 35863 14569
rect 35894 14560 35900 14572
rect 35952 14600 35958 14612
rect 36262 14600 36268 14612
rect 35952 14572 36268 14600
rect 35952 14560 35958 14572
rect 36262 14560 36268 14572
rect 36320 14560 36326 14612
rect 41414 14600 41420 14612
rect 41375 14572 41420 14600
rect 41414 14560 41420 14572
rect 41472 14560 41478 14612
rect 41966 14600 41972 14612
rect 41927 14572 41972 14600
rect 41966 14560 41972 14572
rect 42024 14560 42030 14612
rect 23566 14532 23572 14544
rect 15856 14504 17908 14532
rect 23527 14504 23572 14532
rect 15473 14467 15531 14473
rect 15473 14464 15485 14467
rect 14844 14436 15485 14464
rect 14844 14405 14872 14436
rect 15473 14433 15485 14436
rect 15519 14433 15531 14467
rect 15672 14464 15700 14492
rect 15856 14473 15884 14504
rect 15749 14467 15807 14473
rect 15749 14464 15761 14467
rect 15672 14436 15761 14464
rect 15473 14427 15531 14433
rect 15749 14433 15761 14436
rect 15795 14433 15807 14467
rect 15749 14427 15807 14433
rect 15841 14467 15899 14473
rect 15841 14433 15853 14467
rect 15887 14433 15899 14467
rect 15841 14427 15899 14433
rect 17402 14424 17408 14476
rect 17460 14464 17466 14476
rect 17880 14473 17908 14504
rect 23566 14492 23572 14504
rect 23624 14492 23630 14544
rect 31846 14492 31852 14544
rect 31904 14532 31910 14544
rect 31904 14504 41368 14532
rect 31904 14492 31910 14504
rect 17589 14467 17647 14473
rect 17589 14464 17601 14467
rect 17460 14436 17601 14464
rect 17460 14424 17466 14436
rect 17589 14433 17601 14436
rect 17635 14433 17647 14467
rect 17589 14427 17647 14433
rect 17865 14467 17923 14473
rect 17865 14433 17877 14467
rect 17911 14464 17923 14467
rect 18046 14464 18052 14476
rect 17911 14436 18052 14464
rect 17911 14433 17923 14436
rect 17865 14427 17923 14433
rect 18046 14424 18052 14436
rect 18104 14464 18110 14476
rect 19245 14467 19303 14473
rect 19245 14464 19257 14467
rect 18104 14436 19257 14464
rect 18104 14424 18110 14436
rect 19245 14433 19257 14436
rect 19291 14433 19303 14467
rect 19245 14427 19303 14433
rect 20162 14424 20168 14476
rect 20220 14464 20226 14476
rect 20349 14467 20407 14473
rect 20349 14464 20361 14467
rect 20220 14436 20361 14464
rect 20220 14424 20226 14436
rect 20349 14433 20361 14436
rect 20395 14433 20407 14467
rect 20349 14427 20407 14433
rect 34532 14436 36768 14464
rect 14645 14399 14703 14405
rect 14645 14365 14657 14399
rect 14691 14365 14703 14399
rect 14645 14359 14703 14365
rect 14737 14399 14795 14405
rect 14737 14365 14749 14399
rect 14783 14365 14795 14399
rect 14737 14359 14795 14365
rect 14829 14399 14887 14405
rect 14829 14365 14841 14399
rect 14875 14365 14887 14399
rect 15010 14396 15016 14408
rect 14971 14368 15016 14396
rect 14829 14359 14887 14365
rect 14660 14328 14688 14359
rect 15010 14356 15016 14368
rect 15068 14356 15074 14408
rect 15102 14356 15108 14408
rect 15160 14396 15166 14408
rect 15657 14399 15715 14405
rect 15657 14396 15669 14399
rect 15160 14368 15669 14396
rect 15160 14356 15166 14368
rect 15657 14365 15669 14368
rect 15703 14365 15715 14399
rect 15930 14396 15936 14408
rect 15891 14368 15936 14396
rect 15657 14359 15715 14365
rect 15930 14356 15936 14368
rect 15988 14356 15994 14408
rect 19426 14396 19432 14408
rect 19387 14368 19432 14396
rect 19426 14356 19432 14368
rect 19484 14356 19490 14408
rect 20254 14396 20260 14408
rect 20215 14368 20260 14396
rect 20254 14356 20260 14368
rect 20312 14356 20318 14408
rect 20438 14356 20444 14408
rect 20496 14396 20502 14408
rect 20533 14399 20591 14405
rect 20533 14396 20545 14399
rect 20496 14368 20545 14396
rect 20496 14356 20502 14368
rect 20533 14365 20545 14368
rect 20579 14365 20591 14399
rect 20533 14359 20591 14365
rect 21361 14399 21419 14405
rect 21361 14365 21373 14399
rect 21407 14365 21419 14399
rect 23385 14399 23443 14405
rect 23385 14396 23397 14399
rect 21361 14359 21419 14365
rect 22066 14368 23397 14396
rect 16390 14328 16396 14340
rect 14660 14300 16396 14328
rect 16390 14288 16396 14300
rect 16448 14288 16454 14340
rect 21376 14328 21404 14359
rect 21726 14328 21732 14340
rect 20456 14300 21404 14328
rect 21687 14300 21732 14328
rect 20456 14272 20484 14300
rect 21726 14288 21732 14300
rect 21784 14288 21790 14340
rect 16666 14260 16672 14272
rect 14559 14232 16672 14260
rect 16666 14220 16672 14232
rect 16724 14220 16730 14272
rect 20438 14220 20444 14272
rect 20496 14220 20502 14272
rect 21913 14263 21971 14269
rect 21913 14229 21925 14263
rect 21959 14260 21971 14263
rect 22066 14260 22094 14368
rect 23385 14365 23397 14368
rect 23431 14365 23443 14399
rect 26234 14396 26240 14408
rect 26195 14368 26240 14396
rect 23385 14359 23443 14365
rect 26234 14356 26240 14368
rect 26292 14396 26298 14408
rect 26694 14396 26700 14408
rect 26292 14368 26700 14396
rect 26292 14356 26298 14368
rect 26694 14356 26700 14368
rect 26752 14356 26758 14408
rect 26964 14399 27022 14405
rect 26964 14365 26976 14399
rect 27010 14365 27022 14399
rect 26964 14359 27022 14365
rect 29549 14399 29607 14405
rect 29549 14365 29561 14399
rect 29595 14396 29607 14399
rect 29816 14399 29874 14405
rect 29595 14368 29684 14396
rect 29595 14365 29607 14368
rect 29549 14359 29607 14365
rect 25992 14331 26050 14337
rect 25992 14297 26004 14331
rect 26038 14328 26050 14331
rect 26142 14328 26148 14340
rect 26038 14300 26148 14328
rect 26038 14297 26050 14300
rect 25992 14291 26050 14297
rect 26142 14288 26148 14300
rect 26200 14288 26206 14340
rect 26878 14288 26884 14340
rect 26936 14328 26942 14340
rect 26988 14328 27016 14359
rect 26936 14300 27016 14328
rect 26936 14288 26942 14300
rect 21959 14232 22094 14260
rect 28077 14263 28135 14269
rect 21959 14229 21971 14232
rect 21913 14223 21971 14229
rect 28077 14229 28089 14263
rect 28123 14260 28135 14263
rect 28994 14260 29000 14272
rect 28123 14232 29000 14260
rect 28123 14229 28135 14232
rect 28077 14223 28135 14229
rect 28994 14220 29000 14232
rect 29052 14220 29058 14272
rect 29656 14260 29684 14368
rect 29816 14365 29828 14399
rect 29862 14365 29874 14399
rect 29816 14359 29874 14365
rect 29730 14288 29736 14340
rect 29788 14328 29794 14340
rect 29840 14328 29868 14359
rect 31754 14356 31760 14408
rect 31812 14396 31818 14408
rect 32030 14396 32036 14408
rect 31812 14368 32036 14396
rect 31812 14356 31818 14368
rect 32030 14356 32036 14368
rect 32088 14356 32094 14408
rect 32214 14356 32220 14408
rect 32272 14356 32278 14408
rect 33594 14396 33600 14408
rect 33555 14368 33600 14396
rect 33594 14356 33600 14368
rect 33652 14356 33658 14408
rect 33778 14396 33784 14408
rect 33739 14368 33784 14396
rect 33778 14356 33784 14368
rect 33836 14356 33842 14408
rect 34532 14340 34560 14436
rect 34606 14356 34612 14408
rect 34664 14396 34670 14408
rect 34885 14399 34943 14405
rect 34885 14396 34897 14399
rect 34664 14368 34897 14396
rect 34664 14356 34670 14368
rect 34885 14365 34897 14368
rect 34931 14396 34943 14399
rect 35710 14396 35716 14408
rect 34931 14368 35716 14396
rect 34931 14365 34943 14368
rect 34885 14359 34943 14365
rect 35710 14356 35716 14368
rect 35768 14356 35774 14408
rect 36078 14396 36084 14408
rect 36039 14368 36084 14396
rect 36078 14356 36084 14368
rect 36136 14356 36142 14408
rect 36740 14405 36768 14436
rect 36541 14399 36599 14405
rect 36541 14365 36553 14399
rect 36587 14365 36599 14399
rect 36541 14359 36599 14365
rect 36725 14399 36783 14405
rect 36725 14365 36737 14399
rect 36771 14396 36783 14399
rect 37182 14396 37188 14408
rect 36771 14368 37188 14396
rect 36771 14365 36783 14368
rect 36725 14359 36783 14365
rect 30374 14328 30380 14340
rect 29788 14300 29868 14328
rect 29932 14300 30380 14328
rect 29788 14288 29794 14300
rect 29932 14260 29960 14300
rect 30374 14288 30380 14300
rect 30432 14288 30438 14340
rect 33045 14331 33103 14337
rect 33045 14297 33057 14331
rect 33091 14328 33103 14331
rect 34514 14328 34520 14340
rect 33091 14300 34520 14328
rect 33091 14297 33103 14300
rect 33045 14291 33103 14297
rect 34514 14288 34520 14300
rect 34572 14288 34578 14340
rect 35069 14331 35127 14337
rect 35069 14297 35081 14331
rect 35115 14328 35127 14331
rect 35342 14328 35348 14340
rect 35115 14300 35348 14328
rect 35115 14297 35127 14300
rect 35069 14291 35127 14297
rect 35342 14288 35348 14300
rect 35400 14288 35406 14340
rect 35526 14288 35532 14340
rect 35584 14328 35590 14340
rect 36556 14328 36584 14359
rect 37182 14356 37188 14368
rect 37240 14356 37246 14408
rect 41230 14356 41236 14408
rect 41288 14396 41294 14408
rect 41340 14405 41368 14504
rect 41325 14399 41383 14405
rect 41325 14396 41337 14399
rect 41288 14368 41337 14396
rect 41288 14356 41294 14368
rect 41325 14365 41337 14368
rect 41371 14365 41383 14399
rect 41325 14359 41383 14365
rect 35584 14300 36584 14328
rect 35584 14288 35590 14300
rect 29656 14232 29960 14260
rect 30282 14220 30288 14272
rect 30340 14260 30346 14272
rect 30929 14263 30987 14269
rect 30929 14260 30941 14263
rect 30340 14232 30941 14260
rect 30340 14220 30346 14232
rect 30929 14229 30941 14232
rect 30975 14229 30987 14263
rect 30929 14223 30987 14229
rect 33410 14220 33416 14272
rect 33468 14260 33474 14272
rect 33689 14263 33747 14269
rect 33689 14260 33701 14263
rect 33468 14232 33701 14260
rect 33468 14220 33474 14232
rect 33689 14229 33701 14232
rect 33735 14229 33747 14263
rect 34698 14260 34704 14272
rect 34611 14232 34704 14260
rect 33689 14223 33747 14229
rect 34698 14220 34704 14232
rect 34756 14260 34762 14272
rect 34974 14260 34980 14272
rect 34756 14232 34980 14260
rect 34756 14220 34762 14232
rect 34974 14220 34980 14232
rect 35032 14220 35038 14272
rect 36630 14260 36636 14272
rect 36591 14232 36636 14260
rect 36630 14220 36636 14232
rect 36688 14220 36694 14272
rect 1104 14170 42872 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 42872 14170
rect 1104 14096 42872 14118
rect 15473 14059 15531 14065
rect 15473 14025 15485 14059
rect 15519 14056 15531 14059
rect 15930 14056 15936 14068
rect 15519 14028 15936 14056
rect 15519 14025 15531 14028
rect 15473 14019 15531 14025
rect 15930 14016 15936 14028
rect 15988 14016 15994 14068
rect 16669 14059 16727 14065
rect 16669 14056 16681 14059
rect 16040 14028 16681 14056
rect 14366 13997 14372 14000
rect 14360 13988 14372 13997
rect 14327 13960 14372 13988
rect 14360 13951 14372 13960
rect 14366 13948 14372 13951
rect 14424 13948 14430 14000
rect 15654 13948 15660 14000
rect 15712 13988 15718 14000
rect 16040 13988 16068 14028
rect 16669 14025 16681 14028
rect 16715 14025 16727 14059
rect 16669 14019 16727 14025
rect 19889 14059 19947 14065
rect 19889 14025 19901 14059
rect 19935 14056 19947 14059
rect 20254 14056 20260 14068
rect 19935 14028 20260 14056
rect 19935 14025 19947 14028
rect 19889 14019 19947 14025
rect 20254 14016 20260 14028
rect 20312 14016 20318 14068
rect 24394 14016 24400 14068
rect 24452 14056 24458 14068
rect 24581 14059 24639 14065
rect 24581 14056 24593 14059
rect 24452 14028 24593 14056
rect 24452 14016 24458 14028
rect 24581 14025 24593 14028
rect 24627 14025 24639 14059
rect 26142 14056 26148 14068
rect 26103 14028 26148 14056
rect 24581 14019 24639 14025
rect 26142 14016 26148 14028
rect 26200 14016 26206 14068
rect 31846 14056 31852 14068
rect 26252 14028 31852 14056
rect 15712 13960 16068 13988
rect 15712 13948 15718 13960
rect 16574 13948 16580 14000
rect 16632 13988 16638 14000
rect 16821 13991 16879 13997
rect 16821 13988 16833 13991
rect 16632 13960 16833 13988
rect 16632 13948 16638 13960
rect 16821 13957 16833 13960
rect 16867 13957 16879 13991
rect 16821 13951 16879 13957
rect 17037 13991 17095 13997
rect 17037 13957 17049 13991
rect 17083 13957 17095 13991
rect 20162 13988 20168 14000
rect 17037 13951 17095 13957
rect 18064 13960 20168 13988
rect 11790 13920 11796 13932
rect 11751 13892 11796 13920
rect 11790 13880 11796 13892
rect 11848 13880 11854 13932
rect 14090 13920 14096 13932
rect 14051 13892 14096 13920
rect 14090 13880 14096 13892
rect 14148 13880 14154 13932
rect 1946 13852 1952 13864
rect 1907 13824 1952 13852
rect 1946 13812 1952 13824
rect 2004 13812 2010 13864
rect 2133 13855 2191 13861
rect 2133 13821 2145 13855
rect 2179 13852 2191 13855
rect 2774 13852 2780 13864
rect 2179 13824 2780 13852
rect 2179 13821 2191 13824
rect 2133 13815 2191 13821
rect 2774 13812 2780 13824
rect 2832 13812 2838 13864
rect 2866 13812 2872 13864
rect 2924 13852 2930 13864
rect 11974 13852 11980 13864
rect 2924 13824 2969 13852
rect 11935 13824 11980 13852
rect 2924 13812 2930 13824
rect 11974 13812 11980 13824
rect 12032 13812 12038 13864
rect 13630 13852 13636 13864
rect 13591 13824 13636 13852
rect 13630 13812 13636 13824
rect 13688 13812 13694 13864
rect 16942 13812 16948 13864
rect 17000 13852 17006 13864
rect 17052 13852 17080 13951
rect 18064 13929 18092 13960
rect 20162 13948 20168 13960
rect 20220 13948 20226 14000
rect 20714 13948 20720 14000
rect 20772 13988 20778 14000
rect 21913 13991 21971 13997
rect 21913 13988 21925 13991
rect 20772 13960 21925 13988
rect 20772 13948 20778 13960
rect 21913 13957 21925 13960
rect 21959 13957 21971 13991
rect 21913 13951 21971 13957
rect 22094 13948 22100 14000
rect 22152 13988 22158 14000
rect 22152 13960 22197 13988
rect 22152 13948 22158 13960
rect 22278 13948 22284 14000
rect 22336 13988 22342 14000
rect 22802 13991 22860 13997
rect 22802 13988 22814 13991
rect 22336 13960 22814 13988
rect 22336 13948 22342 13960
rect 22802 13957 22814 13960
rect 22848 13957 22860 13991
rect 22802 13951 22860 13957
rect 23106 13948 23112 14000
rect 23164 13988 23170 14000
rect 26252 13988 26280 14028
rect 31846 14016 31852 14028
rect 31904 14016 31910 14068
rect 32214 14056 32220 14068
rect 32175 14028 32220 14056
rect 32214 14016 32220 14028
rect 32272 14016 32278 14068
rect 33321 14059 33379 14065
rect 33321 14025 33333 14059
rect 33367 14056 33379 14059
rect 35986 14056 35992 14068
rect 33367 14028 35992 14056
rect 33367 14025 33379 14028
rect 33321 14019 33379 14025
rect 35986 14016 35992 14028
rect 36044 14016 36050 14068
rect 23164 13960 26280 13988
rect 27709 13991 27767 13997
rect 23164 13948 23170 13960
rect 27709 13957 27721 13991
rect 27755 13988 27767 13991
rect 30006 13988 30012 14000
rect 27755 13960 30012 13988
rect 27755 13957 27767 13960
rect 27709 13951 27767 13957
rect 30006 13948 30012 13960
rect 30064 13948 30070 14000
rect 31573 13991 31631 13997
rect 31573 13957 31585 13991
rect 31619 13988 31631 13991
rect 31619 13960 31708 13988
rect 31619 13957 31631 13960
rect 31573 13951 31631 13957
rect 18049 13923 18107 13929
rect 18049 13889 18061 13923
rect 18095 13889 18107 13923
rect 19797 13923 19855 13929
rect 19797 13920 19809 13923
rect 18049 13883 18107 13889
rect 18156 13892 19809 13920
rect 18156 13852 18184 13892
rect 19797 13889 19809 13892
rect 19843 13889 19855 13923
rect 19797 13883 19855 13889
rect 17000 13824 18184 13852
rect 18233 13855 18291 13861
rect 17000 13812 17006 13824
rect 18233 13821 18245 13855
rect 18279 13852 18291 13855
rect 18322 13852 18328 13864
rect 18279 13824 18328 13852
rect 18279 13821 18291 13824
rect 18233 13815 18291 13821
rect 18322 13812 18328 13824
rect 18380 13812 18386 13864
rect 19812 13784 19840 13883
rect 19978 13880 19984 13932
rect 20036 13920 20042 13932
rect 20036 13892 20081 13920
rect 20036 13880 20042 13892
rect 20346 13880 20352 13932
rect 20404 13920 20410 13932
rect 20441 13923 20499 13929
rect 20441 13920 20453 13923
rect 20404 13892 20453 13920
rect 20404 13880 20410 13892
rect 20441 13889 20453 13892
rect 20487 13889 20499 13923
rect 21358 13920 21364 13932
rect 20441 13883 20499 13889
rect 20640 13892 21364 13920
rect 20346 13784 20352 13796
rect 19812 13756 20352 13784
rect 20346 13744 20352 13756
rect 20404 13744 20410 13796
rect 20640 13793 20668 13892
rect 21358 13880 21364 13892
rect 21416 13880 21422 13932
rect 22112 13920 22140 13948
rect 31680 13932 31708 13960
rect 33594 13948 33600 14000
rect 33652 13988 33658 14000
rect 34701 13991 34759 13997
rect 34701 13988 34713 13991
rect 33652 13960 34713 13988
rect 33652 13948 33658 13960
rect 34701 13957 34713 13960
rect 34747 13957 34759 13991
rect 34701 13951 34759 13957
rect 22462 13920 22468 13932
rect 22112 13892 22468 13920
rect 22462 13880 22468 13892
rect 22520 13920 22526 13932
rect 22557 13923 22615 13929
rect 22557 13920 22569 13923
rect 22520 13892 22569 13920
rect 22520 13880 22526 13892
rect 22557 13889 22569 13892
rect 22603 13889 22615 13923
rect 22557 13883 22615 13889
rect 24578 13880 24584 13932
rect 24636 13920 24642 13932
rect 24765 13923 24823 13929
rect 24765 13920 24777 13923
rect 24636 13892 24777 13920
rect 24636 13880 24642 13892
rect 24765 13889 24777 13892
rect 24811 13889 24823 13923
rect 25222 13920 25228 13932
rect 25183 13892 25228 13920
rect 24765 13883 24823 13889
rect 25222 13880 25228 13892
rect 25280 13880 25286 13932
rect 25409 13923 25467 13929
rect 25409 13889 25421 13923
rect 25455 13889 25467 13923
rect 25409 13883 25467 13889
rect 26329 13923 26387 13929
rect 26329 13889 26341 13923
rect 26375 13920 26387 13923
rect 28166 13920 28172 13932
rect 26375 13892 28172 13920
rect 26375 13889 26387 13892
rect 26329 13883 26387 13889
rect 20714 13812 20720 13864
rect 20772 13852 20778 13864
rect 24670 13852 24676 13864
rect 20772 13824 20817 13852
rect 23952 13824 24676 13852
rect 20772 13812 20778 13824
rect 23952 13793 23980 13824
rect 24670 13812 24676 13824
rect 24728 13852 24734 13864
rect 25424 13852 25452 13883
rect 28166 13880 28172 13892
rect 28224 13880 28230 13932
rect 30098 13920 30104 13932
rect 30059 13892 30104 13920
rect 30098 13880 30104 13892
rect 30156 13880 30162 13932
rect 30282 13920 30288 13932
rect 30243 13892 30288 13920
rect 30282 13880 30288 13892
rect 30340 13880 30346 13932
rect 31113 13923 31171 13929
rect 31113 13889 31125 13923
rect 31159 13920 31171 13923
rect 31159 13892 31616 13920
rect 31159 13889 31171 13892
rect 31113 13883 31171 13889
rect 24728 13824 25452 13852
rect 24728 13812 24734 13824
rect 30190 13812 30196 13864
rect 30248 13852 30254 13864
rect 31205 13855 31263 13861
rect 31205 13852 31217 13855
rect 30248 13824 31217 13852
rect 30248 13812 30254 13824
rect 31205 13821 31217 13824
rect 31251 13852 31263 13855
rect 31588 13852 31616 13892
rect 31662 13880 31668 13932
rect 31720 13920 31726 13932
rect 32125 13923 32183 13929
rect 32125 13920 32137 13923
rect 31720 13892 32137 13920
rect 31720 13880 31726 13892
rect 32125 13889 32137 13892
rect 32171 13889 32183 13923
rect 32125 13883 32183 13889
rect 32309 13923 32367 13929
rect 32309 13889 32321 13923
rect 32355 13889 32367 13923
rect 33226 13920 33232 13932
rect 33187 13892 33232 13920
rect 32309 13883 32367 13889
rect 31754 13852 31760 13864
rect 31251 13824 31524 13852
rect 31588 13824 31760 13852
rect 31251 13821 31263 13824
rect 31205 13815 31263 13821
rect 20625 13787 20683 13793
rect 20625 13753 20637 13787
rect 20671 13753 20683 13787
rect 20625 13747 20683 13753
rect 23937 13787 23995 13793
rect 23937 13753 23949 13787
rect 23983 13753 23995 13787
rect 27522 13784 27528 13796
rect 27483 13756 27528 13784
rect 23937 13747 23995 13753
rect 27522 13744 27528 13756
rect 27580 13744 27586 13796
rect 31496 13784 31524 13824
rect 31754 13812 31760 13824
rect 31812 13812 31818 13864
rect 32324 13852 32352 13883
rect 33226 13880 33232 13892
rect 33284 13880 33290 13932
rect 34422 13880 34428 13932
rect 34480 13920 34486 13932
rect 34517 13923 34575 13929
rect 34517 13920 34529 13923
rect 34480 13892 34529 13920
rect 34480 13880 34486 13892
rect 34517 13889 34529 13892
rect 34563 13889 34575 13923
rect 34517 13883 34575 13889
rect 34609 13923 34667 13929
rect 34609 13889 34621 13923
rect 34655 13889 34667 13923
rect 34609 13883 34667 13889
rect 31864 13824 32352 13852
rect 33413 13855 33471 13861
rect 31864 13784 31892 13824
rect 33413 13821 33425 13855
rect 33459 13821 33471 13855
rect 33413 13815 33471 13821
rect 31496 13756 31892 13784
rect 33042 13744 33048 13796
rect 33100 13784 33106 13796
rect 33428 13784 33456 13815
rect 34624 13796 34652 13883
rect 34790 13880 34796 13932
rect 34848 13929 34854 13932
rect 34848 13923 34877 13929
rect 34865 13889 34877 13923
rect 34848 13883 34877 13889
rect 35621 13923 35679 13929
rect 35621 13889 35633 13923
rect 35667 13920 35679 13923
rect 35710 13920 35716 13932
rect 35667 13892 35716 13920
rect 35667 13889 35679 13892
rect 35621 13883 35679 13889
rect 34848 13880 34854 13883
rect 35710 13880 35716 13892
rect 35768 13880 35774 13932
rect 35802 13880 35808 13932
rect 35860 13920 35866 13932
rect 37366 13920 37372 13932
rect 35860 13892 37372 13920
rect 35860 13880 35866 13892
rect 37366 13880 37372 13892
rect 37424 13880 37430 13932
rect 34974 13812 34980 13864
rect 35032 13852 35038 13864
rect 35897 13855 35955 13861
rect 35032 13824 35077 13852
rect 35032 13812 35038 13824
rect 35897 13821 35909 13855
rect 35943 13852 35955 13855
rect 36170 13852 36176 13864
rect 35943 13824 36176 13852
rect 35943 13821 35955 13824
rect 35897 13815 35955 13821
rect 36170 13812 36176 13824
rect 36228 13812 36234 13864
rect 34606 13784 34612 13796
rect 33100 13756 33456 13784
rect 34519 13756 34612 13784
rect 33100 13744 33106 13756
rect 34606 13744 34612 13756
rect 34664 13784 34670 13796
rect 36814 13784 36820 13796
rect 34664 13756 36820 13784
rect 34664 13744 34670 13756
rect 36814 13744 36820 13756
rect 36872 13744 36878 13796
rect 16850 13716 16856 13728
rect 16811 13688 16856 13716
rect 16850 13676 16856 13688
rect 16908 13676 16914 13728
rect 17862 13716 17868 13728
rect 17823 13688 17868 13716
rect 17862 13676 17868 13688
rect 17920 13676 17926 13728
rect 19978 13676 19984 13728
rect 20036 13716 20042 13728
rect 20438 13716 20444 13728
rect 20036 13688 20444 13716
rect 20036 13676 20042 13688
rect 20438 13676 20444 13688
rect 20496 13716 20502 13728
rect 20533 13719 20591 13725
rect 20533 13716 20545 13719
rect 20496 13688 20545 13716
rect 20496 13676 20502 13688
rect 20533 13685 20545 13688
rect 20579 13685 20591 13719
rect 25314 13716 25320 13728
rect 25275 13688 25320 13716
rect 20533 13679 20591 13685
rect 25314 13676 25320 13688
rect 25372 13676 25378 13728
rect 30101 13719 30159 13725
rect 30101 13685 30113 13719
rect 30147 13716 30159 13719
rect 30742 13716 30748 13728
rect 30147 13688 30748 13716
rect 30147 13685 30159 13688
rect 30101 13679 30159 13685
rect 30742 13676 30748 13688
rect 30800 13676 30806 13728
rect 30929 13719 30987 13725
rect 30929 13685 30941 13719
rect 30975 13716 30987 13719
rect 31018 13716 31024 13728
rect 30975 13688 31024 13716
rect 30975 13685 30987 13688
rect 30929 13679 30987 13685
rect 31018 13676 31024 13688
rect 31076 13676 31082 13728
rect 32858 13716 32864 13728
rect 32819 13688 32864 13716
rect 32858 13676 32864 13688
rect 32916 13676 32922 13728
rect 34330 13716 34336 13728
rect 34291 13688 34336 13716
rect 34330 13676 34336 13688
rect 34388 13676 34394 13728
rect 41782 13716 41788 13728
rect 41743 13688 41788 13716
rect 41782 13676 41788 13688
rect 41840 13676 41846 13728
rect 1104 13626 42872 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 42872 13626
rect 1104 13552 42872 13574
rect 1946 13472 1952 13524
rect 2004 13512 2010 13524
rect 2041 13515 2099 13521
rect 2041 13512 2053 13515
rect 2004 13484 2053 13512
rect 2004 13472 2010 13484
rect 2041 13481 2053 13484
rect 2087 13481 2099 13515
rect 2774 13512 2780 13524
rect 2735 13484 2780 13512
rect 2041 13475 2099 13481
rect 2774 13472 2780 13484
rect 2832 13472 2838 13524
rect 11974 13472 11980 13524
rect 12032 13512 12038 13524
rect 12069 13515 12127 13521
rect 12069 13512 12081 13515
rect 12032 13484 12081 13512
rect 12032 13472 12038 13484
rect 12069 13481 12081 13484
rect 12115 13481 12127 13515
rect 12069 13475 12127 13481
rect 21545 13515 21603 13521
rect 21545 13481 21557 13515
rect 21591 13481 21603 13515
rect 21545 13475 21603 13481
rect 21913 13515 21971 13521
rect 21913 13481 21925 13515
rect 21959 13512 21971 13515
rect 22646 13512 22652 13524
rect 21959 13484 22652 13512
rect 21959 13481 21971 13484
rect 21913 13475 21971 13481
rect 15194 13404 15200 13456
rect 15252 13444 15258 13456
rect 16298 13444 16304 13456
rect 15252 13416 16304 13444
rect 15252 13404 15258 13416
rect 16298 13404 16304 13416
rect 16356 13444 16362 13456
rect 17681 13447 17739 13453
rect 16356 13416 16804 13444
rect 16356 13404 16362 13416
rect 16666 13376 16672 13388
rect 16408 13348 16672 13376
rect 2869 13311 2927 13317
rect 2869 13277 2881 13311
rect 2915 13308 2927 13311
rect 9398 13308 9404 13320
rect 2915 13280 9404 13308
rect 2915 13277 2927 13280
rect 2869 13271 2927 13277
rect 9398 13268 9404 13280
rect 9456 13268 9462 13320
rect 10686 13268 10692 13320
rect 10744 13308 10750 13320
rect 12161 13311 12219 13317
rect 12161 13308 12173 13311
rect 10744 13280 12173 13308
rect 10744 13268 10750 13280
rect 12161 13277 12173 13280
rect 12207 13308 12219 13311
rect 12802 13308 12808 13320
rect 12207 13280 12808 13308
rect 12207 13277 12219 13280
rect 12161 13271 12219 13277
rect 12802 13268 12808 13280
rect 12860 13268 12866 13320
rect 16114 13308 16120 13320
rect 16027 13280 16120 13308
rect 16114 13268 16120 13280
rect 16172 13308 16178 13320
rect 16408 13317 16436 13348
rect 16666 13336 16672 13348
rect 16724 13336 16730 13388
rect 16393 13311 16451 13317
rect 16172 13280 16344 13308
rect 16172 13268 16178 13280
rect 16209 13243 16267 13249
rect 16209 13209 16221 13243
rect 16255 13209 16267 13243
rect 16316 13240 16344 13280
rect 16393 13277 16405 13311
rect 16439 13277 16451 13311
rect 16574 13308 16580 13320
rect 16535 13280 16580 13308
rect 16393 13271 16451 13277
rect 16574 13268 16580 13280
rect 16632 13268 16638 13320
rect 16776 13308 16804 13416
rect 17681 13413 17693 13447
rect 17727 13444 17739 13447
rect 17862 13444 17868 13456
rect 17727 13416 17868 13444
rect 17727 13413 17739 13416
rect 17681 13407 17739 13413
rect 17862 13404 17868 13416
rect 17920 13404 17926 13456
rect 16850 13336 16856 13388
rect 16908 13376 16914 13388
rect 17589 13379 17647 13385
rect 17589 13376 17601 13379
rect 16908 13348 17601 13376
rect 16908 13336 16914 13348
rect 17589 13345 17601 13348
rect 17635 13376 17647 13379
rect 20254 13376 20260 13388
rect 17635 13348 18000 13376
rect 20167 13348 20260 13376
rect 17635 13345 17647 13348
rect 17589 13339 17647 13345
rect 17865 13311 17923 13317
rect 17865 13308 17877 13311
rect 16776 13280 17877 13308
rect 17865 13277 17877 13280
rect 17911 13277 17923 13311
rect 17972 13308 18000 13348
rect 20254 13336 20260 13348
rect 20312 13376 20318 13388
rect 21560 13376 21588 13475
rect 22646 13472 22652 13484
rect 22704 13472 22710 13524
rect 24857 13515 24915 13521
rect 24857 13481 24869 13515
rect 24903 13512 24915 13515
rect 25130 13512 25136 13524
rect 24903 13484 25136 13512
rect 24903 13481 24915 13484
rect 24857 13475 24915 13481
rect 25130 13472 25136 13484
rect 25188 13512 25194 13524
rect 25409 13515 25467 13521
rect 25409 13512 25421 13515
rect 25188 13484 25421 13512
rect 25188 13472 25194 13484
rect 25409 13481 25421 13484
rect 25455 13481 25467 13515
rect 28166 13512 28172 13524
rect 28127 13484 28172 13512
rect 25409 13475 25467 13481
rect 28166 13472 28172 13484
rect 28224 13472 28230 13524
rect 28353 13515 28411 13521
rect 28353 13481 28365 13515
rect 28399 13512 28411 13515
rect 28902 13512 28908 13524
rect 28399 13484 28908 13512
rect 28399 13481 28411 13484
rect 28353 13475 28411 13481
rect 28902 13472 28908 13484
rect 28960 13472 28966 13524
rect 34701 13515 34759 13521
rect 34701 13481 34713 13515
rect 34747 13512 34759 13515
rect 34790 13512 34796 13524
rect 34747 13484 34796 13512
rect 34747 13481 34759 13484
rect 34701 13475 34759 13481
rect 34790 13472 34796 13484
rect 34848 13472 34854 13524
rect 36538 13512 36544 13524
rect 34900 13484 36544 13512
rect 33042 13444 33048 13456
rect 32048 13416 33048 13444
rect 22462 13376 22468 13388
rect 20312 13348 21588 13376
rect 22423 13348 22468 13376
rect 20312 13336 20318 13348
rect 22462 13336 22468 13348
rect 22520 13336 22526 13388
rect 25222 13376 25228 13388
rect 24872 13348 25228 13376
rect 20533 13311 20591 13317
rect 20533 13308 20545 13311
rect 17972 13280 20545 13308
rect 17865 13271 17923 13277
rect 20533 13277 20545 13280
rect 20579 13308 20591 13311
rect 20714 13308 20720 13320
rect 20579 13280 20720 13308
rect 20579 13277 20591 13280
rect 20533 13271 20591 13277
rect 20714 13268 20720 13280
rect 20772 13268 20778 13320
rect 21542 13308 21548 13320
rect 21503 13280 21548 13308
rect 21542 13268 21548 13280
rect 21600 13268 21606 13320
rect 21637 13311 21695 13317
rect 21637 13277 21649 13311
rect 21683 13277 21695 13311
rect 21637 13271 21695 13277
rect 16482 13240 16488 13252
rect 16316 13212 16488 13240
rect 16209 13203 16267 13209
rect 12342 13132 12348 13184
rect 12400 13172 12406 13184
rect 12713 13175 12771 13181
rect 12713 13172 12725 13175
rect 12400 13144 12725 13172
rect 12400 13132 12406 13144
rect 12713 13141 12725 13144
rect 12759 13141 12771 13175
rect 16224 13172 16252 13203
rect 16482 13200 16488 13212
rect 16540 13200 16546 13252
rect 16390 13172 16396 13184
rect 16224 13144 16396 13172
rect 12713 13135 12771 13141
rect 16390 13132 16396 13144
rect 16448 13132 16454 13184
rect 18046 13172 18052 13184
rect 18007 13144 18052 13172
rect 18046 13132 18052 13144
rect 18104 13132 18110 13184
rect 20530 13132 20536 13184
rect 20588 13172 20594 13184
rect 21652 13172 21680 13271
rect 22370 13268 22376 13320
rect 22428 13308 22434 13320
rect 22721 13311 22779 13317
rect 22721 13308 22733 13311
rect 22428 13280 22733 13308
rect 22428 13268 22434 13280
rect 22721 13277 22733 13280
rect 22767 13277 22779 13311
rect 24670 13308 24676 13320
rect 24631 13280 24676 13308
rect 22721 13271 22779 13277
rect 24670 13268 24676 13280
rect 24728 13268 24734 13320
rect 24872 13317 24900 13348
rect 25222 13336 25228 13348
rect 25280 13336 25286 13388
rect 25777 13379 25835 13385
rect 25777 13345 25789 13379
rect 25823 13345 25835 13379
rect 25777 13339 25835 13345
rect 29917 13379 29975 13385
rect 29917 13345 29929 13379
rect 29963 13376 29975 13379
rect 30282 13376 30288 13388
rect 29963 13348 30288 13376
rect 29963 13345 29975 13348
rect 29917 13339 29975 13345
rect 24857 13311 24915 13317
rect 24857 13277 24869 13311
rect 24903 13277 24915 13311
rect 25314 13308 25320 13320
rect 25275 13280 25320 13308
rect 24857 13271 24915 13277
rect 25314 13268 25320 13280
rect 25372 13268 25378 13320
rect 25792 13308 25820 13339
rect 30282 13336 30288 13348
rect 30340 13336 30346 13388
rect 32048 13385 32076 13416
rect 33042 13404 33048 13416
rect 33100 13444 33106 13456
rect 33100 13416 33548 13444
rect 33100 13404 33106 13416
rect 32033 13379 32091 13385
rect 32033 13345 32045 13379
rect 32079 13345 32091 13379
rect 33410 13376 33416 13388
rect 33371 13348 33416 13376
rect 32033 13339 32091 13345
rect 33410 13336 33416 13348
rect 33468 13336 33474 13388
rect 33520 13385 33548 13416
rect 33505 13379 33563 13385
rect 33505 13345 33517 13379
rect 33551 13345 33563 13379
rect 33505 13339 33563 13345
rect 26329 13311 26387 13317
rect 26329 13308 26341 13311
rect 25792 13280 26341 13308
rect 26329 13277 26341 13280
rect 26375 13277 26387 13311
rect 26329 13271 26387 13277
rect 28721 13311 28779 13317
rect 28721 13277 28733 13311
rect 28767 13308 28779 13311
rect 29270 13308 29276 13320
rect 28767 13280 29276 13308
rect 28767 13277 28779 13280
rect 28721 13271 28779 13277
rect 29270 13268 29276 13280
rect 29328 13268 29334 13320
rect 30098 13308 30104 13320
rect 30059 13280 30104 13308
rect 30098 13268 30104 13280
rect 30156 13268 30162 13320
rect 31018 13308 31024 13320
rect 30979 13280 31024 13308
rect 31018 13268 31024 13280
rect 31076 13268 31082 13320
rect 31389 13311 31447 13317
rect 31389 13277 31401 13311
rect 31435 13308 31447 13311
rect 32214 13308 32220 13320
rect 31435 13280 32220 13308
rect 31435 13277 31447 13280
rect 31389 13271 31447 13277
rect 32214 13268 32220 13280
rect 32272 13268 32278 13320
rect 33321 13311 33379 13317
rect 33321 13277 33333 13311
rect 33367 13308 33379 13311
rect 34330 13308 34336 13320
rect 33367 13280 34336 13308
rect 33367 13277 33379 13280
rect 33321 13271 33379 13277
rect 34330 13268 34336 13280
rect 34388 13268 34394 13320
rect 34514 13268 34520 13320
rect 34572 13308 34578 13320
rect 34701 13311 34759 13317
rect 34701 13308 34713 13311
rect 34572 13280 34713 13308
rect 34572 13268 34578 13280
rect 34701 13277 34713 13280
rect 34747 13277 34759 13311
rect 34701 13271 34759 13277
rect 27246 13240 27252 13252
rect 26528 13212 27252 13240
rect 20588 13144 21680 13172
rect 23845 13175 23903 13181
rect 20588 13132 20594 13144
rect 23845 13141 23857 13175
rect 23891 13172 23903 13175
rect 24210 13172 24216 13184
rect 23891 13144 24216 13172
rect 23891 13141 23903 13144
rect 23845 13135 23903 13141
rect 24210 13132 24216 13144
rect 24268 13132 24274 13184
rect 26528 13181 26556 13212
rect 27246 13200 27252 13212
rect 27304 13240 27310 13252
rect 30116 13240 30144 13268
rect 30282 13240 30288 13252
rect 27304 13212 30144 13240
rect 30243 13212 30288 13240
rect 27304 13200 27310 13212
rect 30282 13200 30288 13212
rect 30340 13200 30346 13252
rect 34900 13240 34928 13484
rect 36538 13472 36544 13484
rect 36596 13472 36602 13524
rect 36814 13512 36820 13524
rect 36775 13484 36820 13512
rect 36814 13472 36820 13484
rect 36872 13472 36878 13524
rect 35710 13404 35716 13456
rect 35768 13404 35774 13456
rect 35437 13379 35495 13385
rect 35437 13345 35449 13379
rect 35483 13376 35495 13379
rect 35728 13376 35756 13404
rect 41322 13376 41328 13388
rect 35483 13348 35756 13376
rect 41283 13348 41328 13376
rect 35483 13345 35495 13348
rect 35437 13339 35495 13345
rect 41322 13336 41328 13348
rect 41380 13336 41386 13388
rect 41782 13336 41788 13388
rect 41840 13376 41846 13388
rect 42153 13379 42211 13385
rect 42153 13376 42165 13379
rect 41840 13348 42165 13376
rect 41840 13336 41846 13348
rect 42153 13345 42165 13348
rect 42199 13345 42211 13379
rect 42153 13339 42211 13345
rect 34977 13311 35035 13317
rect 34977 13277 34989 13311
rect 35023 13277 35035 13311
rect 35710 13308 35716 13320
rect 35671 13280 35716 13308
rect 34977 13271 35035 13277
rect 31726 13212 34928 13240
rect 34992 13240 35020 13271
rect 35710 13268 35716 13280
rect 35768 13268 35774 13320
rect 36170 13268 36176 13320
rect 36228 13308 36234 13320
rect 36725 13311 36783 13317
rect 36725 13308 36737 13311
rect 36228 13280 36737 13308
rect 36228 13268 36234 13280
rect 36725 13277 36737 13280
rect 36771 13277 36783 13311
rect 36725 13271 36783 13277
rect 36909 13311 36967 13317
rect 36909 13277 36921 13311
rect 36955 13277 36967 13311
rect 37366 13308 37372 13320
rect 37327 13280 37372 13308
rect 36909 13271 36967 13277
rect 35342 13240 35348 13252
rect 34992 13212 35348 13240
rect 26513 13175 26571 13181
rect 26513 13141 26525 13175
rect 26559 13141 26571 13175
rect 28350 13172 28356 13184
rect 28311 13144 28356 13172
rect 26513 13135 26571 13141
rect 28350 13132 28356 13144
rect 28408 13132 28414 13184
rect 28442 13132 28448 13184
rect 28500 13172 28506 13184
rect 31726 13172 31754 13212
rect 35342 13200 35348 13212
rect 35400 13240 35406 13252
rect 35526 13240 35532 13252
rect 35400 13212 35532 13240
rect 35400 13200 35406 13212
rect 35526 13200 35532 13212
rect 35584 13200 35590 13252
rect 36262 13200 36268 13252
rect 36320 13240 36326 13252
rect 36924 13240 36952 13271
rect 37366 13268 37372 13280
rect 37424 13268 37430 13320
rect 36320 13212 36952 13240
rect 36320 13200 36326 13212
rect 41506 13200 41512 13252
rect 41564 13240 41570 13252
rect 41969 13243 42027 13249
rect 41969 13240 41981 13243
rect 41564 13212 41981 13240
rect 41564 13200 41570 13212
rect 41969 13209 41981 13212
rect 42015 13209 42027 13243
rect 41969 13203 42027 13209
rect 28500 13144 31754 13172
rect 28500 13132 28506 13144
rect 32306 13132 32312 13184
rect 32364 13172 32370 13184
rect 32953 13175 33011 13181
rect 32953 13172 32965 13175
rect 32364 13144 32965 13172
rect 32364 13132 32370 13144
rect 32953 13141 32965 13144
rect 32999 13141 33011 13175
rect 32953 13135 33011 13141
rect 34885 13175 34943 13181
rect 34885 13141 34897 13175
rect 34931 13172 34943 13175
rect 35250 13172 35256 13184
rect 34931 13144 35256 13172
rect 34931 13141 34943 13144
rect 34885 13135 34943 13141
rect 35250 13132 35256 13144
rect 35308 13172 35314 13184
rect 36170 13172 36176 13184
rect 35308 13144 36176 13172
rect 35308 13132 35314 13144
rect 36170 13132 36176 13144
rect 36228 13132 36234 13184
rect 37458 13172 37464 13184
rect 37419 13144 37464 13172
rect 37458 13132 37464 13144
rect 37516 13132 37522 13184
rect 1104 13082 42872 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 42872 13082
rect 1104 13008 42872 13030
rect 12802 12928 12808 12980
rect 12860 12968 12866 12980
rect 19705 12971 19763 12977
rect 12860 12940 19564 12968
rect 12860 12928 12866 12940
rect 12342 12900 12348 12912
rect 12303 12872 12348 12900
rect 12342 12860 12348 12872
rect 12400 12860 12406 12912
rect 15013 12903 15071 12909
rect 15013 12869 15025 12903
rect 15059 12900 15071 12903
rect 17218 12900 17224 12912
rect 15059 12872 17224 12900
rect 15059 12869 15071 12872
rect 15013 12863 15071 12869
rect 17218 12860 17224 12872
rect 17276 12860 17282 12912
rect 18046 12860 18052 12912
rect 18104 12900 18110 12912
rect 18570 12903 18628 12909
rect 18570 12900 18582 12903
rect 18104 12872 18582 12900
rect 18104 12860 18110 12872
rect 18570 12869 18582 12872
rect 18616 12869 18628 12903
rect 18570 12863 18628 12869
rect 15194 12832 15200 12844
rect 15155 12804 15200 12832
rect 15194 12792 15200 12804
rect 15252 12792 15258 12844
rect 15841 12835 15899 12841
rect 15841 12801 15853 12835
rect 15887 12832 15899 12835
rect 16117 12835 16175 12841
rect 15887 12804 16068 12832
rect 15887 12801 15899 12804
rect 15841 12795 15899 12801
rect 12161 12767 12219 12773
rect 12161 12733 12173 12767
rect 12207 12764 12219 12767
rect 12710 12764 12716 12776
rect 12207 12736 12716 12764
rect 12207 12733 12219 12736
rect 12161 12727 12219 12733
rect 12710 12724 12716 12736
rect 12768 12724 12774 12776
rect 13722 12764 13728 12776
rect 13683 12736 13728 12764
rect 13722 12724 13728 12736
rect 13780 12724 13786 12776
rect 15930 12764 15936 12776
rect 15891 12736 15936 12764
rect 15930 12724 15936 12736
rect 15988 12724 15994 12776
rect 16040 12764 16068 12804
rect 16117 12801 16129 12835
rect 16163 12832 16175 12835
rect 16298 12832 16304 12844
rect 16163 12804 16304 12832
rect 16163 12801 16175 12804
rect 16117 12795 16175 12801
rect 16298 12792 16304 12804
rect 16356 12792 16362 12844
rect 16482 12792 16488 12844
rect 16540 12832 16546 12844
rect 16669 12835 16727 12841
rect 16669 12832 16681 12835
rect 16540 12804 16681 12832
rect 16540 12792 16546 12804
rect 16669 12801 16681 12804
rect 16715 12832 16727 12835
rect 16715 12804 17908 12832
rect 16715 12801 16727 12804
rect 16669 12795 16727 12801
rect 16942 12764 16948 12776
rect 16040 12736 16948 12764
rect 16942 12724 16948 12736
rect 17000 12724 17006 12776
rect 17880 12764 17908 12804
rect 17954 12792 17960 12844
rect 18012 12832 18018 12844
rect 18325 12835 18383 12841
rect 18325 12832 18337 12835
rect 18012 12804 18337 12832
rect 18012 12792 18018 12804
rect 18325 12801 18337 12804
rect 18371 12801 18383 12835
rect 18325 12795 18383 12801
rect 18432 12804 19380 12832
rect 18432 12764 18460 12804
rect 17880 12736 18460 12764
rect 13814 12656 13820 12708
rect 13872 12696 13878 12708
rect 15657 12699 15715 12705
rect 15657 12696 15669 12699
rect 13872 12668 15669 12696
rect 13872 12656 13878 12668
rect 15657 12665 15669 12668
rect 15703 12665 15715 12699
rect 15657 12659 15715 12665
rect 16298 12656 16304 12708
rect 16356 12696 16362 12708
rect 19352 12696 19380 12804
rect 19536 12764 19564 12940
rect 19705 12937 19717 12971
rect 19751 12968 19763 12971
rect 20254 12968 20260 12980
rect 19751 12940 20260 12968
rect 19751 12937 19763 12940
rect 19705 12931 19763 12937
rect 20254 12928 20260 12940
rect 20312 12928 20318 12980
rect 21174 12968 21180 12980
rect 21087 12940 21180 12968
rect 21174 12928 21180 12940
rect 21232 12968 21238 12980
rect 21542 12968 21548 12980
rect 21232 12940 21548 12968
rect 21232 12928 21238 12940
rect 21542 12928 21548 12940
rect 21600 12928 21606 12980
rect 28442 12968 28448 12980
rect 23768 12940 28448 12968
rect 22005 12903 22063 12909
rect 22005 12900 22017 12903
rect 20916 12872 22017 12900
rect 20346 12792 20352 12844
rect 20404 12832 20410 12844
rect 20916 12841 20944 12872
rect 22005 12869 22017 12872
rect 22051 12869 22063 12903
rect 22005 12863 22063 12869
rect 20901 12835 20959 12841
rect 20901 12832 20913 12835
rect 20404 12804 20913 12832
rect 20404 12792 20410 12804
rect 20901 12801 20913 12804
rect 20947 12801 20959 12835
rect 20901 12795 20959 12801
rect 20993 12835 21051 12841
rect 20993 12801 21005 12835
rect 21039 12832 21051 12835
rect 21082 12832 21088 12844
rect 21039 12804 21088 12832
rect 21039 12801 21051 12804
rect 20993 12795 21051 12801
rect 21082 12792 21088 12804
rect 21140 12832 21146 12844
rect 21821 12835 21879 12841
rect 21821 12832 21833 12835
rect 21140 12804 21833 12832
rect 21140 12792 21146 12804
rect 21821 12801 21833 12804
rect 21867 12801 21879 12835
rect 21821 12795 21879 12801
rect 23768 12764 23796 12940
rect 28442 12928 28448 12940
rect 28500 12928 28506 12980
rect 29270 12968 29276 12980
rect 29231 12940 29276 12968
rect 29270 12928 29276 12940
rect 29328 12928 29334 12980
rect 30282 12968 30288 12980
rect 30195 12940 30288 12968
rect 30282 12928 30288 12940
rect 30340 12968 30346 12980
rect 32214 12968 32220 12980
rect 30340 12940 31432 12968
rect 32175 12940 32220 12968
rect 30340 12928 30346 12940
rect 26329 12903 26387 12909
rect 26329 12869 26341 12903
rect 26375 12900 26387 12903
rect 27522 12900 27528 12912
rect 26375 12872 27528 12900
rect 26375 12869 26387 12872
rect 26329 12863 26387 12869
rect 27522 12860 27528 12872
rect 27580 12900 27586 12912
rect 27580 12872 29224 12900
rect 27580 12860 27586 12872
rect 23934 12832 23940 12844
rect 23895 12804 23940 12832
rect 23934 12792 23940 12804
rect 23992 12792 23998 12844
rect 24210 12832 24216 12844
rect 24171 12804 24216 12832
rect 24210 12792 24216 12804
rect 24268 12832 24274 12844
rect 27246 12841 27252 12844
rect 25041 12835 25099 12841
rect 25041 12832 25053 12835
rect 24268 12804 25053 12832
rect 24268 12792 24274 12804
rect 25041 12801 25053 12804
rect 25087 12801 25099 12835
rect 27240 12832 27252 12841
rect 27207 12804 27252 12832
rect 25041 12795 25099 12801
rect 27240 12795 27252 12804
rect 27246 12792 27252 12795
rect 27304 12792 27310 12844
rect 28810 12832 28816 12844
rect 28771 12804 28816 12832
rect 28810 12792 28816 12804
rect 28868 12792 28874 12844
rect 29086 12832 29092 12844
rect 29047 12804 29092 12832
rect 29086 12792 29092 12804
rect 29144 12792 29150 12844
rect 24118 12764 24124 12776
rect 19536 12736 23796 12764
rect 24079 12736 24124 12764
rect 24118 12724 24124 12736
rect 24176 12724 24182 12776
rect 25130 12764 25136 12776
rect 25091 12736 25136 12764
rect 25130 12724 25136 12736
rect 25188 12724 25194 12776
rect 26970 12764 26976 12776
rect 26931 12736 26976 12764
rect 26970 12724 26976 12736
rect 27028 12724 27034 12776
rect 28994 12764 29000 12776
rect 28955 12736 29000 12764
rect 28994 12724 29000 12736
rect 29052 12724 29058 12776
rect 29196 12764 29224 12872
rect 30300 12841 30328 12928
rect 31297 12903 31355 12909
rect 31297 12900 31309 12903
rect 30392 12872 31309 12900
rect 30285 12835 30343 12841
rect 30285 12801 30297 12835
rect 30331 12801 30343 12835
rect 30285 12795 30343 12801
rect 30392 12764 30420 12872
rect 31297 12869 31309 12872
rect 31343 12869 31355 12903
rect 31404 12900 31432 12940
rect 32214 12928 32220 12940
rect 32272 12928 32278 12980
rect 33226 12928 33232 12980
rect 33284 12968 33290 12980
rect 33597 12971 33655 12977
rect 33597 12968 33609 12971
rect 33284 12940 33609 12968
rect 33284 12928 33290 12940
rect 33597 12937 33609 12940
rect 33643 12937 33655 12971
rect 33597 12931 33655 12937
rect 33778 12928 33784 12980
rect 33836 12968 33842 12980
rect 34057 12971 34115 12977
rect 34057 12968 34069 12971
rect 33836 12940 34069 12968
rect 33836 12928 33842 12940
rect 34057 12937 34069 12940
rect 34103 12937 34115 12971
rect 34057 12931 34115 12937
rect 34072 12900 34100 12931
rect 34698 12928 34704 12980
rect 34756 12968 34762 12980
rect 34885 12971 34943 12977
rect 34885 12968 34897 12971
rect 34756 12940 34897 12968
rect 34756 12928 34762 12940
rect 34885 12937 34897 12940
rect 34931 12937 34943 12971
rect 35529 12971 35587 12977
rect 35529 12968 35541 12971
rect 34885 12931 34943 12937
rect 34992 12940 35541 12968
rect 34992 12900 35020 12940
rect 35529 12937 35541 12940
rect 35575 12937 35587 12971
rect 35986 12968 35992 12980
rect 35947 12940 35992 12968
rect 35529 12931 35587 12937
rect 35986 12928 35992 12940
rect 36044 12928 36050 12980
rect 41506 12968 41512 12980
rect 41467 12940 41512 12968
rect 41506 12928 41512 12940
rect 41564 12928 41570 12980
rect 37458 12900 37464 12912
rect 31404 12872 32352 12900
rect 34072 12872 35020 12900
rect 35360 12872 37464 12900
rect 31297 12863 31355 12869
rect 30561 12835 30619 12841
rect 30561 12801 30573 12835
rect 30607 12801 30619 12835
rect 30742 12832 30748 12844
rect 30703 12804 30748 12832
rect 30561 12795 30619 12801
rect 29196 12736 30420 12764
rect 30576 12764 30604 12795
rect 30742 12792 30748 12804
rect 30800 12832 30806 12844
rect 31202 12832 31208 12844
rect 30800 12804 31208 12832
rect 30800 12792 30806 12804
rect 31202 12792 31208 12804
rect 31260 12792 31266 12844
rect 31478 12792 31484 12844
rect 31536 12832 31542 12844
rect 32324 12841 32352 12872
rect 32125 12835 32183 12841
rect 32125 12832 32137 12835
rect 31536 12804 32137 12832
rect 31536 12792 31542 12804
rect 32125 12801 32137 12804
rect 32171 12801 32183 12835
rect 32125 12795 32183 12801
rect 32309 12835 32367 12841
rect 32309 12801 32321 12835
rect 32355 12801 32367 12835
rect 32309 12795 32367 12801
rect 33965 12835 34023 12841
rect 33965 12801 33977 12835
rect 34011 12832 34023 12835
rect 34790 12832 34796 12844
rect 34011 12804 34796 12832
rect 34011 12801 34023 12804
rect 33965 12795 34023 12801
rect 34790 12792 34796 12804
rect 34848 12792 34854 12844
rect 35360 12841 35388 12872
rect 37458 12860 37464 12872
rect 37516 12860 37522 12912
rect 35345 12835 35403 12841
rect 35345 12801 35357 12835
rect 35391 12801 35403 12835
rect 35345 12795 35403 12801
rect 35710 12792 35716 12844
rect 35768 12832 35774 12844
rect 36127 12835 36185 12841
rect 36127 12832 36139 12835
rect 35768 12804 36139 12832
rect 35768 12792 35774 12804
rect 36127 12801 36139 12804
rect 36173 12801 36185 12835
rect 36262 12832 36268 12844
rect 36223 12804 36268 12832
rect 36127 12795 36185 12801
rect 36262 12792 36268 12804
rect 36320 12792 36326 12844
rect 36357 12835 36415 12841
rect 36357 12801 36369 12835
rect 36403 12801 36415 12835
rect 36485 12835 36543 12841
rect 36485 12832 36497 12835
rect 36357 12795 36415 12801
rect 36464 12801 36497 12832
rect 36531 12801 36543 12835
rect 36464 12795 36543 12801
rect 31018 12764 31024 12776
rect 30576 12736 31024 12764
rect 31018 12724 31024 12736
rect 31076 12724 31082 12776
rect 34241 12767 34299 12773
rect 34241 12733 34253 12767
rect 34287 12733 34299 12767
rect 35250 12764 35256 12776
rect 35211 12736 35256 12764
rect 34241 12727 34299 12733
rect 20530 12696 20536 12708
rect 16356 12668 16988 12696
rect 19352 12668 20536 12696
rect 16356 12656 16362 12668
rect 1670 12628 1676 12640
rect 1631 12600 1676 12628
rect 1670 12588 1676 12600
rect 1728 12588 1734 12640
rect 16117 12631 16175 12637
rect 16117 12597 16129 12631
rect 16163 12628 16175 12631
rect 16666 12628 16672 12640
rect 16163 12600 16672 12628
rect 16163 12597 16175 12600
rect 16117 12591 16175 12597
rect 16666 12588 16672 12600
rect 16724 12588 16730 12640
rect 16960 12628 16988 12668
rect 20530 12656 20536 12668
rect 20588 12656 20594 12708
rect 24670 12696 24676 12708
rect 24228 12668 24676 12696
rect 22186 12628 22192 12640
rect 16960 12600 22192 12628
rect 22186 12588 22192 12600
rect 22244 12588 22250 12640
rect 24228 12637 24256 12668
rect 24670 12656 24676 12668
rect 24728 12656 24734 12708
rect 26050 12656 26056 12708
rect 26108 12696 26114 12708
rect 26145 12699 26203 12705
rect 26145 12696 26157 12699
rect 26108 12668 26157 12696
rect 26108 12656 26114 12668
rect 26145 12665 26157 12668
rect 26191 12696 26203 12699
rect 26234 12696 26240 12708
rect 26191 12668 26240 12696
rect 26191 12665 26203 12668
rect 26145 12659 26203 12665
rect 26234 12656 26240 12668
rect 26292 12656 26298 12708
rect 30374 12696 30380 12708
rect 28276 12668 30380 12696
rect 24213 12631 24271 12637
rect 24213 12597 24225 12631
rect 24259 12597 24271 12631
rect 24394 12628 24400 12640
rect 24355 12600 24400 12628
rect 24213 12591 24271 12597
rect 24394 12588 24400 12600
rect 24452 12588 24458 12640
rect 25409 12631 25467 12637
rect 25409 12597 25421 12631
rect 25455 12628 25467 12631
rect 26326 12628 26332 12640
rect 25455 12600 26332 12628
rect 25455 12597 25467 12600
rect 25409 12591 25467 12597
rect 26326 12588 26332 12600
rect 26384 12588 26390 12640
rect 26970 12588 26976 12640
rect 27028 12628 27034 12640
rect 28276 12628 28304 12668
rect 30374 12656 30380 12668
rect 30432 12696 30438 12708
rect 30834 12696 30840 12708
rect 30432 12668 30840 12696
rect 30432 12656 30438 12668
rect 30834 12656 30840 12668
rect 30892 12696 30898 12708
rect 31481 12699 31539 12705
rect 31481 12696 31493 12699
rect 30892 12668 31493 12696
rect 30892 12656 30898 12668
rect 31481 12665 31493 12668
rect 31527 12665 31539 12699
rect 31481 12659 31539 12665
rect 27028 12600 28304 12628
rect 28353 12631 28411 12637
rect 27028 12588 27034 12600
rect 28353 12597 28365 12631
rect 28399 12628 28411 12631
rect 28813 12631 28871 12637
rect 28813 12628 28825 12631
rect 28399 12600 28825 12628
rect 28399 12597 28411 12600
rect 28353 12591 28411 12597
rect 28813 12597 28825 12600
rect 28859 12597 28871 12631
rect 28813 12591 28871 12597
rect 30466 12588 30472 12640
rect 30524 12628 30530 12640
rect 30561 12631 30619 12637
rect 30561 12628 30573 12631
rect 30524 12600 30573 12628
rect 30524 12588 30530 12600
rect 30561 12597 30573 12600
rect 30607 12597 30619 12631
rect 34256 12628 34284 12727
rect 35250 12724 35256 12736
rect 35308 12724 35314 12776
rect 35526 12724 35532 12776
rect 35584 12764 35590 12776
rect 36372 12764 36400 12795
rect 35584 12736 36400 12764
rect 35584 12724 35590 12736
rect 36354 12696 36360 12708
rect 35544 12668 36360 12696
rect 35544 12628 35572 12668
rect 36354 12656 36360 12668
rect 36412 12696 36418 12708
rect 36464 12696 36492 12795
rect 36630 12792 36636 12844
rect 36688 12832 36694 12844
rect 36688 12804 36733 12832
rect 36688 12792 36694 12804
rect 37182 12792 37188 12844
rect 37240 12832 37246 12844
rect 37829 12835 37887 12841
rect 37829 12832 37841 12835
rect 37240 12804 37841 12832
rect 37240 12792 37246 12804
rect 37829 12801 37841 12804
rect 37875 12801 37887 12835
rect 41414 12832 41420 12844
rect 41375 12804 41420 12832
rect 37829 12795 37887 12801
rect 41414 12792 41420 12804
rect 41472 12832 41478 12844
rect 41690 12832 41696 12844
rect 41472 12804 41696 12832
rect 41472 12792 41478 12804
rect 41690 12792 41696 12804
rect 41748 12792 41754 12844
rect 37645 12699 37703 12705
rect 37645 12696 37657 12699
rect 36412 12668 37657 12696
rect 36412 12656 36418 12668
rect 37645 12665 37657 12668
rect 37691 12665 37703 12699
rect 37645 12659 37703 12665
rect 40770 12628 40776 12640
rect 34256 12600 35572 12628
rect 40731 12600 40776 12628
rect 30561 12591 30619 12597
rect 40770 12588 40776 12600
rect 40828 12588 40834 12640
rect 1104 12538 42872 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 42872 12538
rect 1104 12464 42872 12486
rect 9398 12384 9404 12436
rect 9456 12424 9462 12436
rect 11698 12424 11704 12436
rect 9456 12396 11704 12424
rect 9456 12384 9462 12396
rect 11698 12384 11704 12396
rect 11756 12384 11762 12436
rect 12710 12424 12716 12436
rect 12671 12396 12716 12424
rect 12710 12384 12716 12396
rect 12768 12384 12774 12436
rect 15657 12427 15715 12433
rect 15657 12393 15669 12427
rect 15703 12424 15715 12427
rect 16114 12424 16120 12436
rect 15703 12396 16120 12424
rect 15703 12393 15715 12396
rect 15657 12387 15715 12393
rect 16114 12384 16120 12396
rect 16172 12384 16178 12436
rect 16209 12427 16267 12433
rect 16209 12393 16221 12427
rect 16255 12424 16267 12427
rect 16574 12424 16580 12436
rect 16255 12396 16580 12424
rect 16255 12393 16267 12396
rect 16209 12387 16267 12393
rect 16574 12384 16580 12396
rect 16632 12384 16638 12436
rect 17218 12424 17224 12436
rect 17179 12396 17224 12424
rect 17218 12384 17224 12396
rect 17276 12384 17282 12436
rect 20162 12424 20168 12436
rect 20123 12396 20168 12424
rect 20162 12384 20168 12396
rect 20220 12384 20226 12436
rect 20346 12424 20352 12436
rect 20307 12396 20352 12424
rect 20346 12384 20352 12396
rect 20404 12384 20410 12436
rect 24394 12424 24400 12436
rect 24355 12396 24400 12424
rect 24394 12384 24400 12396
rect 24452 12384 24458 12436
rect 24762 12424 24768 12436
rect 24723 12396 24768 12424
rect 24762 12384 24768 12396
rect 24820 12384 24826 12436
rect 27433 12427 27491 12433
rect 27433 12393 27445 12427
rect 27479 12424 27491 12427
rect 28810 12424 28816 12436
rect 27479 12396 28816 12424
rect 27479 12393 27491 12396
rect 27433 12387 27491 12393
rect 28810 12384 28816 12396
rect 28868 12384 28874 12436
rect 34698 12384 34704 12436
rect 34756 12424 34762 12436
rect 34885 12427 34943 12433
rect 34885 12424 34897 12427
rect 34756 12396 34897 12424
rect 34756 12384 34762 12396
rect 34885 12393 34897 12396
rect 34931 12393 34943 12427
rect 34885 12387 34943 12393
rect 17589 12359 17647 12365
rect 17589 12325 17601 12359
rect 17635 12356 17647 12359
rect 17862 12356 17868 12368
rect 17635 12328 17868 12356
rect 17635 12325 17647 12328
rect 17589 12319 17647 12325
rect 17862 12316 17868 12328
rect 17920 12316 17926 12368
rect 19334 12356 19340 12368
rect 19295 12328 19340 12356
rect 19334 12316 19340 12328
rect 19392 12316 19398 12368
rect 1397 12291 1455 12297
rect 1397 12257 1409 12291
rect 1443 12288 1455 12291
rect 1670 12288 1676 12300
rect 1443 12260 1676 12288
rect 1443 12257 1455 12260
rect 1397 12251 1455 12257
rect 1670 12248 1676 12260
rect 1728 12248 1734 12300
rect 2774 12248 2780 12300
rect 2832 12288 2838 12300
rect 2832 12260 2877 12288
rect 2832 12248 2838 12260
rect 14090 12248 14096 12300
rect 14148 12288 14154 12300
rect 14277 12291 14335 12297
rect 14277 12288 14289 12291
rect 14148 12260 14289 12288
rect 14148 12248 14154 12260
rect 14277 12257 14289 12260
rect 14323 12257 14335 12291
rect 20438 12288 20444 12300
rect 14277 12251 14335 12257
rect 19168 12260 20444 12288
rect 12897 12223 12955 12229
rect 12897 12189 12909 12223
rect 12943 12220 12955 12223
rect 13814 12220 13820 12232
rect 12943 12192 13820 12220
rect 12943 12189 12955 12192
rect 12897 12183 12955 12189
rect 13814 12180 13820 12192
rect 13872 12180 13878 12232
rect 16298 12180 16304 12232
rect 16356 12220 16362 12232
rect 16393 12223 16451 12229
rect 16393 12220 16405 12223
rect 16356 12192 16405 12220
rect 16356 12180 16362 12192
rect 16393 12189 16405 12192
rect 16439 12189 16451 12223
rect 16393 12183 16451 12189
rect 16942 12180 16948 12232
rect 17000 12220 17006 12232
rect 18233 12223 18291 12229
rect 18233 12220 18245 12223
rect 17000 12192 18245 12220
rect 17000 12180 17006 12192
rect 18233 12189 18245 12192
rect 18279 12189 18291 12223
rect 18233 12183 18291 12189
rect 18322 12180 18328 12232
rect 18380 12220 18386 12232
rect 18509 12223 18567 12229
rect 18509 12220 18521 12223
rect 18380 12192 18521 12220
rect 18380 12180 18386 12192
rect 18509 12189 18521 12192
rect 18555 12189 18567 12223
rect 18509 12183 18567 12189
rect 19168 12222 19196 12260
rect 20438 12248 20444 12260
rect 20496 12288 20502 12300
rect 20993 12291 21051 12297
rect 20993 12288 21005 12291
rect 20496 12260 21005 12288
rect 20496 12248 20502 12260
rect 20993 12257 21005 12260
rect 21039 12257 21051 12291
rect 28537 12291 28595 12297
rect 28537 12288 28549 12291
rect 20993 12251 21051 12257
rect 27172 12260 28549 12288
rect 19245 12223 19303 12229
rect 19245 12222 19257 12223
rect 19168 12194 19257 12222
rect 1581 12155 1639 12161
rect 1581 12121 1593 12155
rect 1627 12152 1639 12155
rect 2130 12152 2136 12164
rect 1627 12124 2136 12152
rect 1627 12121 1639 12124
rect 1581 12115 1639 12121
rect 2130 12112 2136 12124
rect 2188 12112 2194 12164
rect 14544 12155 14602 12161
rect 14544 12121 14556 12155
rect 14590 12152 14602 12155
rect 14734 12152 14740 12164
rect 14590 12124 14740 12152
rect 14590 12121 14602 12124
rect 14544 12115 14602 12121
rect 14734 12112 14740 12124
rect 14792 12112 14798 12164
rect 16577 12155 16635 12161
rect 16577 12121 16589 12155
rect 16623 12152 16635 12155
rect 17494 12152 17500 12164
rect 16623 12124 17500 12152
rect 16623 12121 16635 12124
rect 16577 12115 16635 12121
rect 17494 12112 17500 12124
rect 17552 12152 17558 12164
rect 18340 12152 18368 12180
rect 17552 12124 18368 12152
rect 18417 12155 18475 12161
rect 17552 12112 17558 12124
rect 18417 12121 18429 12155
rect 18463 12152 18475 12155
rect 19168 12152 19196 12194
rect 19245 12189 19257 12194
rect 19291 12189 19303 12223
rect 19429 12223 19487 12229
rect 19429 12220 19441 12223
rect 19245 12183 19303 12189
rect 19352 12192 19441 12220
rect 18463 12124 19196 12152
rect 18463 12121 18475 12124
rect 18417 12115 18475 12121
rect 16298 12044 16304 12096
rect 16356 12084 16362 12096
rect 17037 12087 17095 12093
rect 17037 12084 17049 12087
rect 16356 12056 17049 12084
rect 16356 12044 16362 12056
rect 17037 12053 17049 12056
rect 17083 12053 17095 12087
rect 17037 12047 17095 12053
rect 17221 12087 17279 12093
rect 17221 12053 17233 12087
rect 17267 12084 17279 12087
rect 18049 12087 18107 12093
rect 18049 12084 18061 12087
rect 17267 12056 18061 12084
rect 17267 12053 17279 12056
rect 17221 12047 17279 12053
rect 18049 12053 18061 12056
rect 18095 12053 18107 12087
rect 18049 12047 18107 12053
rect 19150 12044 19156 12096
rect 19208 12084 19214 12096
rect 19352 12084 19380 12192
rect 19429 12189 19441 12192
rect 19475 12189 19487 12223
rect 21174 12220 21180 12232
rect 21135 12192 21180 12220
rect 19429 12183 19487 12189
rect 21174 12180 21180 12192
rect 21232 12180 21238 12232
rect 21266 12180 21272 12232
rect 21324 12220 21330 12232
rect 24397 12223 24455 12229
rect 24397 12220 24409 12223
rect 21324 12192 24409 12220
rect 21324 12180 21330 12192
rect 24397 12189 24409 12192
rect 24443 12189 24455 12223
rect 24397 12183 24455 12189
rect 24581 12223 24639 12229
rect 24581 12189 24593 12223
rect 24627 12220 24639 12223
rect 25130 12220 25136 12232
rect 24627 12192 25136 12220
rect 24627 12189 24639 12192
rect 24581 12183 24639 12189
rect 25130 12180 25136 12192
rect 25188 12180 25194 12232
rect 26050 12220 26056 12232
rect 26011 12192 26056 12220
rect 26050 12180 26056 12192
rect 26108 12180 26114 12232
rect 26326 12229 26332 12232
rect 26320 12220 26332 12229
rect 26239 12192 26332 12220
rect 26320 12183 26332 12192
rect 26384 12220 26390 12232
rect 27172 12220 27200 12260
rect 28537 12257 28549 12260
rect 28583 12257 28595 12291
rect 28537 12251 28595 12257
rect 28997 12291 29055 12297
rect 28997 12257 29009 12291
rect 29043 12288 29055 12291
rect 30193 12291 30251 12297
rect 30193 12288 30205 12291
rect 29043 12260 30205 12288
rect 29043 12257 29055 12260
rect 28997 12251 29055 12257
rect 30193 12257 30205 12260
rect 30239 12257 30251 12291
rect 30193 12251 30251 12257
rect 31113 12291 31171 12297
rect 31113 12257 31125 12291
rect 31159 12288 31171 12291
rect 32493 12291 32551 12297
rect 32493 12288 32505 12291
rect 31159 12260 32505 12288
rect 31159 12257 31171 12260
rect 31113 12251 31171 12257
rect 32493 12257 32505 12260
rect 32539 12288 32551 12291
rect 33410 12288 33416 12300
rect 32539 12260 33416 12288
rect 32539 12257 32551 12260
rect 32493 12251 32551 12257
rect 33410 12248 33416 12260
rect 33468 12248 33474 12300
rect 33594 12248 33600 12300
rect 33652 12288 33658 12300
rect 33873 12291 33931 12297
rect 33873 12288 33885 12291
rect 33652 12260 33885 12288
rect 33652 12248 33658 12260
rect 33873 12257 33885 12260
rect 33919 12257 33931 12291
rect 33873 12251 33931 12257
rect 34149 12291 34207 12297
rect 34149 12257 34161 12291
rect 34195 12288 34207 12291
rect 34514 12288 34520 12300
rect 34195 12260 34520 12288
rect 34195 12257 34207 12260
rect 34149 12251 34207 12257
rect 28626 12220 28632 12232
rect 26384 12192 27200 12220
rect 28587 12192 28632 12220
rect 26326 12180 26332 12183
rect 26384 12180 26390 12192
rect 28626 12180 28632 12192
rect 28684 12180 28690 12232
rect 30466 12220 30472 12232
rect 30427 12192 30472 12220
rect 30466 12180 30472 12192
rect 30524 12180 30530 12232
rect 32306 12220 32312 12232
rect 32267 12192 32312 12220
rect 32306 12180 32312 12192
rect 32364 12180 32370 12232
rect 32401 12223 32459 12229
rect 32401 12189 32413 12223
rect 32447 12220 32459 12223
rect 32858 12220 32864 12232
rect 32447 12192 32864 12220
rect 32447 12189 32459 12192
rect 32401 12183 32459 12189
rect 32858 12180 32864 12192
rect 32916 12180 32922 12232
rect 33888 12220 33916 12251
rect 34514 12248 34520 12260
rect 34572 12248 34578 12300
rect 34790 12248 34796 12300
rect 34848 12288 34854 12300
rect 36909 12291 36967 12297
rect 36909 12288 36921 12291
rect 34848 12260 36921 12288
rect 34848 12248 34854 12260
rect 33888 12192 34836 12220
rect 20530 12152 20536 12164
rect 20491 12124 20536 12152
rect 20530 12112 20536 12124
rect 20588 12112 20594 12164
rect 19208 12056 19380 12084
rect 20333 12087 20391 12093
rect 19208 12044 19214 12056
rect 20333 12053 20345 12087
rect 20379 12084 20391 12087
rect 20990 12084 20996 12096
rect 20379 12056 20996 12084
rect 20379 12053 20391 12056
rect 20333 12047 20391 12053
rect 20990 12044 20996 12056
rect 21048 12084 21054 12096
rect 21634 12084 21640 12096
rect 21048 12056 21640 12084
rect 21048 12044 21054 12056
rect 21634 12044 21640 12056
rect 21692 12044 21698 12096
rect 31938 12084 31944 12096
rect 31899 12056 31944 12084
rect 31938 12044 31944 12056
rect 31996 12044 32002 12096
rect 33502 12044 33508 12096
rect 33560 12084 33566 12096
rect 34701 12087 34759 12093
rect 34701 12084 34713 12087
rect 33560 12056 34713 12084
rect 33560 12044 33566 12056
rect 34701 12053 34713 12056
rect 34747 12053 34759 12087
rect 34808 12084 34836 12192
rect 34869 12155 34927 12161
rect 34869 12121 34881 12155
rect 34915 12152 34927 12155
rect 34992 12152 35020 12260
rect 36909 12257 36921 12260
rect 36955 12257 36967 12291
rect 36909 12251 36967 12257
rect 40313 12291 40371 12297
rect 40313 12257 40325 12291
rect 40359 12288 40371 12291
rect 40770 12288 40776 12300
rect 40359 12260 40776 12288
rect 40359 12257 40371 12260
rect 40313 12251 40371 12257
rect 40770 12248 40776 12260
rect 40828 12248 40834 12300
rect 42150 12288 42156 12300
rect 42111 12260 42156 12288
rect 42150 12248 42156 12260
rect 42208 12248 42214 12300
rect 35989 12223 36047 12229
rect 35989 12189 36001 12223
rect 36035 12220 36047 12223
rect 36078 12220 36084 12232
rect 36035 12192 36084 12220
rect 36035 12189 36047 12192
rect 35989 12183 36047 12189
rect 36078 12180 36084 12192
rect 36136 12180 36142 12232
rect 36817 12223 36875 12229
rect 36817 12220 36829 12223
rect 36372 12192 36829 12220
rect 34915 12124 35020 12152
rect 35069 12155 35127 12161
rect 34915 12121 34927 12124
rect 34869 12115 34927 12121
rect 35069 12121 35081 12155
rect 35115 12121 35127 12155
rect 35069 12115 35127 12121
rect 35084 12084 35112 12115
rect 35618 12112 35624 12164
rect 35676 12152 35682 12164
rect 35802 12152 35808 12164
rect 35676 12124 35808 12152
rect 35676 12112 35682 12124
rect 35802 12112 35808 12124
rect 35860 12112 35866 12164
rect 36173 12155 36231 12161
rect 36173 12121 36185 12155
rect 36219 12152 36231 12155
rect 36262 12152 36268 12164
rect 36219 12124 36268 12152
rect 36219 12121 36231 12124
rect 36173 12115 36231 12121
rect 36262 12112 36268 12124
rect 36320 12112 36326 12164
rect 36372 12096 36400 12192
rect 36817 12189 36829 12192
rect 36863 12189 36875 12223
rect 36998 12220 37004 12232
rect 36959 12192 37004 12220
rect 36817 12183 36875 12189
rect 36998 12180 37004 12192
rect 37056 12180 37062 12232
rect 40497 12155 40555 12161
rect 40497 12121 40509 12155
rect 40543 12152 40555 12155
rect 41506 12152 41512 12164
rect 40543 12124 41512 12152
rect 40543 12121 40555 12124
rect 40497 12115 40555 12121
rect 41506 12112 41512 12124
rect 41564 12112 41570 12164
rect 34808 12056 35112 12084
rect 34701 12047 34759 12053
rect 35158 12044 35164 12096
rect 35216 12084 35222 12096
rect 35986 12084 35992 12096
rect 35216 12056 35992 12084
rect 35216 12044 35222 12056
rect 35986 12044 35992 12056
rect 36044 12044 36050 12096
rect 36354 12084 36360 12096
rect 36315 12056 36360 12084
rect 36354 12044 36360 12056
rect 36412 12044 36418 12096
rect 1104 11994 42872 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 42872 11994
rect 1104 11920 42872 11942
rect 2130 11880 2136 11892
rect 2091 11852 2136 11880
rect 2130 11840 2136 11852
rect 2188 11840 2194 11892
rect 14734 11880 14740 11892
rect 14695 11852 14740 11880
rect 14734 11840 14740 11852
rect 14792 11840 14798 11892
rect 16761 11883 16819 11889
rect 16761 11849 16773 11883
rect 16807 11880 16819 11883
rect 17218 11880 17224 11892
rect 16807 11852 17224 11880
rect 16807 11849 16819 11852
rect 16761 11843 16819 11849
rect 17218 11840 17224 11852
rect 17276 11840 17282 11892
rect 19889 11883 19947 11889
rect 19889 11849 19901 11883
rect 19935 11880 19947 11883
rect 20346 11880 20352 11892
rect 19935 11852 20352 11880
rect 19935 11849 19947 11852
rect 19889 11843 19947 11849
rect 2225 11747 2283 11753
rect 2225 11713 2237 11747
rect 2271 11744 2283 11747
rect 2314 11744 2320 11756
rect 2271 11716 2320 11744
rect 2271 11713 2283 11716
rect 2225 11707 2283 11713
rect 2314 11704 2320 11716
rect 2372 11704 2378 11756
rect 9398 11744 9404 11756
rect 9359 11716 9404 11744
rect 9398 11704 9404 11716
rect 9456 11704 9462 11756
rect 14921 11747 14979 11753
rect 14921 11713 14933 11747
rect 14967 11744 14979 11747
rect 16298 11744 16304 11756
rect 14967 11716 16304 11744
rect 14967 11713 14979 11716
rect 14921 11707 14979 11713
rect 16298 11704 16304 11716
rect 16356 11704 16362 11756
rect 16482 11704 16488 11756
rect 16540 11744 16546 11756
rect 16945 11747 17003 11753
rect 16945 11744 16957 11747
rect 16540 11716 16957 11744
rect 16540 11704 16546 11716
rect 16945 11713 16957 11716
rect 16991 11713 17003 11747
rect 17236 11744 17264 11840
rect 19061 11815 19119 11821
rect 19061 11781 19073 11815
rect 19107 11781 19119 11815
rect 19061 11775 19119 11781
rect 19277 11815 19335 11821
rect 19277 11781 19289 11815
rect 19323 11812 19335 11815
rect 19518 11812 19524 11824
rect 19323 11784 19524 11812
rect 19323 11781 19335 11784
rect 19277 11775 19335 11781
rect 17681 11747 17739 11753
rect 17681 11744 17693 11747
rect 17236 11716 17693 11744
rect 16945 11707 17003 11713
rect 17681 11713 17693 11716
rect 17727 11713 17739 11747
rect 17681 11707 17739 11713
rect 17129 11679 17187 11685
rect 17129 11645 17141 11679
rect 17175 11645 17187 11679
rect 17129 11639 17187 11645
rect 17957 11679 18015 11685
rect 17957 11645 17969 11679
rect 18003 11676 18015 11679
rect 18230 11676 18236 11688
rect 18003 11648 18236 11676
rect 18003 11645 18015 11648
rect 17957 11639 18015 11645
rect 17144 11608 17172 11639
rect 18230 11636 18236 11648
rect 18288 11676 18294 11688
rect 19076 11676 19104 11775
rect 19518 11772 19524 11784
rect 19576 11772 19582 11824
rect 19702 11772 19708 11824
rect 19760 11812 19766 11824
rect 19904 11812 19932 11843
rect 20346 11840 20352 11852
rect 20404 11840 20410 11892
rect 23845 11883 23903 11889
rect 23845 11849 23857 11883
rect 23891 11880 23903 11883
rect 23934 11880 23940 11892
rect 23891 11852 23940 11880
rect 23891 11849 23903 11852
rect 23845 11843 23903 11849
rect 23934 11840 23940 11852
rect 23992 11840 23998 11892
rect 24118 11840 24124 11892
rect 24176 11880 24182 11892
rect 24305 11883 24363 11889
rect 24305 11880 24317 11883
rect 24176 11852 24317 11880
rect 24176 11840 24182 11852
rect 24305 11849 24317 11852
rect 24351 11849 24363 11883
rect 24305 11843 24363 11849
rect 28353 11883 28411 11889
rect 28353 11849 28365 11883
rect 28399 11880 28411 11883
rect 29086 11880 29092 11892
rect 28399 11852 29092 11880
rect 28399 11849 28411 11852
rect 28353 11843 28411 11849
rect 29086 11840 29092 11852
rect 29144 11840 29150 11892
rect 36170 11880 36176 11892
rect 35084 11852 36176 11880
rect 19760 11784 19932 11812
rect 19760 11772 19766 11784
rect 27154 11772 27160 11824
rect 27212 11821 27218 11824
rect 27212 11815 27276 11821
rect 27212 11781 27230 11815
rect 27264 11781 27276 11815
rect 27212 11775 27276 11781
rect 27212 11772 27218 11775
rect 33594 11772 33600 11824
rect 33652 11812 33658 11824
rect 34422 11812 34428 11824
rect 33652 11784 34428 11812
rect 33652 11772 33658 11784
rect 34422 11772 34428 11784
rect 34480 11772 34486 11824
rect 34974 11812 34980 11824
rect 34532 11784 34980 11812
rect 21013 11747 21071 11753
rect 21013 11713 21025 11747
rect 21059 11744 21071 11747
rect 21174 11744 21180 11756
rect 21059 11716 21180 11744
rect 21059 11713 21071 11716
rect 21013 11707 21071 11713
rect 21174 11704 21180 11716
rect 21232 11704 21238 11756
rect 21269 11747 21327 11753
rect 21269 11713 21281 11747
rect 21315 11744 21327 11747
rect 22462 11744 22468 11756
rect 21315 11716 22468 11744
rect 21315 11713 21327 11716
rect 21269 11707 21327 11713
rect 22462 11704 22468 11716
rect 22520 11704 22526 11756
rect 22554 11704 22560 11756
rect 22612 11744 22618 11756
rect 22721 11747 22779 11753
rect 22721 11744 22733 11747
rect 22612 11716 22733 11744
rect 22612 11704 22618 11716
rect 22721 11713 22733 11716
rect 22767 11713 22779 11747
rect 22721 11707 22779 11713
rect 23474 11704 23480 11756
rect 23532 11744 23538 11756
rect 25418 11747 25476 11753
rect 25418 11744 25430 11747
rect 23532 11716 25430 11744
rect 23532 11704 23538 11716
rect 25418 11713 25430 11716
rect 25464 11713 25476 11747
rect 26970 11744 26976 11756
rect 26931 11716 26976 11744
rect 25418 11707 25476 11713
rect 26970 11704 26976 11716
rect 27028 11704 27034 11756
rect 30653 11747 30711 11753
rect 30653 11713 30665 11747
rect 30699 11744 30711 11747
rect 31938 11744 31944 11756
rect 30699 11716 31944 11744
rect 30699 11713 30711 11716
rect 30653 11707 30711 11713
rect 31938 11704 31944 11716
rect 31996 11704 32002 11756
rect 33042 11704 33048 11756
rect 33100 11744 33106 11756
rect 33413 11747 33471 11753
rect 33413 11744 33425 11747
rect 33100 11716 33425 11744
rect 33100 11704 33106 11716
rect 33413 11713 33425 11716
rect 33459 11713 33471 11747
rect 33686 11744 33692 11756
rect 33647 11716 33692 11744
rect 33413 11707 33471 11713
rect 33686 11704 33692 11716
rect 33744 11704 33750 11756
rect 33873 11747 33931 11753
rect 33873 11713 33885 11747
rect 33919 11744 33931 11747
rect 34333 11747 34391 11753
rect 34333 11744 34345 11747
rect 33919 11716 34345 11744
rect 33919 11713 33931 11716
rect 33873 11707 33931 11713
rect 34333 11713 34345 11716
rect 34379 11744 34391 11747
rect 34532 11744 34560 11784
rect 34974 11772 34980 11784
rect 35032 11772 35038 11824
rect 35084 11775 35112 11852
rect 36170 11840 36176 11852
rect 36228 11880 36234 11892
rect 36998 11880 37004 11892
rect 36228 11852 37004 11880
rect 36228 11840 36234 11852
rect 36998 11840 37004 11852
rect 37056 11840 37062 11892
rect 41506 11880 41512 11892
rect 41467 11852 41512 11880
rect 41506 11840 41512 11852
rect 41564 11840 41570 11892
rect 36078 11812 36084 11824
rect 35820 11784 36084 11812
rect 35070 11769 35128 11775
rect 34379 11716 34560 11744
rect 34379 11713 34391 11716
rect 34333 11707 34391 11713
rect 34606 11704 34612 11756
rect 34664 11744 34670 11756
rect 34664 11716 34709 11744
rect 35070 11735 35082 11769
rect 35116 11735 35128 11769
rect 35820 11753 35848 11784
rect 36078 11772 36084 11784
rect 36136 11772 36142 11824
rect 35070 11729 35128 11735
rect 35805 11747 35863 11753
rect 34664 11704 34670 11716
rect 35805 11713 35817 11747
rect 35851 11713 35863 11747
rect 35805 11707 35863 11713
rect 36262 11704 36268 11756
rect 36320 11744 36326 11756
rect 36998 11744 37004 11756
rect 36320 11716 37004 11744
rect 36320 11704 36326 11716
rect 36998 11704 37004 11716
rect 37056 11704 37062 11756
rect 41414 11704 41420 11756
rect 41472 11744 41478 11756
rect 41601 11747 41659 11753
rect 41601 11744 41613 11747
rect 41472 11716 41613 11744
rect 41472 11704 41478 11716
rect 41601 11713 41613 11716
rect 41647 11713 41659 11747
rect 41601 11707 41659 11713
rect 18288 11648 19104 11676
rect 25685 11679 25743 11685
rect 18288 11636 18294 11648
rect 25685 11645 25697 11679
rect 25731 11676 25743 11679
rect 26050 11676 26056 11688
rect 25731 11648 26056 11676
rect 25731 11645 25743 11648
rect 25685 11639 25743 11645
rect 17144 11580 20024 11608
rect 9214 11500 9220 11552
rect 9272 11540 9278 11552
rect 9309 11543 9367 11549
rect 9309 11540 9321 11543
rect 9272 11512 9321 11540
rect 9272 11500 9278 11512
rect 9309 11509 9321 11512
rect 9355 11509 9367 11543
rect 9309 11503 9367 11509
rect 19245 11543 19303 11549
rect 19245 11509 19257 11543
rect 19291 11540 19303 11543
rect 19334 11540 19340 11552
rect 19291 11512 19340 11540
rect 19291 11509 19303 11512
rect 19245 11503 19303 11509
rect 19334 11500 19340 11512
rect 19392 11500 19398 11552
rect 19426 11500 19432 11552
rect 19484 11540 19490 11552
rect 19996 11540 20024 11580
rect 24578 11540 24584 11552
rect 19484 11512 19529 11540
rect 19996 11512 24584 11540
rect 19484 11500 19490 11512
rect 24578 11500 24584 11512
rect 24636 11500 24642 11552
rect 25314 11500 25320 11552
rect 25372 11540 25378 11552
rect 25700 11540 25728 11639
rect 26050 11636 26056 11648
rect 26108 11636 26114 11688
rect 34624 11676 34652 11704
rect 35345 11679 35403 11685
rect 35345 11676 35357 11679
rect 34624 11648 35357 11676
rect 35345 11645 35357 11648
rect 35391 11645 35403 11679
rect 35345 11639 35403 11645
rect 35986 11636 35992 11688
rect 36044 11676 36050 11688
rect 36081 11679 36139 11685
rect 36081 11676 36093 11679
rect 36044 11648 36093 11676
rect 36044 11636 36050 11648
rect 36081 11645 36093 11648
rect 36127 11676 36139 11679
rect 36814 11676 36820 11688
rect 36127 11648 36820 11676
rect 36127 11645 36139 11648
rect 36081 11639 36139 11645
rect 36814 11636 36820 11648
rect 36872 11636 36878 11688
rect 35161 11611 35219 11617
rect 35161 11577 35173 11611
rect 35207 11608 35219 11611
rect 35618 11608 35624 11620
rect 35207 11580 35624 11608
rect 35207 11577 35219 11580
rect 35161 11571 35219 11577
rect 35618 11568 35624 11580
rect 35676 11608 35682 11620
rect 36262 11608 36268 11620
rect 35676 11580 36268 11608
rect 35676 11568 35682 11580
rect 36262 11568 36268 11580
rect 36320 11568 36326 11620
rect 30466 11540 30472 11552
rect 25372 11512 25728 11540
rect 30427 11512 30472 11540
rect 25372 11500 25378 11512
rect 30466 11500 30472 11512
rect 30524 11500 30530 11552
rect 33226 11540 33232 11552
rect 33187 11512 33232 11540
rect 33226 11500 33232 11512
rect 33284 11500 33290 11552
rect 34330 11540 34336 11552
rect 34291 11512 34336 11540
rect 34330 11500 34336 11512
rect 34388 11500 34394 11552
rect 35253 11543 35311 11549
rect 35253 11509 35265 11543
rect 35299 11540 35311 11543
rect 35986 11540 35992 11552
rect 35299 11512 35992 11540
rect 35299 11509 35311 11512
rect 35253 11503 35311 11509
rect 35986 11500 35992 11512
rect 36044 11500 36050 11552
rect 40310 11500 40316 11552
rect 40368 11540 40374 11552
rect 40773 11543 40831 11549
rect 40773 11540 40785 11543
rect 40368 11512 40785 11540
rect 40368 11500 40374 11512
rect 40773 11509 40785 11512
rect 40819 11509 40831 11543
rect 40773 11503 40831 11509
rect 1104 11450 42872 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 42872 11450
rect 1104 11376 42872 11398
rect 19518 11336 19524 11348
rect 19479 11308 19524 11336
rect 19518 11296 19524 11308
rect 19576 11296 19582 11348
rect 20990 11336 20996 11348
rect 20951 11308 20996 11336
rect 20990 11296 20996 11308
rect 21048 11296 21054 11348
rect 21174 11296 21180 11348
rect 21232 11336 21238 11348
rect 21637 11339 21695 11345
rect 21637 11336 21649 11339
rect 21232 11308 21649 11336
rect 21232 11296 21238 11308
rect 21637 11305 21649 11308
rect 21683 11305 21695 11339
rect 22830 11336 22836 11348
rect 22743 11308 22836 11336
rect 21637 11299 21695 11305
rect 22830 11296 22836 11308
rect 22888 11336 22894 11348
rect 24026 11336 24032 11348
rect 22888 11308 24032 11336
rect 22888 11296 22894 11308
rect 24026 11296 24032 11308
rect 24084 11296 24090 11348
rect 36817 11339 36875 11345
rect 36817 11336 36829 11339
rect 35912 11308 36829 11336
rect 35912 11280 35940 11308
rect 36817 11305 36829 11308
rect 36863 11305 36875 11339
rect 36817 11299 36875 11305
rect 33873 11271 33931 11277
rect 33873 11237 33885 11271
rect 33919 11268 33931 11271
rect 35894 11268 35900 11280
rect 33919 11240 35900 11268
rect 33919 11237 33931 11240
rect 33873 11231 33931 11237
rect 35894 11228 35900 11240
rect 35952 11228 35958 11280
rect 36354 11268 36360 11280
rect 36096 11240 36360 11268
rect 19426 11160 19432 11212
rect 19484 11200 19490 11212
rect 19484 11172 21864 11200
rect 19484 11160 19490 11172
rect 1670 11132 1676 11144
rect 1631 11104 1676 11132
rect 1670 11092 1676 11104
rect 1728 11092 1734 11144
rect 17218 11132 17224 11144
rect 17179 11104 17224 11132
rect 17218 11092 17224 11104
rect 17276 11092 17282 11144
rect 17494 11092 17500 11144
rect 17552 11132 17558 11144
rect 17773 11135 17831 11141
rect 17773 11132 17785 11135
rect 17552 11104 17785 11132
rect 17552 11092 17558 11104
rect 17773 11101 17785 11104
rect 17819 11101 17831 11135
rect 17773 11095 17831 11101
rect 18049 11135 18107 11141
rect 18049 11101 18061 11135
rect 18095 11132 18107 11135
rect 18506 11132 18512 11144
rect 18095 11104 18512 11132
rect 18095 11101 18107 11104
rect 18049 11095 18107 11101
rect 18506 11092 18512 11104
rect 18564 11092 18570 11144
rect 19702 11132 19708 11144
rect 19663 11104 19708 11132
rect 19702 11092 19708 11104
rect 19760 11092 19766 11144
rect 19981 11135 20039 11141
rect 19981 11101 19993 11135
rect 20027 11101 20039 11135
rect 21082 11132 21088 11144
rect 21043 11104 21088 11132
rect 19981 11095 20039 11101
rect 18524 11064 18552 11092
rect 19150 11064 19156 11076
rect 18524 11036 19156 11064
rect 19150 11024 19156 11036
rect 19208 11064 19214 11076
rect 19996 11064 20024 11095
rect 21082 11092 21088 11104
rect 21140 11092 21146 11144
rect 21836 11141 21864 11172
rect 33686 11160 33692 11212
rect 33744 11200 33750 11212
rect 36096 11209 36124 11240
rect 36354 11228 36360 11240
rect 36412 11228 36418 11280
rect 36446 11228 36452 11280
rect 36504 11268 36510 11280
rect 36504 11240 37688 11268
rect 36504 11228 36510 11240
rect 33965 11203 34023 11209
rect 33965 11200 33977 11203
rect 33744 11172 33977 11200
rect 33744 11160 33750 11172
rect 33965 11169 33977 11172
rect 34011 11200 34023 11203
rect 34701 11203 34759 11209
rect 34701 11200 34713 11203
rect 34011 11172 34713 11200
rect 34011 11169 34023 11172
rect 33965 11163 34023 11169
rect 34701 11169 34713 11172
rect 34747 11169 34759 11203
rect 34701 11163 34759 11169
rect 36081 11203 36139 11209
rect 36081 11169 36093 11203
rect 36127 11169 36139 11203
rect 36081 11163 36139 11169
rect 36170 11160 36176 11212
rect 36228 11200 36234 11212
rect 36228 11172 36273 11200
rect 36228 11160 36234 11172
rect 21821 11135 21879 11141
rect 21821 11101 21833 11135
rect 21867 11101 21879 11135
rect 21821 11095 21879 11101
rect 22186 11092 22192 11144
rect 22244 11132 22250 11144
rect 22649 11135 22707 11141
rect 22649 11132 22661 11135
rect 22244 11104 22661 11132
rect 22244 11092 22250 11104
rect 22649 11101 22661 11104
rect 22695 11132 22707 11135
rect 23382 11132 23388 11144
rect 22695 11104 23388 11132
rect 22695 11101 22707 11104
rect 22649 11095 22707 11101
rect 23382 11092 23388 11104
rect 23440 11092 23446 11144
rect 25774 11092 25780 11144
rect 25832 11132 25838 11144
rect 26329 11135 26387 11141
rect 26329 11132 26341 11135
rect 25832 11104 26341 11132
rect 25832 11092 25838 11104
rect 26329 11101 26341 11104
rect 26375 11101 26387 11135
rect 33502 11132 33508 11144
rect 33463 11104 33508 11132
rect 26329 11095 26387 11101
rect 33502 11092 33508 11104
rect 33560 11092 33566 11144
rect 34422 11092 34428 11144
rect 34480 11132 34486 11144
rect 34885 11135 34943 11141
rect 34885 11132 34897 11135
rect 34480 11104 34897 11132
rect 34480 11092 34486 11104
rect 34885 11101 34897 11104
rect 34931 11101 34943 11135
rect 34885 11095 34943 11101
rect 35069 11135 35127 11141
rect 35069 11101 35081 11135
rect 35115 11132 35127 11135
rect 35434 11132 35440 11144
rect 35115 11104 35440 11132
rect 35115 11101 35127 11104
rect 35069 11095 35127 11101
rect 35434 11092 35440 11104
rect 35492 11132 35498 11144
rect 35710 11132 35716 11144
rect 35492 11104 35716 11132
rect 35492 11092 35498 11104
rect 35710 11092 35716 11104
rect 35768 11092 35774 11144
rect 35986 11132 35992 11144
rect 35947 11104 35992 11132
rect 35986 11092 35992 11104
rect 36044 11092 36050 11144
rect 36188 11132 36216 11160
rect 36446 11132 36452 11144
rect 36188 11104 36452 11132
rect 36446 11092 36452 11104
rect 36504 11092 36510 11144
rect 36814 11132 36820 11144
rect 36775 11104 36820 11132
rect 36814 11092 36820 11104
rect 36872 11092 36878 11144
rect 36998 11132 37004 11144
rect 36959 11104 37004 11132
rect 36998 11092 37004 11104
rect 37056 11092 37062 11144
rect 37660 11141 37688 11240
rect 40310 11200 40316 11212
rect 40271 11172 40316 11200
rect 40310 11160 40316 11172
rect 40368 11160 40374 11212
rect 37461 11135 37519 11141
rect 37461 11101 37473 11135
rect 37507 11101 37519 11135
rect 37461 11095 37519 11101
rect 37645 11135 37703 11141
rect 37645 11101 37657 11135
rect 37691 11101 37703 11135
rect 37645 11095 37703 11101
rect 20990 11064 20996 11076
rect 19208 11036 20024 11064
rect 20364 11036 20996 11064
rect 19208 11024 19214 11036
rect 14550 10956 14556 11008
rect 14608 10996 14614 11008
rect 17126 10996 17132 11008
rect 14608 10968 17132 10996
rect 14608 10956 14614 10968
rect 17126 10956 17132 10968
rect 17184 10956 17190 11008
rect 17310 10956 17316 11008
rect 17368 10996 17374 11008
rect 19242 10996 19248 11008
rect 17368 10968 19248 10996
rect 17368 10956 17374 10968
rect 19242 10956 19248 10968
rect 19300 10956 19306 11008
rect 19426 10956 19432 11008
rect 19484 10996 19490 11008
rect 19889 10999 19947 11005
rect 19889 10996 19901 10999
rect 19484 10968 19901 10996
rect 19484 10956 19490 10968
rect 19889 10965 19901 10968
rect 19935 10996 19947 10999
rect 20364 10996 20392 11036
rect 20990 11024 20996 11036
rect 21048 11024 21054 11076
rect 35728 11064 35756 11092
rect 37476 11064 37504 11095
rect 35728 11036 37504 11064
rect 40497 11067 40555 11073
rect 40497 11033 40509 11067
rect 40543 11064 40555 11067
rect 41414 11064 41420 11076
rect 40543 11036 41420 11064
rect 40543 11033 40555 11036
rect 40497 11027 40555 11033
rect 41414 11024 41420 11036
rect 41472 11024 41478 11076
rect 42150 11064 42156 11076
rect 42111 11036 42156 11064
rect 42150 11024 42156 11036
rect 42208 11024 42214 11076
rect 25682 10996 25688 11008
rect 19935 10968 20392 10996
rect 25643 10968 25688 10996
rect 19935 10965 19947 10968
rect 19889 10959 19947 10965
rect 25682 10956 25688 10968
rect 25740 10956 25746 11008
rect 33318 10996 33324 11008
rect 33279 10968 33324 10996
rect 33318 10956 33324 10968
rect 33376 10956 33382 11008
rect 33410 10956 33416 11008
rect 33468 10996 33474 11008
rect 33505 10999 33563 11005
rect 33505 10996 33517 10999
rect 33468 10968 33517 10996
rect 33468 10956 33474 10968
rect 33505 10965 33517 10968
rect 33551 10965 33563 10999
rect 35618 10996 35624 11008
rect 35579 10968 35624 10996
rect 33505 10959 33563 10965
rect 35618 10956 35624 10968
rect 35676 10956 35682 11008
rect 37550 10996 37556 11008
rect 37511 10968 37556 10996
rect 37550 10956 37556 10968
rect 37608 10956 37614 11008
rect 1104 10906 42872 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 42872 10906
rect 1104 10832 42872 10854
rect 18690 10752 18696 10804
rect 18748 10792 18754 10804
rect 18748 10764 20024 10792
rect 18748 10752 18754 10764
rect 18138 10724 18144 10736
rect 18099 10696 18144 10724
rect 18138 10684 18144 10696
rect 18196 10684 18202 10736
rect 19242 10684 19248 10736
rect 19300 10724 19306 10736
rect 19996 10724 20024 10764
rect 21082 10752 21088 10804
rect 21140 10792 21146 10804
rect 21269 10795 21327 10801
rect 21269 10792 21281 10795
rect 21140 10764 21281 10792
rect 21140 10752 21146 10764
rect 21269 10761 21281 10764
rect 21315 10761 21327 10795
rect 21269 10755 21327 10761
rect 23845 10795 23903 10801
rect 23845 10761 23857 10795
rect 23891 10761 23903 10795
rect 23845 10755 23903 10761
rect 25685 10795 25743 10801
rect 25685 10761 25697 10795
rect 25731 10792 25743 10795
rect 25774 10792 25780 10804
rect 25731 10764 25780 10792
rect 25731 10761 25743 10764
rect 25685 10755 25743 10761
rect 23860 10724 23888 10755
rect 25774 10752 25780 10764
rect 25832 10752 25838 10804
rect 28350 10792 28356 10804
rect 28311 10764 28356 10792
rect 28350 10752 28356 10764
rect 28408 10752 28414 10804
rect 32861 10795 32919 10801
rect 32861 10761 32873 10795
rect 32907 10792 32919 10795
rect 33318 10792 33324 10804
rect 32907 10764 33324 10792
rect 32907 10761 32919 10764
rect 32861 10755 32919 10761
rect 33318 10752 33324 10764
rect 33376 10752 33382 10804
rect 34977 10795 35035 10801
rect 34977 10761 34989 10795
rect 35023 10792 35035 10795
rect 35618 10792 35624 10804
rect 35023 10764 35624 10792
rect 35023 10761 35035 10764
rect 34977 10755 35035 10761
rect 35618 10752 35624 10764
rect 35676 10752 35682 10804
rect 41414 10792 41420 10804
rect 41375 10764 41420 10792
rect 41414 10752 41420 10764
rect 41472 10752 41478 10804
rect 24550 10727 24608 10733
rect 24550 10724 24562 10727
rect 19300 10696 19932 10724
rect 19996 10696 22094 10724
rect 23860 10696 24562 10724
rect 19300 10684 19306 10696
rect 1670 10656 1676 10668
rect 1631 10628 1676 10656
rect 1670 10616 1676 10628
rect 1728 10616 1734 10668
rect 14090 10616 14096 10668
rect 14148 10656 14154 10668
rect 14734 10656 14740 10668
rect 14148 10628 14740 10656
rect 14148 10616 14154 10628
rect 14734 10616 14740 10628
rect 14792 10616 14798 10668
rect 14826 10616 14832 10668
rect 14884 10656 14890 10668
rect 14993 10659 15051 10665
rect 14993 10656 15005 10659
rect 14884 10628 15005 10656
rect 14884 10616 14890 10628
rect 14993 10625 15005 10628
rect 15039 10625 15051 10659
rect 18506 10656 18512 10668
rect 18467 10628 18512 10656
rect 14993 10619 15051 10625
rect 18506 10616 18512 10628
rect 18564 10656 18570 10668
rect 19058 10656 19064 10668
rect 18564 10628 19064 10656
rect 18564 10616 18570 10628
rect 19058 10616 19064 10628
rect 19116 10656 19122 10668
rect 19337 10659 19395 10665
rect 19337 10656 19349 10659
rect 19116 10628 19349 10656
rect 19116 10616 19122 10628
rect 19337 10625 19349 10628
rect 19383 10625 19395 10659
rect 19337 10619 19395 10625
rect 19426 10616 19432 10668
rect 19484 10656 19490 10668
rect 19904 10665 19932 10696
rect 19889 10659 19947 10665
rect 19484 10628 19529 10656
rect 19484 10616 19490 10628
rect 19889 10625 19901 10659
rect 19935 10625 19947 10659
rect 19889 10619 19947 10625
rect 19978 10616 19984 10668
rect 20036 10656 20042 10668
rect 20145 10659 20203 10665
rect 20145 10656 20157 10659
rect 20036 10628 20157 10656
rect 20036 10616 20042 10628
rect 20145 10625 20157 10628
rect 20191 10625 20203 10659
rect 22066 10656 22094 10696
rect 24550 10693 24562 10696
rect 24596 10693 24608 10727
rect 24550 10687 24608 10693
rect 28813 10727 28871 10733
rect 28813 10693 28825 10727
rect 28859 10724 28871 10727
rect 30282 10724 30288 10736
rect 28859 10696 30288 10724
rect 28859 10693 28871 10696
rect 28813 10687 28871 10693
rect 30282 10684 30288 10696
rect 30340 10684 30346 10736
rect 30466 10684 30472 10736
rect 30524 10724 30530 10736
rect 30662 10727 30720 10733
rect 30662 10724 30674 10727
rect 30524 10696 30674 10724
rect 30524 10684 30530 10696
rect 30662 10693 30674 10696
rect 30708 10693 30720 10727
rect 30662 10687 30720 10693
rect 35434 10684 35440 10736
rect 35492 10724 35498 10736
rect 35492 10696 36308 10724
rect 35492 10684 35498 10696
rect 23017 10659 23075 10665
rect 23017 10656 23029 10659
rect 22066 10628 23029 10656
rect 20145 10619 20203 10625
rect 23017 10625 23029 10628
rect 23063 10625 23075 10659
rect 23017 10619 23075 10625
rect 23201 10659 23259 10665
rect 23201 10625 23213 10659
rect 23247 10656 23259 10659
rect 23661 10659 23719 10665
rect 23661 10656 23673 10659
rect 23247 10628 23673 10656
rect 23247 10625 23259 10628
rect 23201 10619 23259 10625
rect 23661 10625 23673 10628
rect 23707 10625 23719 10659
rect 23661 10619 23719 10625
rect 28721 10659 28779 10665
rect 28721 10625 28733 10659
rect 28767 10656 28779 10659
rect 29914 10656 29920 10668
rect 28767 10628 29920 10656
rect 28767 10625 28779 10628
rect 28721 10619 28779 10625
rect 29914 10616 29920 10628
rect 29972 10616 29978 10668
rect 30834 10616 30840 10668
rect 30892 10656 30898 10668
rect 30929 10659 30987 10665
rect 30929 10656 30941 10659
rect 30892 10628 30941 10656
rect 30892 10616 30898 10628
rect 30929 10625 30941 10628
rect 30975 10625 30987 10659
rect 30929 10619 30987 10625
rect 31573 10659 31631 10665
rect 31573 10625 31585 10659
rect 31619 10656 31631 10659
rect 32582 10656 32588 10668
rect 31619 10628 32588 10656
rect 31619 10625 31631 10628
rect 31573 10619 31631 10625
rect 32582 10616 32588 10628
rect 32640 10616 32646 10668
rect 32953 10659 33011 10665
rect 32953 10625 32965 10659
rect 32999 10656 33011 10659
rect 33318 10656 33324 10668
rect 32999 10628 33324 10656
rect 32999 10625 33011 10628
rect 32953 10619 33011 10625
rect 33318 10616 33324 10628
rect 33376 10616 33382 10668
rect 34885 10659 34943 10665
rect 34885 10625 34897 10659
rect 34931 10656 34943 10659
rect 35342 10656 35348 10668
rect 34931 10628 35348 10656
rect 34931 10625 34943 10628
rect 34885 10619 34943 10625
rect 35342 10616 35348 10628
rect 35400 10616 35406 10668
rect 35894 10616 35900 10668
rect 35952 10656 35958 10668
rect 35989 10659 36047 10665
rect 35989 10656 36001 10659
rect 35952 10628 36001 10656
rect 35952 10616 35958 10628
rect 35989 10625 36001 10628
rect 36035 10625 36047 10659
rect 35989 10619 36047 10625
rect 36081 10659 36139 10665
rect 36081 10625 36093 10659
rect 36127 10625 36139 10659
rect 36081 10619 36139 10625
rect 36173 10659 36231 10665
rect 36173 10625 36185 10659
rect 36219 10656 36231 10659
rect 36280 10656 36308 10696
rect 36219 10628 36308 10656
rect 36357 10659 36415 10665
rect 36219 10625 36231 10628
rect 36173 10619 36231 10625
rect 36357 10625 36369 10659
rect 36403 10656 36415 10659
rect 37182 10656 37188 10668
rect 36403 10628 37188 10656
rect 36403 10625 36415 10628
rect 36357 10619 36415 10625
rect 1857 10591 1915 10597
rect 1857 10557 1869 10591
rect 1903 10588 1915 10591
rect 2038 10588 2044 10600
rect 1903 10560 2044 10588
rect 1903 10557 1915 10560
rect 1857 10551 1915 10557
rect 2038 10548 2044 10560
rect 2096 10548 2102 10600
rect 2774 10548 2780 10600
rect 2832 10588 2838 10600
rect 16669 10591 16727 10597
rect 2832 10560 2877 10588
rect 2832 10548 2838 10560
rect 16669 10557 16681 10591
rect 16715 10557 16727 10591
rect 16942 10588 16948 10600
rect 16903 10560 16948 10588
rect 16669 10551 16727 10557
rect 16117 10523 16175 10529
rect 16117 10489 16129 10523
rect 16163 10520 16175 10523
rect 16482 10520 16488 10532
rect 16163 10492 16488 10520
rect 16163 10489 16175 10492
rect 16117 10483 16175 10489
rect 16482 10480 16488 10492
rect 16540 10520 16546 10532
rect 16684 10520 16712 10551
rect 16942 10548 16948 10560
rect 17000 10548 17006 10600
rect 19150 10588 19156 10600
rect 19111 10560 19156 10588
rect 19150 10548 19156 10560
rect 19208 10548 19214 10600
rect 22830 10588 22836 10600
rect 22791 10560 22836 10588
rect 22830 10548 22836 10560
rect 22888 10548 22894 10600
rect 24305 10591 24363 10597
rect 24305 10557 24317 10591
rect 24351 10557 24363 10591
rect 24305 10551 24363 10557
rect 18230 10520 18236 10532
rect 16540 10492 16712 10520
rect 18143 10492 18236 10520
rect 16540 10480 16546 10492
rect 17957 10455 18015 10461
rect 17957 10421 17969 10455
rect 18003 10452 18015 10455
rect 18046 10452 18052 10464
rect 18003 10424 18052 10452
rect 18003 10421 18015 10424
rect 17957 10415 18015 10421
rect 18046 10412 18052 10424
rect 18104 10412 18110 10464
rect 18156 10461 18184 10492
rect 18230 10480 18236 10492
rect 18288 10520 18294 10532
rect 19168 10520 19196 10548
rect 18288 10492 19196 10520
rect 18288 10480 18294 10492
rect 18141 10455 18199 10461
rect 18141 10421 18153 10455
rect 18187 10421 18199 10455
rect 19242 10452 19248 10464
rect 19203 10424 19248 10452
rect 18141 10415 18199 10421
rect 19242 10412 19248 10424
rect 19300 10412 19306 10464
rect 24320 10452 24348 10551
rect 28902 10548 28908 10600
rect 28960 10588 28966 10600
rect 33042 10588 33048 10600
rect 28960 10560 29005 10588
rect 32955 10560 33048 10588
rect 28960 10548 28966 10560
rect 33042 10548 33048 10560
rect 33100 10588 33106 10600
rect 35069 10591 35127 10597
rect 35069 10588 35081 10591
rect 33100 10560 35081 10588
rect 33100 10548 33106 10560
rect 35069 10557 35081 10560
rect 35115 10557 35127 10591
rect 36096 10588 36124 10619
rect 37182 10616 37188 10628
rect 37240 10616 37246 10668
rect 41509 10659 41567 10665
rect 41509 10625 41521 10659
rect 41555 10656 41567 10659
rect 42242 10656 42248 10668
rect 41555 10628 42248 10656
rect 41555 10625 41567 10628
rect 41509 10619 41567 10625
rect 42242 10616 42248 10628
rect 42300 10616 42306 10668
rect 36262 10588 36268 10600
rect 36096 10560 36268 10588
rect 35069 10551 35127 10557
rect 36262 10548 36268 10560
rect 36320 10548 36326 10600
rect 25314 10452 25320 10464
rect 24320 10424 25320 10452
rect 25314 10412 25320 10424
rect 25372 10412 25378 10464
rect 29549 10455 29607 10461
rect 29549 10421 29561 10455
rect 29595 10452 29607 10455
rect 30558 10452 30564 10464
rect 29595 10424 30564 10452
rect 29595 10421 29607 10424
rect 29549 10415 29607 10421
rect 30558 10412 30564 10424
rect 30616 10412 30622 10464
rect 31110 10412 31116 10464
rect 31168 10452 31174 10464
rect 31389 10455 31447 10461
rect 31389 10452 31401 10455
rect 31168 10424 31401 10452
rect 31168 10412 31174 10424
rect 31389 10421 31401 10424
rect 31435 10421 31447 10455
rect 31389 10415 31447 10421
rect 32306 10412 32312 10464
rect 32364 10452 32370 10464
rect 32493 10455 32551 10461
rect 32493 10452 32505 10455
rect 32364 10424 32505 10452
rect 32364 10412 32370 10424
rect 32493 10421 32505 10424
rect 32539 10421 32551 10455
rect 32493 10415 32551 10421
rect 33042 10412 33048 10464
rect 33100 10452 33106 10464
rect 34517 10455 34575 10461
rect 34517 10452 34529 10455
rect 33100 10424 34529 10452
rect 33100 10412 33106 10424
rect 34517 10421 34529 10424
rect 34563 10421 34575 10455
rect 35710 10452 35716 10464
rect 35671 10424 35716 10452
rect 34517 10415 34575 10421
rect 35710 10412 35716 10424
rect 35768 10412 35774 10464
rect 40310 10412 40316 10464
rect 40368 10452 40374 10464
rect 40681 10455 40739 10461
rect 40681 10452 40693 10455
rect 40368 10424 40693 10452
rect 40368 10412 40374 10424
rect 40681 10421 40693 10424
rect 40727 10421 40739 10455
rect 40681 10415 40739 10421
rect 1104 10362 42872 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 42872 10362
rect 1104 10288 42872 10310
rect 2038 10248 2044 10260
rect 1999 10220 2044 10248
rect 2038 10208 2044 10220
rect 2096 10208 2102 10260
rect 14826 10248 14832 10260
rect 14787 10220 14832 10248
rect 14826 10208 14832 10220
rect 14884 10208 14890 10260
rect 15841 10251 15899 10257
rect 15841 10217 15853 10251
rect 15887 10248 15899 10251
rect 15930 10248 15936 10260
rect 15887 10220 15936 10248
rect 15887 10217 15899 10220
rect 15841 10211 15899 10217
rect 15930 10208 15936 10220
rect 15988 10208 15994 10260
rect 16482 10248 16488 10260
rect 16443 10220 16488 10248
rect 16482 10208 16488 10220
rect 16540 10208 16546 10260
rect 16669 10251 16727 10257
rect 16669 10217 16681 10251
rect 16715 10248 16727 10251
rect 17494 10248 17500 10260
rect 16715 10220 17500 10248
rect 16715 10217 16727 10220
rect 16669 10211 16727 10217
rect 17494 10208 17500 10220
rect 17552 10208 17558 10260
rect 18230 10208 18236 10260
rect 18288 10248 18294 10260
rect 18690 10248 18696 10260
rect 18288 10220 18696 10248
rect 18288 10208 18294 10220
rect 18690 10208 18696 10220
rect 18748 10208 18754 10260
rect 19613 10251 19671 10257
rect 19613 10217 19625 10251
rect 19659 10248 19671 10251
rect 19978 10248 19984 10260
rect 19659 10220 19984 10248
rect 19659 10217 19671 10220
rect 19613 10211 19671 10217
rect 19978 10208 19984 10220
rect 20036 10208 20042 10260
rect 22554 10248 22560 10260
rect 22515 10220 22560 10248
rect 22554 10208 22560 10220
rect 22612 10208 22618 10260
rect 23201 10251 23259 10257
rect 23201 10217 23213 10251
rect 23247 10248 23259 10251
rect 23474 10248 23480 10260
rect 23247 10220 23480 10248
rect 23247 10217 23259 10220
rect 23201 10211 23259 10217
rect 23474 10208 23480 10220
rect 23532 10208 23538 10260
rect 32582 10248 32588 10260
rect 32543 10220 32588 10248
rect 32582 10208 32588 10220
rect 32640 10208 32646 10260
rect 35161 10251 35219 10257
rect 35161 10217 35173 10251
rect 35207 10217 35219 10251
rect 35161 10211 35219 10217
rect 35176 10180 35204 10211
rect 35342 10208 35348 10260
rect 35400 10248 35406 10260
rect 35713 10251 35771 10257
rect 35713 10248 35725 10251
rect 35400 10220 35725 10248
rect 35400 10208 35406 10220
rect 35713 10217 35725 10220
rect 35759 10217 35771 10251
rect 35713 10211 35771 10217
rect 36170 10180 36176 10192
rect 35176 10152 36176 10180
rect 36170 10140 36176 10152
rect 36228 10140 36234 10192
rect 14734 10072 14740 10124
rect 14792 10112 14798 10124
rect 16850 10112 16856 10124
rect 14792 10084 16856 10112
rect 14792 10072 14798 10084
rect 16850 10072 16856 10084
rect 16908 10112 16914 10124
rect 17310 10112 17316 10124
rect 16908 10084 17316 10112
rect 16908 10072 16914 10084
rect 17310 10072 17316 10084
rect 17368 10072 17374 10124
rect 19058 10072 19064 10124
rect 19116 10112 19122 10124
rect 33042 10112 33048 10124
rect 19116 10084 19932 10112
rect 33003 10084 33048 10112
rect 19116 10072 19122 10084
rect 2130 10044 2136 10056
rect 2091 10016 2136 10044
rect 2130 10004 2136 10016
rect 2188 10004 2194 10056
rect 2777 10047 2835 10053
rect 2777 10013 2789 10047
rect 2823 10044 2835 10047
rect 3234 10044 3240 10056
rect 2823 10016 3240 10044
rect 2823 10013 2835 10016
rect 2777 10007 2835 10013
rect 3234 10004 3240 10016
rect 3292 10004 3298 10056
rect 15105 10047 15163 10053
rect 15105 10013 15117 10047
rect 15151 10044 15163 10047
rect 15378 10044 15384 10056
rect 15151 10016 15384 10044
rect 15151 10013 15163 10016
rect 15105 10007 15163 10013
rect 15378 10004 15384 10016
rect 15436 10004 15442 10056
rect 15565 10047 15623 10053
rect 15565 10013 15577 10047
rect 15611 10044 15623 10047
rect 15654 10044 15660 10056
rect 15611 10016 15660 10044
rect 15611 10013 15623 10016
rect 15565 10007 15623 10013
rect 14829 9979 14887 9985
rect 14829 9945 14841 9979
rect 14875 9976 14887 9979
rect 15470 9976 15476 9988
rect 14875 9948 15476 9976
rect 14875 9945 14887 9948
rect 14829 9939 14887 9945
rect 15470 9936 15476 9948
rect 15528 9936 15534 9988
rect 15013 9911 15071 9917
rect 15013 9877 15025 9911
rect 15059 9908 15071 9911
rect 15580 9908 15608 10007
rect 15654 10004 15660 10016
rect 15712 10004 15718 10056
rect 15841 10047 15899 10053
rect 15841 10013 15853 10047
rect 15887 10013 15899 10047
rect 15841 10007 15899 10013
rect 15856 9976 15884 10007
rect 19242 10004 19248 10056
rect 19300 10044 19306 10056
rect 19904 10053 19932 10084
rect 33042 10072 33048 10084
rect 33100 10072 33106 10124
rect 33137 10115 33195 10121
rect 33137 10081 33149 10115
rect 33183 10112 33195 10115
rect 33410 10112 33416 10124
rect 33183 10084 33416 10112
rect 33183 10081 33195 10084
rect 33137 10075 33195 10081
rect 33410 10072 33416 10084
rect 33468 10072 33474 10124
rect 34977 10115 35035 10121
rect 34977 10081 34989 10115
rect 35023 10112 35035 10115
rect 36814 10112 36820 10124
rect 35023 10084 36820 10112
rect 35023 10081 35035 10084
rect 34977 10075 35035 10081
rect 19613 10047 19671 10053
rect 19613 10044 19625 10047
rect 19300 10016 19625 10044
rect 19300 10004 19306 10016
rect 19613 10013 19625 10016
rect 19659 10013 19671 10047
rect 19613 10007 19671 10013
rect 19889 10047 19947 10053
rect 19889 10013 19901 10047
rect 19935 10013 19947 10047
rect 19889 10007 19947 10013
rect 21913 10047 21971 10053
rect 21913 10013 21925 10047
rect 21959 10044 21971 10047
rect 22186 10044 22192 10056
rect 21959 10016 22192 10044
rect 21959 10013 21971 10016
rect 21913 10007 21971 10013
rect 22186 10004 22192 10016
rect 22244 10004 22250 10056
rect 22370 10044 22376 10056
rect 22331 10016 22376 10044
rect 22370 10004 22376 10016
rect 22428 10004 22434 10056
rect 22554 10004 22560 10056
rect 22612 10044 22618 10056
rect 23017 10047 23075 10053
rect 23017 10044 23029 10047
rect 22612 10016 23029 10044
rect 22612 10004 22618 10016
rect 23017 10013 23029 10016
rect 23063 10013 23075 10047
rect 23017 10007 23075 10013
rect 25314 10004 25320 10056
rect 25372 10044 25378 10056
rect 25409 10047 25467 10053
rect 25409 10044 25421 10047
rect 25372 10016 25421 10044
rect 25372 10004 25378 10016
rect 25409 10013 25421 10016
rect 25455 10044 25467 10047
rect 27338 10044 27344 10056
rect 25455 10016 27344 10044
rect 25455 10013 25467 10016
rect 25409 10007 25467 10013
rect 27338 10004 27344 10016
rect 27396 10004 27402 10056
rect 30834 10004 30840 10056
rect 30892 10044 30898 10056
rect 31389 10047 31447 10053
rect 31389 10044 31401 10047
rect 30892 10016 31401 10044
rect 30892 10004 30898 10016
rect 31389 10013 31401 10016
rect 31435 10044 31447 10047
rect 31478 10044 31484 10056
rect 31435 10016 31484 10044
rect 31435 10013 31447 10016
rect 31389 10007 31447 10013
rect 31478 10004 31484 10016
rect 31536 10004 31542 10056
rect 32953 10047 33011 10053
rect 32953 10013 32965 10047
rect 32999 10044 33011 10047
rect 33226 10044 33232 10056
rect 32999 10016 33232 10044
rect 32999 10013 33011 10016
rect 32953 10007 33011 10013
rect 33226 10004 33232 10016
rect 33284 10004 33290 10056
rect 35253 10047 35311 10053
rect 35253 10013 35265 10047
rect 35299 10044 35311 10047
rect 35434 10044 35440 10056
rect 35299 10016 35440 10044
rect 35299 10013 35311 10016
rect 35253 10007 35311 10013
rect 35434 10004 35440 10016
rect 35492 10004 35498 10056
rect 35710 10044 35716 10056
rect 35671 10016 35716 10044
rect 35710 10004 35716 10016
rect 35768 10004 35774 10056
rect 35912 10053 35940 10084
rect 36814 10072 36820 10084
rect 36872 10072 36878 10124
rect 40310 10112 40316 10124
rect 40271 10084 40316 10112
rect 40310 10072 40316 10084
rect 40368 10072 40374 10124
rect 42150 10112 42156 10124
rect 42111 10084 42156 10112
rect 42150 10072 42156 10084
rect 42208 10072 42214 10124
rect 35897 10047 35955 10053
rect 35897 10013 35909 10047
rect 35943 10013 35955 10047
rect 35897 10007 35955 10013
rect 35989 10047 36047 10053
rect 35989 10013 36001 10047
rect 36035 10044 36047 10047
rect 37550 10044 37556 10056
rect 36035 10016 37556 10044
rect 36035 10013 36047 10016
rect 35989 10007 36047 10013
rect 37550 10004 37556 10016
rect 37608 10004 37614 10056
rect 16301 9979 16359 9985
rect 16301 9976 16313 9979
rect 15856 9948 16313 9976
rect 16301 9945 16313 9948
rect 16347 9976 16359 9979
rect 17580 9979 17638 9985
rect 16347 9948 17540 9976
rect 16347 9945 16359 9948
rect 16301 9939 16359 9945
rect 15059 9880 15608 9908
rect 15657 9911 15715 9917
rect 15059 9877 15071 9880
rect 15013 9871 15071 9877
rect 15657 9877 15669 9911
rect 15703 9908 15715 9911
rect 16114 9908 16120 9920
rect 15703 9880 16120 9908
rect 15703 9877 15715 9880
rect 15657 9871 15715 9877
rect 16114 9868 16120 9880
rect 16172 9868 16178 9920
rect 16482 9868 16488 9920
rect 16540 9917 16546 9920
rect 16540 9911 16559 9917
rect 16547 9877 16559 9911
rect 17512 9908 17540 9948
rect 17580 9945 17592 9979
rect 17626 9976 17638 9979
rect 17954 9976 17960 9988
rect 17626 9948 17960 9976
rect 17626 9945 17638 9948
rect 17580 9939 17638 9945
rect 17954 9936 17960 9948
rect 18012 9936 18018 9988
rect 19426 9936 19432 9988
rect 19484 9976 19490 9988
rect 25682 9985 25688 9988
rect 19797 9979 19855 9985
rect 19797 9976 19809 9979
rect 19484 9948 19809 9976
rect 19484 9936 19490 9948
rect 19797 9945 19809 9948
rect 19843 9945 19855 9979
rect 25676 9976 25688 9985
rect 25643 9948 25688 9976
rect 19797 9939 19855 9945
rect 25676 9939 25688 9948
rect 25682 9936 25688 9939
rect 25740 9936 25746 9988
rect 27614 9985 27620 9988
rect 27608 9939 27620 9985
rect 27672 9976 27678 9988
rect 27672 9948 27708 9976
rect 27614 9936 27620 9939
rect 27672 9936 27678 9948
rect 31110 9936 31116 9988
rect 31168 9985 31174 9988
rect 31168 9976 31180 9985
rect 40497 9979 40555 9985
rect 31168 9948 31213 9976
rect 31168 9939 31180 9948
rect 40497 9945 40509 9979
rect 40543 9976 40555 9979
rect 41414 9976 41420 9988
rect 40543 9948 41420 9976
rect 40543 9945 40555 9948
rect 40497 9939 40555 9945
rect 31168 9936 31174 9939
rect 41414 9936 41420 9948
rect 41472 9936 41478 9988
rect 18230 9908 18236 9920
rect 17512 9880 18236 9908
rect 16540 9871 16559 9877
rect 16540 9868 16546 9871
rect 18230 9868 18236 9880
rect 18288 9868 18294 9920
rect 21726 9908 21732 9920
rect 21687 9880 21732 9908
rect 21726 9868 21732 9880
rect 21784 9868 21790 9920
rect 28721 9911 28779 9917
rect 28721 9877 28733 9911
rect 28767 9908 28779 9911
rect 29546 9908 29552 9920
rect 28767 9880 29552 9908
rect 28767 9877 28779 9880
rect 28721 9871 28779 9877
rect 29546 9868 29552 9880
rect 29604 9868 29610 9920
rect 30009 9911 30067 9917
rect 30009 9877 30021 9911
rect 30055 9908 30067 9911
rect 30374 9908 30380 9920
rect 30055 9880 30380 9908
rect 30055 9877 30067 9880
rect 30009 9871 30067 9877
rect 30374 9868 30380 9880
rect 30432 9868 30438 9920
rect 34698 9908 34704 9920
rect 34659 9880 34704 9908
rect 34698 9868 34704 9880
rect 34756 9868 34762 9920
rect 1104 9818 42872 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 42872 9818
rect 1104 9744 42872 9766
rect 18138 9664 18144 9716
rect 18196 9704 18202 9716
rect 18601 9707 18659 9713
rect 18601 9704 18613 9707
rect 18196 9676 18613 9704
rect 18196 9664 18202 9676
rect 18601 9673 18613 9676
rect 18647 9673 18659 9707
rect 18601 9667 18659 9673
rect 27893 9707 27951 9713
rect 27893 9673 27905 9707
rect 27939 9704 27951 9707
rect 28902 9704 28908 9716
rect 27939 9676 28908 9704
rect 27939 9673 27951 9676
rect 27893 9667 27951 9673
rect 28902 9664 28908 9676
rect 28960 9664 28966 9716
rect 29914 9664 29920 9716
rect 29972 9704 29978 9716
rect 30009 9707 30067 9713
rect 30009 9704 30021 9707
rect 29972 9676 30021 9704
rect 29972 9664 29978 9676
rect 30009 9673 30021 9676
rect 30055 9673 30067 9707
rect 30009 9667 30067 9673
rect 30469 9707 30527 9713
rect 30469 9673 30481 9707
rect 30515 9704 30527 9707
rect 30558 9704 30564 9716
rect 30515 9676 30564 9704
rect 30515 9673 30527 9676
rect 30469 9667 30527 9673
rect 30558 9664 30564 9676
rect 30616 9664 30622 9716
rect 15470 9596 15476 9648
rect 15528 9636 15534 9648
rect 15565 9639 15623 9645
rect 15565 9636 15577 9639
rect 15528 9608 15577 9636
rect 15528 9596 15534 9608
rect 15565 9605 15577 9608
rect 15611 9605 15623 9639
rect 15565 9599 15623 9605
rect 15654 9596 15660 9648
rect 15712 9636 15718 9648
rect 16942 9636 16948 9648
rect 15712 9608 16948 9636
rect 15712 9596 15718 9608
rect 2317 9571 2375 9577
rect 2317 9537 2329 9571
rect 2363 9568 2375 9571
rect 2961 9571 3019 9577
rect 2961 9568 2973 9571
rect 2363 9540 2973 9568
rect 2363 9537 2375 9540
rect 2317 9531 2375 9537
rect 2961 9537 2973 9540
rect 3007 9568 3019 9571
rect 4706 9568 4712 9580
rect 3007 9540 4712 9568
rect 3007 9537 3019 9540
rect 2961 9531 3019 9537
rect 4706 9528 4712 9540
rect 4764 9528 4770 9580
rect 15378 9528 15384 9580
rect 15436 9568 15442 9580
rect 15856 9577 15884 9608
rect 16942 9596 16948 9608
rect 17000 9636 17006 9648
rect 17000 9608 18552 9636
rect 17000 9596 17006 9608
rect 15749 9571 15807 9577
rect 15749 9568 15761 9571
rect 15436 9540 15761 9568
rect 15436 9528 15442 9540
rect 15749 9537 15761 9540
rect 15795 9537 15807 9571
rect 15749 9531 15807 9537
rect 15841 9571 15899 9577
rect 15841 9537 15853 9571
rect 15887 9537 15899 9571
rect 15841 9531 15899 9537
rect 16298 9528 16304 9580
rect 16356 9568 16362 9580
rect 18417 9571 18475 9577
rect 18417 9568 18429 9571
rect 16356 9540 18429 9568
rect 16356 9528 16362 9540
rect 18417 9537 18429 9540
rect 18463 9537 18475 9571
rect 18417 9531 18475 9537
rect 18524 9512 18552 9608
rect 18782 9596 18788 9648
rect 18840 9636 18846 9648
rect 25774 9636 25780 9648
rect 18840 9608 22048 9636
rect 18840 9596 18846 9608
rect 21726 9528 21732 9580
rect 21784 9568 21790 9580
rect 22020 9577 22048 9608
rect 25424 9608 25780 9636
rect 21821 9571 21879 9577
rect 21821 9568 21833 9571
rect 21784 9540 21833 9568
rect 21784 9528 21790 9540
rect 21821 9537 21833 9540
rect 21867 9537 21879 9571
rect 21821 9531 21879 9537
rect 22005 9571 22063 9577
rect 22005 9537 22017 9571
rect 22051 9537 22063 9571
rect 22005 9531 22063 9537
rect 22186 9528 22192 9580
rect 22244 9568 22250 9580
rect 23566 9577 23572 9580
rect 22649 9571 22707 9577
rect 22649 9568 22661 9571
rect 22244 9540 22661 9568
rect 22244 9528 22250 9540
rect 22649 9537 22661 9540
rect 22695 9537 22707 9571
rect 22649 9531 22707 9537
rect 23560 9531 23572 9577
rect 23624 9568 23630 9580
rect 25424 9577 25452 9608
rect 25774 9596 25780 9608
rect 25832 9636 25838 9648
rect 26237 9639 26295 9645
rect 26237 9636 26249 9639
rect 25832 9608 26249 9636
rect 25832 9596 25838 9608
rect 26237 9605 26249 9608
rect 26283 9605 26295 9639
rect 27154 9636 27160 9648
rect 26237 9599 26295 9605
rect 26344 9608 27160 9636
rect 25317 9571 25375 9577
rect 25317 9568 25329 9571
rect 23624 9540 23660 9568
rect 24688 9540 25329 9568
rect 23566 9528 23572 9531
rect 23624 9528 23630 9540
rect 15565 9503 15623 9509
rect 15565 9469 15577 9503
rect 15611 9500 15623 9503
rect 15930 9500 15936 9512
rect 15611 9472 15936 9500
rect 15611 9469 15623 9472
rect 15565 9463 15623 9469
rect 15930 9460 15936 9472
rect 15988 9500 15994 9512
rect 17126 9500 17132 9512
rect 15988 9472 17132 9500
rect 15988 9460 15994 9472
rect 17126 9460 17132 9472
rect 17184 9460 17190 9512
rect 18138 9500 18144 9512
rect 18099 9472 18144 9500
rect 18138 9460 18144 9472
rect 18196 9460 18202 9512
rect 18233 9503 18291 9509
rect 18233 9469 18245 9503
rect 18279 9469 18291 9503
rect 18233 9463 18291 9469
rect 18325 9503 18383 9509
rect 18325 9469 18337 9503
rect 18371 9500 18383 9503
rect 18506 9500 18512 9512
rect 18371 9472 18512 9500
rect 18371 9469 18383 9472
rect 18325 9463 18383 9469
rect 16114 9392 16120 9444
rect 16172 9432 16178 9444
rect 18248 9432 18276 9463
rect 18506 9460 18512 9472
rect 18564 9460 18570 9512
rect 18690 9460 18696 9512
rect 18748 9500 18754 9512
rect 18748 9472 22094 9500
rect 18748 9460 18754 9472
rect 18782 9432 18788 9444
rect 16172 9404 18788 9432
rect 16172 9392 16178 9404
rect 18782 9392 18788 9404
rect 18840 9392 18846 9444
rect 1673 9367 1731 9373
rect 1673 9333 1685 9367
rect 1719 9364 1731 9367
rect 1762 9364 1768 9376
rect 1719 9336 1768 9364
rect 1719 9333 1731 9336
rect 1673 9327 1731 9333
rect 1762 9324 1768 9336
rect 1820 9324 1826 9376
rect 2222 9364 2228 9376
rect 2183 9336 2228 9364
rect 2222 9324 2228 9336
rect 2280 9324 2286 9376
rect 2866 9364 2872 9376
rect 2827 9336 2872 9364
rect 2866 9324 2872 9336
rect 2924 9324 2930 9376
rect 22066 9364 22094 9472
rect 22462 9460 22468 9512
rect 22520 9500 22526 9512
rect 23014 9500 23020 9512
rect 22520 9472 23020 9500
rect 22520 9460 22526 9472
rect 23014 9460 23020 9472
rect 23072 9500 23078 9512
rect 23293 9503 23351 9509
rect 23293 9500 23305 9503
rect 23072 9472 23305 9500
rect 23072 9460 23078 9472
rect 23293 9469 23305 9472
rect 23339 9469 23351 9503
rect 23293 9463 23351 9469
rect 22189 9435 22247 9441
rect 22189 9401 22201 9435
rect 22235 9432 22247 9435
rect 22922 9432 22928 9444
rect 22235 9404 22928 9432
rect 22235 9401 22247 9404
rect 22189 9395 22247 9401
rect 22922 9392 22928 9404
rect 22980 9392 22986 9444
rect 24688 9441 24716 9540
rect 25317 9537 25329 9540
rect 25363 9537 25375 9571
rect 25317 9531 25375 9537
rect 25409 9571 25467 9577
rect 25409 9537 25421 9571
rect 25455 9537 25467 9571
rect 25409 9531 25467 9537
rect 25498 9528 25504 9580
rect 25556 9568 25562 9580
rect 25593 9571 25651 9577
rect 25593 9568 25605 9571
rect 25556 9540 25605 9568
rect 25556 9528 25562 9540
rect 25593 9537 25605 9540
rect 25639 9537 25651 9571
rect 25593 9531 25651 9537
rect 26053 9571 26111 9577
rect 26053 9537 26065 9571
rect 26099 9568 26111 9571
rect 26344 9568 26372 9608
rect 27154 9596 27160 9608
rect 27212 9596 27218 9648
rect 30834 9636 30840 9648
rect 29288 9608 30840 9636
rect 26099 9540 26372 9568
rect 26421 9571 26479 9577
rect 26099 9537 26111 9540
rect 26053 9531 26111 9537
rect 26252 9512 26280 9540
rect 26421 9537 26433 9571
rect 26467 9568 26479 9571
rect 26973 9571 27031 9577
rect 26973 9568 26985 9571
rect 26467 9540 26985 9568
rect 26467 9537 26479 9540
rect 26421 9531 26479 9537
rect 26973 9537 26985 9540
rect 27019 9537 27031 9571
rect 26973 9531 27031 9537
rect 29017 9571 29075 9577
rect 29017 9537 29029 9571
rect 29063 9568 29075 9571
rect 29178 9568 29184 9580
rect 29063 9540 29184 9568
rect 29063 9537 29075 9540
rect 29017 9531 29075 9537
rect 29178 9528 29184 9540
rect 29236 9528 29242 9580
rect 29288 9577 29316 9608
rect 30834 9596 30840 9608
rect 30892 9596 30898 9648
rect 33318 9636 33324 9648
rect 33279 9608 33324 9636
rect 33318 9596 33324 9608
rect 33376 9596 33382 9648
rect 33965 9639 34023 9645
rect 33965 9605 33977 9639
rect 34011 9636 34023 9639
rect 34698 9636 34704 9648
rect 34011 9608 34704 9636
rect 34011 9605 34023 9608
rect 33965 9599 34023 9605
rect 34698 9596 34704 9608
rect 34756 9596 34762 9648
rect 41414 9636 41420 9648
rect 41375 9608 41420 9636
rect 41414 9596 41420 9608
rect 41472 9596 41478 9648
rect 29273 9571 29331 9577
rect 29273 9537 29285 9571
rect 29319 9537 29331 9571
rect 30374 9568 30380 9580
rect 30335 9540 30380 9568
rect 29273 9531 29331 9537
rect 30374 9528 30380 9540
rect 30432 9528 30438 9580
rect 32306 9568 32312 9580
rect 32267 9540 32312 9568
rect 32306 9528 32312 9540
rect 32364 9528 32370 9580
rect 33505 9571 33563 9577
rect 33505 9537 33517 9571
rect 33551 9568 33563 9571
rect 34330 9568 34336 9580
rect 33551 9540 34336 9568
rect 33551 9537 33563 9540
rect 33505 9531 33563 9537
rect 34330 9528 34336 9540
rect 34388 9528 34394 9580
rect 41138 9528 41144 9580
rect 41196 9568 41202 9580
rect 41325 9571 41383 9577
rect 41325 9568 41337 9571
rect 41196 9540 41337 9568
rect 41196 9528 41202 9540
rect 41325 9537 41337 9540
rect 41371 9537 41383 9571
rect 41325 9531 41383 9537
rect 26234 9460 26240 9512
rect 26292 9460 26298 9512
rect 30558 9460 30564 9512
rect 30616 9500 30622 9512
rect 30616 9472 30661 9500
rect 30616 9460 30622 9472
rect 33410 9460 33416 9512
rect 33468 9500 33474 9512
rect 33597 9503 33655 9509
rect 33597 9500 33609 9503
rect 33468 9472 33609 9500
rect 33468 9460 33474 9472
rect 33597 9469 33609 9472
rect 33643 9469 33655 9503
rect 33597 9463 33655 9469
rect 24673 9435 24731 9441
rect 24673 9401 24685 9435
rect 24719 9401 24731 9435
rect 25130 9432 25136 9444
rect 25091 9404 25136 9432
rect 24673 9395 24731 9401
rect 25130 9392 25136 9404
rect 25188 9392 25194 9444
rect 27157 9435 27215 9441
rect 27157 9401 27169 9435
rect 27203 9432 27215 9435
rect 27614 9432 27620 9444
rect 27203 9404 27620 9432
rect 27203 9401 27215 9404
rect 27157 9395 27215 9401
rect 27614 9392 27620 9404
rect 27672 9392 27678 9444
rect 22646 9364 22652 9376
rect 22066 9336 22652 9364
rect 22646 9324 22652 9336
rect 22704 9324 22710 9376
rect 22830 9364 22836 9376
rect 22791 9336 22836 9364
rect 22830 9324 22836 9336
rect 22888 9324 22894 9376
rect 25222 9324 25228 9376
rect 25280 9364 25286 9376
rect 25317 9367 25375 9373
rect 25317 9364 25329 9367
rect 25280 9336 25329 9364
rect 25280 9324 25286 9336
rect 25317 9333 25329 9336
rect 25363 9333 25375 9367
rect 32122 9364 32128 9376
rect 32083 9336 32128 9364
rect 25317 9327 25375 9333
rect 32122 9324 32128 9336
rect 32180 9324 32186 9376
rect 1104 9274 42872 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 42872 9274
rect 1104 9200 42872 9222
rect 17954 9160 17960 9172
rect 17915 9132 17960 9160
rect 17954 9120 17960 9132
rect 18012 9120 18018 9172
rect 19889 9163 19947 9169
rect 19889 9160 19901 9163
rect 18064 9132 19901 9160
rect 17862 9052 17868 9104
rect 17920 9092 17926 9104
rect 18064 9092 18092 9132
rect 19889 9129 19901 9132
rect 19935 9160 19947 9163
rect 21542 9160 21548 9172
rect 19935 9132 21548 9160
rect 19935 9129 19947 9132
rect 19889 9123 19947 9129
rect 21542 9120 21548 9132
rect 21600 9120 21606 9172
rect 21637 9163 21695 9169
rect 21637 9129 21649 9163
rect 21683 9160 21695 9163
rect 22370 9160 22376 9172
rect 21683 9132 22376 9160
rect 21683 9129 21695 9132
rect 21637 9123 21695 9129
rect 22370 9120 22376 9132
rect 22428 9120 22434 9172
rect 22465 9163 22523 9169
rect 22465 9129 22477 9163
rect 22511 9160 22523 9163
rect 22554 9160 22560 9172
rect 22511 9132 22560 9160
rect 22511 9129 22523 9132
rect 22465 9123 22523 9129
rect 22554 9120 22560 9132
rect 22612 9120 22618 9172
rect 29178 9120 29184 9172
rect 29236 9160 29242 9172
rect 30193 9163 30251 9169
rect 30193 9160 30205 9163
rect 29236 9132 30205 9160
rect 29236 9120 29242 9132
rect 30193 9129 30205 9132
rect 30239 9129 30251 9163
rect 30193 9123 30251 9129
rect 17920 9064 18092 9092
rect 17920 9052 17926 9064
rect 2222 8984 2228 9036
rect 2280 9024 2286 9036
rect 3053 9027 3111 9033
rect 3053 9024 3065 9027
rect 2280 8996 3065 9024
rect 2280 8984 2286 8996
rect 3053 8993 3065 8996
rect 3099 8993 3111 9027
rect 3234 9024 3240 9036
rect 3195 8996 3240 9024
rect 3053 8987 3111 8993
rect 3234 8984 3240 8996
rect 3292 8984 3298 9036
rect 16482 9024 16488 9036
rect 15488 8996 16488 9024
rect 1394 8956 1400 8968
rect 1355 8928 1400 8956
rect 1394 8916 1400 8928
rect 1452 8916 1458 8968
rect 15378 8916 15384 8968
rect 15436 8956 15442 8968
rect 15488 8965 15516 8996
rect 16482 8984 16488 8996
rect 16540 8984 16546 9036
rect 21269 9027 21327 9033
rect 21269 8993 21281 9027
rect 21315 9024 21327 9027
rect 21726 9024 21732 9036
rect 21315 8996 21732 9024
rect 21315 8993 21327 8996
rect 21269 8987 21327 8993
rect 21726 8984 21732 8996
rect 21784 9024 21790 9036
rect 22097 9027 22155 9033
rect 22097 9024 22109 9027
rect 21784 8996 22109 9024
rect 21784 8984 21790 8996
rect 22097 8993 22109 8996
rect 22143 9024 22155 9027
rect 22925 9027 22983 9033
rect 22925 9024 22937 9027
rect 22143 8996 22937 9024
rect 22143 8993 22155 8996
rect 22097 8987 22155 8993
rect 22925 8993 22937 8996
rect 22971 8993 22983 9027
rect 31478 9024 31484 9036
rect 31439 8996 31484 9024
rect 22925 8987 22983 8993
rect 31478 8984 31484 8996
rect 31536 8984 31542 9036
rect 15473 8959 15531 8965
rect 15473 8956 15485 8959
rect 15436 8928 15485 8956
rect 15436 8916 15442 8928
rect 15473 8925 15485 8928
rect 15519 8925 15531 8959
rect 15654 8956 15660 8968
rect 15615 8928 15660 8956
rect 15473 8919 15531 8925
rect 15654 8916 15660 8928
rect 15712 8916 15718 8968
rect 16114 8956 16120 8968
rect 16075 8928 16120 8956
rect 16114 8916 16120 8928
rect 16172 8916 16178 8968
rect 16298 8956 16304 8968
rect 16259 8928 16304 8956
rect 16298 8916 16304 8928
rect 16356 8916 16362 8968
rect 18046 8916 18052 8968
rect 18104 8956 18110 8968
rect 18141 8959 18199 8965
rect 18141 8956 18153 8959
rect 18104 8928 18153 8956
rect 18104 8916 18110 8928
rect 18141 8925 18153 8928
rect 18187 8925 18199 8959
rect 18141 8919 18199 8925
rect 20990 8916 20996 8968
rect 21048 8956 21054 8968
rect 21453 8959 21511 8965
rect 21453 8956 21465 8959
rect 21048 8928 21465 8956
rect 21048 8916 21054 8928
rect 21453 8925 21465 8928
rect 21499 8925 21511 8959
rect 21453 8919 21511 8925
rect 21542 8916 21548 8968
rect 21600 8956 21606 8968
rect 22281 8959 22339 8965
rect 21600 8928 22094 8956
rect 21600 8916 21606 8928
rect 20073 8891 20131 8897
rect 20073 8857 20085 8891
rect 20119 8888 20131 8891
rect 20714 8888 20720 8900
rect 20119 8860 20720 8888
rect 20119 8857 20131 8860
rect 20073 8851 20131 8857
rect 20714 8848 20720 8860
rect 20772 8848 20778 8900
rect 22066 8888 22094 8928
rect 22281 8925 22293 8959
rect 22327 8925 22339 8959
rect 22281 8919 22339 8925
rect 22296 8888 22324 8919
rect 22646 8916 22652 8968
rect 22704 8956 22710 8968
rect 23109 8959 23167 8965
rect 23109 8956 23121 8959
rect 22704 8928 23121 8956
rect 22704 8916 22710 8928
rect 23109 8925 23121 8928
rect 23155 8925 23167 8959
rect 23109 8919 23167 8925
rect 25498 8916 25504 8968
rect 25556 8956 25562 8968
rect 26329 8959 26387 8965
rect 26329 8956 26341 8959
rect 25556 8928 26341 8956
rect 25556 8916 25562 8928
rect 26329 8925 26341 8928
rect 26375 8925 26387 8959
rect 26329 8919 26387 8925
rect 26513 8959 26571 8965
rect 26513 8925 26525 8959
rect 26559 8956 26571 8959
rect 26973 8959 27031 8965
rect 26973 8956 26985 8959
rect 26559 8928 26985 8956
rect 26559 8925 26571 8928
rect 26513 8919 26571 8925
rect 26973 8925 26985 8928
rect 27019 8925 27031 8959
rect 26973 8919 27031 8925
rect 28353 8959 28411 8965
rect 28353 8925 28365 8959
rect 28399 8956 28411 8959
rect 28626 8956 28632 8968
rect 28399 8928 28632 8956
rect 28399 8925 28411 8928
rect 28353 8919 28411 8925
rect 28626 8916 28632 8928
rect 28684 8916 28690 8968
rect 29546 8956 29552 8968
rect 29507 8928 29552 8956
rect 29546 8916 29552 8928
rect 29604 8916 29610 8968
rect 31748 8959 31806 8965
rect 31748 8925 31760 8959
rect 31794 8956 31806 8959
rect 32122 8956 32128 8968
rect 31794 8928 32128 8956
rect 31794 8925 31806 8928
rect 31748 8919 31806 8925
rect 32122 8916 32128 8928
rect 32180 8916 32186 8968
rect 22066 8860 22324 8888
rect 26145 8891 26203 8897
rect 26145 8857 26157 8891
rect 26191 8888 26203 8891
rect 26234 8888 26240 8900
rect 26191 8860 26240 8888
rect 26191 8857 26203 8860
rect 26145 8851 26203 8857
rect 26234 8848 26240 8860
rect 26292 8848 26298 8900
rect 15562 8820 15568 8832
rect 15523 8792 15568 8820
rect 15562 8780 15568 8792
rect 15620 8780 15626 8832
rect 19426 8780 19432 8832
rect 19484 8820 19490 8832
rect 19705 8823 19763 8829
rect 19705 8820 19717 8823
rect 19484 8792 19717 8820
rect 19484 8780 19490 8792
rect 19705 8789 19717 8792
rect 19751 8789 19763 8823
rect 19705 8783 19763 8789
rect 19873 8823 19931 8829
rect 19873 8789 19885 8823
rect 19919 8820 19931 8823
rect 20622 8820 20628 8832
rect 19919 8792 20628 8820
rect 19919 8789 19931 8792
rect 19873 8783 19931 8789
rect 20622 8780 20628 8792
rect 20680 8780 20686 8832
rect 23293 8823 23351 8829
rect 23293 8789 23305 8823
rect 23339 8820 23351 8823
rect 23750 8820 23756 8832
rect 23339 8792 23756 8820
rect 23339 8789 23351 8792
rect 23293 8783 23351 8789
rect 23750 8780 23756 8792
rect 23808 8780 23814 8832
rect 27154 8820 27160 8832
rect 27115 8792 27160 8820
rect 27154 8780 27160 8792
rect 27212 8780 27218 8832
rect 28997 8823 29055 8829
rect 28997 8789 29009 8823
rect 29043 8820 29055 8823
rect 29178 8820 29184 8832
rect 29043 8792 29184 8820
rect 29043 8789 29055 8792
rect 28997 8783 29055 8789
rect 29178 8780 29184 8792
rect 29236 8780 29242 8832
rect 31294 8780 31300 8832
rect 31352 8820 31358 8832
rect 32861 8823 32919 8829
rect 32861 8820 32873 8823
rect 31352 8792 32873 8820
rect 31352 8780 31358 8792
rect 32861 8789 32873 8792
rect 32907 8789 32919 8823
rect 32861 8783 32919 8789
rect 1104 8730 42872 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 42872 8730
rect 1104 8656 42872 8678
rect 16114 8616 16120 8628
rect 16075 8588 16120 8616
rect 16114 8576 16120 8588
rect 16172 8576 16178 8628
rect 20901 8619 20959 8625
rect 20901 8585 20913 8619
rect 20947 8616 20959 8619
rect 21542 8616 21548 8628
rect 20947 8588 21548 8616
rect 20947 8585 20959 8588
rect 20901 8579 20959 8585
rect 21542 8576 21548 8588
rect 21600 8576 21606 8628
rect 22186 8616 22192 8628
rect 22147 8588 22192 8616
rect 22186 8576 22192 8588
rect 22244 8576 22250 8628
rect 24397 8619 24455 8625
rect 24397 8585 24409 8619
rect 24443 8616 24455 8619
rect 25222 8616 25228 8628
rect 24443 8588 25228 8616
rect 24443 8585 24455 8588
rect 24397 8579 24455 8585
rect 25222 8576 25228 8588
rect 25280 8576 25286 8628
rect 28626 8616 28632 8628
rect 28587 8588 28632 8616
rect 28626 8576 28632 8588
rect 28684 8576 28690 8628
rect 30469 8619 30527 8625
rect 30469 8585 30481 8619
rect 30515 8616 30527 8619
rect 30558 8616 30564 8628
rect 30515 8588 30564 8616
rect 30515 8585 30527 8588
rect 30469 8579 30527 8585
rect 30558 8576 30564 8588
rect 30616 8616 30622 8628
rect 30616 8588 30972 8616
rect 30616 8576 30622 8588
rect 1949 8551 2007 8557
rect 1949 8517 1961 8551
rect 1995 8548 2007 8551
rect 2866 8548 2872 8560
rect 1995 8520 2872 8548
rect 1995 8517 2007 8520
rect 1949 8511 2007 8517
rect 2866 8508 2872 8520
rect 2924 8508 2930 8560
rect 15004 8551 15062 8557
rect 15004 8517 15016 8551
rect 15050 8548 15062 8551
rect 15562 8548 15568 8560
rect 15050 8520 15568 8548
rect 15050 8517 15062 8520
rect 15004 8511 15062 8517
rect 15562 8508 15568 8520
rect 15620 8508 15626 8560
rect 16298 8508 16304 8560
rect 16356 8548 16362 8560
rect 19426 8548 19432 8560
rect 16356 8520 19432 8548
rect 16356 8508 16362 8520
rect 19426 8508 19432 8520
rect 19484 8548 19490 8560
rect 19889 8551 19947 8557
rect 19484 8520 19564 8548
rect 19484 8508 19490 8520
rect 1762 8480 1768 8492
rect 1723 8452 1768 8480
rect 1762 8440 1768 8452
rect 1820 8440 1826 8492
rect 14734 8480 14740 8492
rect 14695 8452 14740 8480
rect 14734 8440 14740 8452
rect 14792 8440 14798 8492
rect 17497 8483 17555 8489
rect 17497 8449 17509 8483
rect 17543 8480 17555 8483
rect 17862 8480 17868 8492
rect 17543 8452 17868 8480
rect 17543 8449 17555 8452
rect 17497 8443 17555 8449
rect 17862 8440 17868 8452
rect 17920 8440 17926 8492
rect 19536 8489 19564 8520
rect 19889 8517 19901 8551
rect 19935 8548 19947 8551
rect 20533 8551 20591 8557
rect 20533 8548 20545 8551
rect 19935 8520 20545 8548
rect 19935 8517 19947 8520
rect 19889 8511 19947 8517
rect 20533 8517 20545 8520
rect 20579 8517 20591 8551
rect 20533 8511 20591 8517
rect 20732 8520 22048 8548
rect 20732 8492 20760 8520
rect 22020 8492 22048 8520
rect 22830 8508 22836 8560
rect 22888 8548 22894 8560
rect 23262 8551 23320 8557
rect 23262 8548 23274 8551
rect 22888 8520 23274 8548
rect 22888 8508 22894 8520
rect 23262 8517 23274 8520
rect 23308 8517 23320 8551
rect 23262 8511 23320 8517
rect 27154 8508 27160 8560
rect 27212 8548 27218 8560
rect 27494 8551 27552 8557
rect 27494 8548 27506 8551
rect 27212 8520 27506 8548
rect 27212 8508 27218 8520
rect 27494 8517 27506 8520
rect 27540 8517 27552 8551
rect 30834 8548 30840 8560
rect 27494 8511 27552 8517
rect 29104 8520 30840 8548
rect 19521 8483 19579 8489
rect 19521 8449 19533 8483
rect 19567 8449 19579 8483
rect 20714 8480 20720 8492
rect 20675 8452 20720 8480
rect 19521 8443 19579 8449
rect 20714 8440 20720 8452
rect 20772 8440 20778 8492
rect 20990 8440 20996 8492
rect 21048 8480 21054 8492
rect 21048 8452 21093 8480
rect 21048 8440 21054 8452
rect 21726 8440 21732 8492
rect 21784 8480 21790 8492
rect 21821 8483 21879 8489
rect 21821 8480 21833 8483
rect 21784 8452 21833 8480
rect 21784 8440 21790 8452
rect 21821 8449 21833 8452
rect 21867 8449 21879 8483
rect 22002 8480 22008 8492
rect 21915 8452 22008 8480
rect 21821 8443 21879 8449
rect 22002 8440 22008 8452
rect 22060 8440 22066 8492
rect 23014 8480 23020 8492
rect 22975 8452 23020 8480
rect 23014 8440 23020 8452
rect 23072 8440 23078 8492
rect 27249 8483 27307 8489
rect 27249 8449 27261 8483
rect 27295 8480 27307 8483
rect 27338 8480 27344 8492
rect 27295 8452 27344 8480
rect 27295 8449 27307 8452
rect 27249 8443 27307 8449
rect 27338 8440 27344 8452
rect 27396 8440 27402 8492
rect 29104 8489 29132 8520
rect 30834 8508 30840 8520
rect 30892 8508 30898 8560
rect 30944 8557 30972 8588
rect 30929 8551 30987 8557
rect 30929 8517 30941 8551
rect 30975 8517 30987 8551
rect 30929 8511 30987 8517
rect 29089 8483 29147 8489
rect 29089 8449 29101 8483
rect 29135 8449 29147 8483
rect 29089 8443 29147 8449
rect 29178 8440 29184 8492
rect 29236 8480 29242 8492
rect 29345 8483 29403 8489
rect 29345 8480 29357 8483
rect 29236 8452 29357 8480
rect 29236 8440 29242 8452
rect 29345 8449 29357 8452
rect 29391 8449 29403 8483
rect 29345 8443 29403 8449
rect 2774 8372 2780 8424
rect 2832 8412 2838 8424
rect 2832 8384 2877 8412
rect 2832 8372 2838 8384
rect 17126 8372 17132 8424
rect 17184 8412 17190 8424
rect 17221 8415 17279 8421
rect 17221 8412 17233 8415
rect 17184 8384 17233 8412
rect 17184 8372 17190 8384
rect 17221 8381 17233 8384
rect 17267 8381 17279 8415
rect 17221 8375 17279 8381
rect 17402 8372 17408 8424
rect 17460 8412 17466 8424
rect 18233 8415 18291 8421
rect 18233 8412 18245 8415
rect 17460 8384 18245 8412
rect 17460 8372 17466 8384
rect 18233 8381 18245 8384
rect 18279 8412 18291 8415
rect 21008 8412 21036 8440
rect 18279 8384 21036 8412
rect 18279 8381 18291 8384
rect 18233 8375 18291 8381
rect 30282 8372 30288 8424
rect 30340 8412 30346 8424
rect 31389 8415 31447 8421
rect 31389 8412 31401 8415
rect 30340 8384 31401 8412
rect 30340 8372 30346 8384
rect 31389 8381 31401 8384
rect 31435 8381 31447 8415
rect 31389 8375 31447 8381
rect 18509 8347 18567 8353
rect 18509 8313 18521 8347
rect 18555 8344 18567 8347
rect 20073 8347 20131 8353
rect 18555 8316 18828 8344
rect 18555 8313 18567 8316
rect 18509 8307 18567 8313
rect 17218 8236 17224 8288
rect 17276 8276 17282 8288
rect 17313 8279 17371 8285
rect 17313 8276 17325 8279
rect 17276 8248 17325 8276
rect 17276 8236 17282 8248
rect 17313 8245 17325 8248
rect 17359 8245 17371 8279
rect 17313 8239 17371 8245
rect 18598 8236 18604 8288
rect 18656 8276 18662 8288
rect 18693 8279 18751 8285
rect 18693 8276 18705 8279
rect 18656 8248 18705 8276
rect 18656 8236 18662 8248
rect 18693 8245 18705 8248
rect 18739 8245 18751 8279
rect 18800 8276 18828 8316
rect 20073 8313 20085 8347
rect 20119 8344 20131 8347
rect 20254 8344 20260 8356
rect 20119 8316 20260 8344
rect 20119 8313 20131 8316
rect 20073 8307 20131 8313
rect 20254 8304 20260 8316
rect 20312 8304 20318 8356
rect 31294 8344 31300 8356
rect 31255 8316 31300 8344
rect 31294 8304 31300 8316
rect 31352 8304 31358 8356
rect 19150 8276 19156 8288
rect 18800 8248 19156 8276
rect 18693 8239 18751 8245
rect 19150 8236 19156 8248
rect 19208 8276 19214 8288
rect 19889 8279 19947 8285
rect 19889 8276 19901 8279
rect 19208 8248 19901 8276
rect 19208 8236 19214 8248
rect 19889 8245 19901 8248
rect 19935 8245 19947 8279
rect 19889 8239 19947 8245
rect 1104 8186 42872 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 42872 8186
rect 1104 8112 42872 8134
rect 15654 8032 15660 8084
rect 15712 8072 15718 8084
rect 16025 8075 16083 8081
rect 16025 8072 16037 8075
rect 15712 8044 16037 8072
rect 15712 8032 15718 8044
rect 16025 8041 16037 8044
rect 16071 8041 16083 8075
rect 16025 8035 16083 8041
rect 16117 8075 16175 8081
rect 16117 8041 16129 8075
rect 16163 8072 16175 8075
rect 16298 8072 16304 8084
rect 16163 8044 16304 8072
rect 16163 8041 16175 8044
rect 16117 8035 16175 8041
rect 16298 8032 16304 8044
rect 16356 8032 16362 8084
rect 17862 8032 17868 8084
rect 17920 8072 17926 8084
rect 18233 8075 18291 8081
rect 18233 8072 18245 8075
rect 17920 8044 18245 8072
rect 17920 8032 17926 8044
rect 18233 8041 18245 8044
rect 18279 8041 18291 8075
rect 20622 8072 20628 8084
rect 20583 8044 20628 8072
rect 18233 8035 18291 8041
rect 20622 8032 20628 8044
rect 20680 8032 20686 8084
rect 22002 8032 22008 8084
rect 22060 8072 22066 8084
rect 22465 8075 22523 8081
rect 22465 8072 22477 8075
rect 22060 8044 22477 8072
rect 22060 8032 22066 8044
rect 22465 8041 22477 8044
rect 22511 8041 22523 8075
rect 22465 8035 22523 8041
rect 23109 8075 23167 8081
rect 23109 8041 23121 8075
rect 23155 8072 23167 8075
rect 23566 8072 23572 8084
rect 23155 8044 23572 8072
rect 23155 8041 23167 8044
rect 23109 8035 23167 8041
rect 23566 8032 23572 8044
rect 23624 8032 23630 8084
rect 15930 7936 15936 7948
rect 15891 7908 15936 7936
rect 15930 7896 15936 7908
rect 15988 7896 15994 7948
rect 16850 7936 16856 7948
rect 16811 7908 16856 7936
rect 16850 7896 16856 7908
rect 16908 7896 16914 7948
rect 23014 7936 23020 7948
rect 22664 7908 23020 7936
rect 16114 7828 16120 7880
rect 16172 7868 16178 7880
rect 16209 7871 16267 7877
rect 16209 7868 16221 7871
rect 16172 7840 16221 7868
rect 16172 7828 16178 7840
rect 16209 7837 16221 7840
rect 16255 7837 16267 7871
rect 16868 7868 16896 7896
rect 19245 7871 19303 7877
rect 19245 7868 19257 7871
rect 16868 7840 19257 7868
rect 16209 7831 16267 7837
rect 19245 7837 19257 7840
rect 19291 7837 19303 7871
rect 19245 7831 19303 7837
rect 21085 7871 21143 7877
rect 21085 7837 21097 7871
rect 21131 7868 21143 7871
rect 22664 7868 22692 7908
rect 23014 7896 23020 7908
rect 23072 7896 23078 7948
rect 25314 7936 25320 7948
rect 25275 7908 25320 7936
rect 25314 7896 25320 7908
rect 25372 7896 25378 7948
rect 22922 7868 22928 7880
rect 21131 7840 22692 7868
rect 22883 7840 22928 7868
rect 21131 7837 21143 7840
rect 21085 7831 21143 7837
rect 22922 7828 22928 7840
rect 22980 7828 22986 7880
rect 23750 7868 23756 7880
rect 23711 7840 23756 7868
rect 23750 7828 23756 7840
rect 23808 7828 23814 7880
rect 41598 7828 41604 7880
rect 41656 7868 41662 7880
rect 41693 7871 41751 7877
rect 41693 7868 41705 7871
rect 41656 7840 41705 7868
rect 41656 7828 41662 7840
rect 41693 7837 41705 7840
rect 41739 7837 41751 7871
rect 41693 7831 41751 7837
rect 17126 7809 17132 7812
rect 17120 7763 17132 7809
rect 17184 7800 17190 7812
rect 17184 7772 17220 7800
rect 17126 7760 17132 7763
rect 17184 7760 17190 7772
rect 18782 7760 18788 7812
rect 18840 7800 18846 7812
rect 19490 7803 19548 7809
rect 19490 7800 19502 7803
rect 18840 7772 19502 7800
rect 18840 7760 18846 7772
rect 19490 7769 19502 7772
rect 19536 7769 19548 7803
rect 19490 7763 19548 7769
rect 20714 7760 20720 7812
rect 20772 7800 20778 7812
rect 25590 7809 25596 7812
rect 21330 7803 21388 7809
rect 21330 7800 21342 7803
rect 20772 7772 21342 7800
rect 20772 7760 20778 7772
rect 21330 7769 21342 7772
rect 21376 7769 21388 7803
rect 21330 7763 21388 7769
rect 25584 7763 25596 7809
rect 25648 7800 25654 7812
rect 25648 7772 25684 7800
rect 25590 7760 25596 7763
rect 25648 7760 25654 7772
rect 23566 7732 23572 7744
rect 23527 7704 23572 7732
rect 23566 7692 23572 7704
rect 23624 7692 23630 7744
rect 40494 7692 40500 7744
rect 40552 7732 40558 7744
rect 41601 7735 41659 7741
rect 41601 7732 41613 7735
rect 40552 7704 41613 7732
rect 40552 7692 40558 7704
rect 41601 7701 41613 7704
rect 41647 7701 41659 7735
rect 41601 7695 41659 7701
rect 1104 7642 42872 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 42872 7642
rect 1104 7568 42872 7590
rect 17313 7531 17371 7537
rect 17313 7497 17325 7531
rect 17359 7528 17371 7531
rect 17862 7528 17868 7540
rect 17359 7500 17868 7528
rect 17359 7497 17371 7500
rect 17313 7491 17371 7497
rect 17862 7488 17868 7500
rect 17920 7488 17926 7540
rect 18782 7528 18788 7540
rect 18743 7500 18788 7528
rect 18782 7488 18788 7500
rect 18840 7488 18846 7540
rect 24397 7531 24455 7537
rect 24397 7497 24409 7531
rect 24443 7497 24455 7531
rect 24397 7491 24455 7497
rect 25501 7531 25559 7537
rect 25501 7497 25513 7531
rect 25547 7528 25559 7531
rect 25590 7528 25596 7540
rect 25547 7500 25596 7528
rect 25547 7497 25559 7500
rect 25501 7491 25559 7497
rect 17129 7463 17187 7469
rect 17129 7429 17141 7463
rect 17175 7460 17187 7463
rect 17218 7460 17224 7472
rect 17175 7432 17224 7460
rect 17175 7429 17187 7432
rect 17129 7423 17187 7429
rect 17218 7420 17224 7432
rect 17276 7420 17282 7472
rect 23284 7463 23342 7469
rect 23284 7429 23296 7463
rect 23330 7460 23342 7463
rect 23566 7460 23572 7472
rect 23330 7432 23572 7460
rect 23330 7429 23342 7432
rect 23284 7423 23342 7429
rect 23566 7420 23572 7432
rect 23624 7420 23630 7472
rect 17402 7352 17408 7404
rect 17460 7392 17466 7404
rect 18598 7392 18604 7404
rect 17460 7364 17505 7392
rect 18559 7364 18604 7392
rect 17460 7352 17466 7364
rect 18598 7352 18604 7364
rect 18656 7352 18662 7404
rect 19981 7395 20039 7401
rect 19981 7361 19993 7395
rect 20027 7392 20039 7395
rect 20622 7392 20628 7404
rect 20027 7364 20628 7392
rect 20027 7361 20039 7364
rect 19981 7355 20039 7361
rect 20622 7352 20628 7364
rect 20680 7352 20686 7404
rect 23014 7392 23020 7404
rect 22975 7364 23020 7392
rect 23014 7352 23020 7364
rect 23072 7352 23078 7404
rect 24412 7392 24440 7491
rect 25590 7488 25596 7500
rect 25648 7488 25654 7540
rect 24857 7395 24915 7401
rect 24857 7392 24869 7395
rect 24412 7364 24869 7392
rect 24857 7361 24869 7364
rect 24903 7392 24915 7395
rect 25498 7392 25504 7404
rect 24903 7364 25504 7392
rect 24903 7361 24915 7364
rect 24857 7355 24915 7361
rect 25498 7352 25504 7364
rect 25556 7352 25562 7404
rect 41874 7392 41880 7404
rect 41835 7364 41880 7392
rect 41874 7352 41880 7364
rect 41932 7352 41938 7404
rect 20257 7327 20315 7333
rect 20257 7293 20269 7327
rect 20303 7324 20315 7327
rect 20990 7324 20996 7336
rect 20303 7296 20996 7324
rect 20303 7293 20315 7296
rect 20257 7287 20315 7293
rect 20990 7284 20996 7296
rect 21048 7284 21054 7336
rect 17126 7256 17132 7268
rect 17087 7228 17132 7256
rect 17126 7216 17132 7228
rect 17184 7216 17190 7268
rect 24578 7216 24584 7268
rect 24636 7256 24642 7268
rect 41693 7259 41751 7265
rect 41693 7256 41705 7259
rect 24636 7228 41705 7256
rect 24636 7216 24642 7228
rect 41693 7225 41705 7228
rect 41739 7225 41751 7259
rect 41693 7219 41751 7225
rect 40954 7188 40960 7200
rect 40915 7160 40960 7188
rect 40954 7148 40960 7160
rect 41012 7148 41018 7200
rect 1104 7098 42872 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 42872 7098
rect 1104 7024 42872 7046
rect 4062 6808 4068 6860
rect 4120 6848 4126 6860
rect 13630 6848 13636 6860
rect 4120 6820 13636 6848
rect 4120 6808 4126 6820
rect 13630 6808 13636 6820
rect 13688 6808 13694 6860
rect 40313 6851 40371 6857
rect 40313 6817 40325 6851
rect 40359 6848 40371 6851
rect 40954 6848 40960 6860
rect 40359 6820 40960 6848
rect 40359 6817 40371 6820
rect 40313 6811 40371 6817
rect 40954 6808 40960 6820
rect 41012 6808 41018 6860
rect 4249 6783 4307 6789
rect 4249 6749 4261 6783
rect 4295 6780 4307 6783
rect 4614 6780 4620 6792
rect 4295 6752 4620 6780
rect 4295 6749 4307 6752
rect 4249 6743 4307 6749
rect 4614 6740 4620 6752
rect 4672 6740 4678 6792
rect 20254 6780 20260 6792
rect 20215 6752 20260 6780
rect 20254 6740 20260 6752
rect 20312 6740 20318 6792
rect 40494 6712 40500 6724
rect 40455 6684 40500 6712
rect 40494 6672 40500 6684
rect 40552 6672 40558 6724
rect 42150 6712 42156 6724
rect 42111 6684 42156 6712
rect 42150 6672 42156 6684
rect 42208 6672 42214 6724
rect 4154 6644 4160 6656
rect 4115 6616 4160 6644
rect 4154 6604 4160 6616
rect 4212 6604 4218 6656
rect 20441 6647 20499 6653
rect 20441 6613 20453 6647
rect 20487 6644 20499 6647
rect 20714 6644 20720 6656
rect 20487 6616 20720 6644
rect 20487 6613 20499 6616
rect 20441 6607 20499 6613
rect 20714 6604 20720 6616
rect 20772 6604 20778 6656
rect 1104 6554 42872 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 42872 6554
rect 1104 6480 42872 6502
rect 7650 6440 7656 6452
rect 2884 6412 7656 6440
rect 2884 6313 2912 6412
rect 7650 6400 7656 6412
rect 7708 6400 7714 6452
rect 4154 6372 4160 6384
rect 4115 6344 4160 6372
rect 4154 6332 4160 6344
rect 4212 6332 4218 6384
rect 2869 6307 2927 6313
rect 2869 6273 2881 6307
rect 2915 6273 2927 6307
rect 2869 6267 2927 6273
rect 3970 6236 3976 6248
rect 3931 6208 3976 6236
rect 3970 6196 3976 6208
rect 4028 6196 4034 6248
rect 5074 6236 5080 6248
rect 5035 6208 5080 6236
rect 5074 6196 5080 6208
rect 5132 6196 5138 6248
rect 1394 6100 1400 6112
rect 1355 6072 1400 6100
rect 1394 6060 1400 6072
rect 1452 6060 1458 6112
rect 1946 6060 1952 6112
rect 2004 6100 2010 6112
rect 2041 6103 2099 6109
rect 2041 6100 2053 6103
rect 2004 6072 2053 6100
rect 2004 6060 2010 6072
rect 2041 6069 2053 6072
rect 2087 6069 2099 6103
rect 2041 6063 2099 6069
rect 2774 6060 2780 6112
rect 2832 6100 2838 6112
rect 2832 6072 2877 6100
rect 2832 6060 2838 6072
rect 40310 6060 40316 6112
rect 40368 6100 40374 6112
rect 40957 6103 41015 6109
rect 40957 6100 40969 6103
rect 40368 6072 40969 6100
rect 40368 6060 40374 6072
rect 40957 6069 40969 6072
rect 41003 6069 41015 6103
rect 41782 6100 41788 6112
rect 41743 6072 41788 6100
rect 40957 6063 41015 6069
rect 41782 6060 41788 6072
rect 41840 6060 41846 6112
rect 1104 6010 42872 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 42872 6010
rect 1104 5936 42872 5958
rect 3970 5856 3976 5908
rect 4028 5896 4034 5908
rect 4433 5899 4491 5905
rect 4433 5896 4445 5899
rect 4028 5868 4445 5896
rect 4028 5856 4034 5868
rect 4433 5865 4445 5868
rect 4479 5865 4491 5899
rect 4433 5859 4491 5865
rect 1394 5760 1400 5772
rect 1355 5732 1400 5760
rect 1394 5720 1400 5732
rect 1452 5720 1458 5772
rect 1854 5760 1860 5772
rect 1815 5732 1860 5760
rect 1854 5720 1860 5732
rect 1912 5720 1918 5772
rect 2130 5720 2136 5772
rect 2188 5760 2194 5772
rect 40865 5763 40923 5769
rect 2188 5732 22094 5760
rect 2188 5720 2194 5732
rect 3973 5695 4031 5701
rect 3973 5661 3985 5695
rect 4019 5692 4031 5695
rect 4982 5692 4988 5704
rect 4019 5664 4988 5692
rect 4019 5661 4031 5664
rect 3973 5655 4031 5661
rect 4982 5652 4988 5664
rect 5040 5652 5046 5704
rect 22066 5692 22094 5732
rect 40865 5729 40877 5763
rect 40911 5760 40923 5763
rect 41690 5760 41696 5772
rect 40911 5732 41696 5760
rect 40911 5729 40923 5732
rect 40865 5723 40923 5729
rect 41690 5720 41696 5732
rect 41748 5720 41754 5772
rect 37829 5695 37887 5701
rect 37829 5692 37841 5695
rect 22066 5664 37841 5692
rect 37829 5661 37841 5664
rect 37875 5661 37887 5695
rect 37829 5655 37887 5661
rect 38470 5652 38476 5704
rect 38528 5692 38534 5704
rect 38565 5695 38623 5701
rect 38565 5692 38577 5695
rect 38528 5664 38577 5692
rect 38528 5652 38534 5664
rect 38565 5661 38577 5664
rect 38611 5661 38623 5695
rect 39850 5692 39856 5704
rect 39811 5664 39856 5692
rect 38565 5655 38623 5661
rect 39850 5652 39856 5664
rect 39908 5652 39914 5704
rect 41230 5652 41236 5704
rect 41288 5692 41294 5704
rect 41325 5695 41383 5701
rect 41325 5692 41337 5695
rect 41288 5664 41337 5692
rect 41288 5652 41294 5664
rect 41325 5661 41337 5664
rect 41371 5661 41383 5695
rect 41966 5692 41972 5704
rect 41927 5664 41972 5692
rect 41325 5655 41383 5661
rect 41966 5652 41972 5664
rect 42024 5652 42030 5704
rect 1578 5624 1584 5636
rect 1539 5596 1584 5624
rect 1578 5584 1584 5596
rect 1636 5584 1642 5636
rect 37921 5559 37979 5565
rect 37921 5525 37933 5559
rect 37967 5556 37979 5559
rect 38654 5556 38660 5568
rect 37967 5528 38660 5556
rect 37967 5525 37979 5528
rect 37921 5519 37979 5525
rect 38654 5516 38660 5528
rect 38712 5516 38718 5568
rect 41417 5559 41475 5565
rect 41417 5525 41429 5559
rect 41463 5556 41475 5559
rect 41966 5556 41972 5568
rect 41463 5528 41972 5556
rect 41463 5525 41475 5528
rect 41417 5519 41475 5525
rect 41966 5516 41972 5528
rect 42024 5516 42030 5568
rect 42058 5516 42064 5568
rect 42116 5556 42122 5568
rect 42116 5528 42161 5556
rect 42116 5516 42122 5528
rect 1104 5466 42872 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 42872 5466
rect 1104 5392 42872 5414
rect 2133 5287 2191 5293
rect 2133 5253 2145 5287
rect 2179 5284 2191 5287
rect 2774 5284 2780 5296
rect 2179 5256 2780 5284
rect 2179 5253 2191 5256
rect 2133 5247 2191 5253
rect 2774 5244 2780 5256
rect 2832 5244 2838 5296
rect 38654 5284 38660 5296
rect 38615 5256 38660 5284
rect 38654 5244 38660 5256
rect 38712 5244 38718 5296
rect 1946 5216 1952 5228
rect 1907 5188 1952 5216
rect 1946 5176 1952 5188
rect 2004 5176 2010 5228
rect 38470 5216 38476 5228
rect 38431 5188 38476 5216
rect 38470 5176 38476 5188
rect 38528 5176 38534 5228
rect 40957 5219 41015 5225
rect 40957 5185 40969 5219
rect 41003 5216 41015 5219
rect 41046 5216 41052 5228
rect 41003 5188 41052 5216
rect 41003 5185 41015 5188
rect 40957 5179 41015 5185
rect 41046 5176 41052 5188
rect 41104 5176 41110 5228
rect 41414 5216 41420 5228
rect 41375 5188 41420 5216
rect 41414 5176 41420 5188
rect 41472 5176 41478 5228
rect 2774 5108 2780 5160
rect 2832 5148 2838 5160
rect 40313 5151 40371 5157
rect 2832 5120 2877 5148
rect 2832 5108 2838 5120
rect 40313 5117 40325 5151
rect 40359 5148 40371 5151
rect 43162 5148 43168 5160
rect 40359 5120 43168 5148
rect 40359 5117 40371 5120
rect 40313 5111 40371 5117
rect 43162 5108 43168 5120
rect 43220 5108 43226 5160
rect 4249 5015 4307 5021
rect 4249 4981 4261 5015
rect 4295 5012 4307 5015
rect 4614 5012 4620 5024
rect 4295 4984 4620 5012
rect 4295 4981 4307 4984
rect 4249 4975 4307 4981
rect 4614 4972 4620 4984
rect 4672 4972 4678 5024
rect 40034 4972 40040 5024
rect 40092 5012 40098 5024
rect 40865 5015 40923 5021
rect 40865 5012 40877 5015
rect 40092 4984 40877 5012
rect 40092 4972 40098 4984
rect 40865 4981 40877 4984
rect 40911 4981 40923 5015
rect 41506 5012 41512 5024
rect 41467 4984 41512 5012
rect 40865 4975 40923 4981
rect 41506 4972 41512 4984
rect 41564 4972 41570 5024
rect 1104 4922 42872 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 42872 4922
rect 1104 4848 42872 4870
rect 1578 4768 1584 4820
rect 1636 4808 1642 4820
rect 2133 4811 2191 4817
rect 2133 4808 2145 4811
rect 1636 4780 2145 4808
rect 1636 4768 1642 4780
rect 2133 4777 2145 4780
rect 2179 4777 2191 4811
rect 2133 4771 2191 4777
rect 4798 4740 4804 4752
rect 2746 4712 4804 4740
rect 2746 4672 2774 4712
rect 4798 4700 4804 4712
rect 4856 4700 4862 4752
rect 2240 4644 2774 4672
rect 4617 4675 4675 4681
rect 1397 4607 1455 4613
rect 1397 4573 1409 4607
rect 1443 4604 1455 4607
rect 1486 4604 1492 4616
rect 1443 4576 1492 4604
rect 1443 4573 1455 4576
rect 1397 4567 1455 4573
rect 1486 4564 1492 4576
rect 1544 4564 1550 4616
rect 2130 4564 2136 4616
rect 2188 4604 2194 4616
rect 2240 4613 2268 4644
rect 4617 4641 4629 4675
rect 4663 4672 4675 4675
rect 5534 4672 5540 4684
rect 4663 4644 5540 4672
rect 4663 4641 4675 4644
rect 4617 4635 4675 4641
rect 5534 4632 5540 4644
rect 5592 4632 5598 4684
rect 40310 4672 40316 4684
rect 40271 4644 40316 4672
rect 40310 4632 40316 4644
rect 40368 4632 40374 4684
rect 40497 4675 40555 4681
rect 40497 4641 40509 4675
rect 40543 4672 40555 4675
rect 41506 4672 41512 4684
rect 40543 4644 41512 4672
rect 40543 4641 40555 4644
rect 40497 4635 40555 4641
rect 41506 4632 41512 4644
rect 41564 4632 41570 4684
rect 41874 4672 41880 4684
rect 41835 4644 41880 4672
rect 41874 4632 41880 4644
rect 41932 4632 41938 4684
rect 2225 4607 2283 4613
rect 2225 4604 2237 4607
rect 2188 4576 2237 4604
rect 2188 4564 2194 4576
rect 2225 4573 2237 4576
rect 2271 4573 2283 4607
rect 2225 4567 2283 4573
rect 2869 4607 2927 4613
rect 2869 4573 2881 4607
rect 2915 4604 2927 4607
rect 3234 4604 3240 4616
rect 2915 4576 3240 4604
rect 2915 4573 2927 4576
rect 2869 4567 2927 4573
rect 3234 4564 3240 4576
rect 3292 4564 3298 4616
rect 3973 4607 4031 4613
rect 3973 4573 3985 4607
rect 4019 4573 4031 4607
rect 3973 4567 4031 4573
rect 3988 4536 4016 4567
rect 4706 4564 4712 4616
rect 4764 4604 4770 4616
rect 5077 4607 5135 4613
rect 5077 4604 5089 4607
rect 4764 4576 5089 4604
rect 4764 4564 4770 4576
rect 5077 4573 5089 4576
rect 5123 4573 5135 4607
rect 36722 4604 36728 4616
rect 36683 4576 36728 4604
rect 5077 4567 5135 4573
rect 36722 4564 36728 4576
rect 36780 4564 36786 4616
rect 37550 4564 37556 4616
rect 37608 4604 37614 4616
rect 37829 4607 37887 4613
rect 37829 4604 37841 4607
rect 37608 4576 37841 4604
rect 37608 4564 37614 4576
rect 37829 4573 37841 4576
rect 37875 4573 37887 4607
rect 37829 4567 37887 4573
rect 38657 4607 38715 4613
rect 38657 4573 38669 4607
rect 38703 4604 38715 4607
rect 39022 4604 39028 4616
rect 38703 4576 39028 4604
rect 38703 4573 38715 4576
rect 38657 4567 38715 4573
rect 39022 4564 39028 4576
rect 39080 4564 39086 4616
rect 39114 4564 39120 4616
rect 39172 4604 39178 4616
rect 39172 4576 39217 4604
rect 39172 4564 39178 4576
rect 5166 4536 5172 4548
rect 3988 4508 5172 4536
rect 5166 4496 5172 4508
rect 5224 4536 5230 4548
rect 11238 4536 11244 4548
rect 5224 4508 11244 4536
rect 5224 4496 5230 4508
rect 11238 4496 11244 4508
rect 11296 4496 11302 4548
rect 3881 4471 3939 4477
rect 3881 4437 3893 4471
rect 3927 4468 3939 4471
rect 4798 4468 4804 4480
rect 3927 4440 4804 4468
rect 3927 4437 3939 4440
rect 3881 4431 3939 4437
rect 4798 4428 4804 4440
rect 4856 4428 4862 4480
rect 39209 4471 39267 4477
rect 39209 4437 39221 4471
rect 39255 4468 39267 4471
rect 39758 4468 39764 4480
rect 39255 4440 39764 4468
rect 39255 4437 39267 4440
rect 39209 4431 39267 4437
rect 39758 4428 39764 4440
rect 39816 4428 39822 4480
rect 1104 4378 42872 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 42872 4378
rect 1104 4304 42872 4326
rect 10134 4156 10140 4208
rect 10192 4196 10198 4208
rect 18598 4196 18604 4208
rect 10192 4168 18604 4196
rect 10192 4156 10198 4168
rect 18598 4156 18604 4168
rect 18656 4156 18662 4208
rect 39758 4196 39764 4208
rect 39719 4168 39764 4196
rect 39758 4156 39764 4168
rect 39816 4156 39822 4208
rect 2133 4131 2191 4137
rect 2133 4097 2145 4131
rect 2179 4128 2191 4131
rect 2406 4128 2412 4140
rect 2179 4100 2412 4128
rect 2179 4097 2191 4100
rect 2133 4091 2191 4097
rect 2406 4088 2412 4100
rect 2464 4088 2470 4140
rect 3142 4128 3148 4140
rect 3103 4100 3148 4128
rect 3142 4088 3148 4100
rect 3200 4088 3206 4140
rect 4982 4088 4988 4140
rect 5040 4128 5046 4140
rect 5629 4131 5687 4137
rect 5040 4100 5085 4128
rect 5040 4088 5046 4100
rect 5629 4097 5641 4131
rect 5675 4128 5687 4131
rect 37826 4128 37832 4140
rect 5675 4100 12434 4128
rect 37787 4100 37832 4128
rect 5675 4097 5687 4100
rect 5629 4091 5687 4097
rect 2424 3992 2452 4088
rect 4798 4060 4804 4072
rect 4759 4032 4804 4060
rect 4798 4020 4804 4032
rect 4856 4020 4862 4072
rect 5644 3992 5672 4091
rect 7558 4020 7564 4072
rect 7616 4060 7622 4072
rect 10134 4060 10140 4072
rect 7616 4032 10140 4060
rect 7616 4020 7622 4032
rect 10134 4020 10140 4032
rect 10192 4020 10198 4072
rect 10226 4020 10232 4072
rect 10284 4060 10290 4072
rect 11422 4060 11428 4072
rect 10284 4032 11428 4060
rect 10284 4020 10290 4032
rect 11422 4020 11428 4032
rect 11480 4020 11486 4072
rect 2424 3964 5672 3992
rect 9401 3995 9459 4001
rect 9401 3961 9413 3995
rect 9447 3992 9459 3995
rect 10686 3992 10692 4004
rect 9447 3964 10692 3992
rect 9447 3961 9459 3964
rect 9401 3955 9459 3961
rect 10686 3952 10692 3964
rect 10744 3952 10750 4004
rect 12406 3992 12434 4100
rect 37826 4088 37832 4100
rect 37884 4088 37890 4140
rect 38749 4131 38807 4137
rect 38749 4097 38761 4131
rect 38795 4097 38807 4131
rect 38749 4091 38807 4097
rect 22462 4020 22468 4072
rect 22520 4060 22526 4072
rect 22649 4063 22707 4069
rect 22649 4060 22661 4063
rect 22520 4032 22661 4060
rect 22520 4020 22526 4032
rect 22649 4029 22661 4032
rect 22695 4029 22707 4063
rect 22830 4060 22836 4072
rect 22791 4032 22836 4060
rect 22649 4023 22707 4029
rect 22830 4020 22836 4032
rect 22888 4020 22894 4072
rect 23198 4060 23204 4072
rect 23159 4032 23204 4060
rect 23198 4020 23204 4032
rect 23256 4020 23262 4072
rect 38764 4060 38792 4091
rect 39022 4088 39028 4140
rect 39080 4128 39086 4140
rect 39577 4131 39635 4137
rect 39577 4128 39589 4131
rect 39080 4100 39589 4128
rect 39080 4088 39086 4100
rect 39577 4097 39589 4100
rect 39623 4097 39635 4131
rect 39577 4091 39635 4097
rect 39114 4060 39120 4072
rect 31726 4032 39120 4060
rect 31726 3992 31754 4032
rect 39114 4020 39120 4032
rect 39172 4020 39178 4072
rect 41322 4060 41328 4072
rect 41283 4032 41328 4060
rect 41322 4020 41328 4032
rect 41380 4020 41386 4072
rect 12406 3964 31754 3992
rect 2041 3927 2099 3933
rect 2041 3893 2053 3927
rect 2087 3924 2099 3927
rect 3050 3924 3056 3936
rect 2087 3896 3056 3924
rect 2087 3893 2099 3896
rect 2041 3887 2099 3893
rect 3050 3884 3056 3896
rect 3108 3884 3114 3936
rect 4890 3884 4896 3936
rect 4948 3924 4954 3936
rect 5537 3927 5595 3933
rect 5537 3924 5549 3927
rect 4948 3896 5549 3924
rect 4948 3884 4954 3896
rect 5537 3893 5549 3896
rect 5583 3893 5595 3927
rect 6362 3924 6368 3936
rect 6323 3896 6368 3924
rect 5537 3887 5595 3893
rect 6362 3884 6368 3896
rect 6420 3884 6426 3936
rect 9858 3924 9864 3936
rect 9819 3896 9864 3924
rect 9858 3884 9864 3896
rect 9916 3884 9922 3936
rect 10965 3927 11023 3933
rect 10965 3893 10977 3927
rect 11011 3924 11023 3927
rect 11330 3924 11336 3936
rect 11011 3896 11336 3924
rect 11011 3893 11023 3896
rect 10965 3887 11023 3893
rect 11330 3884 11336 3896
rect 11388 3884 11394 3936
rect 11514 3924 11520 3936
rect 11475 3896 11520 3924
rect 11514 3884 11520 3896
rect 11572 3884 11578 3936
rect 18138 3924 18144 3936
rect 18099 3896 18144 3924
rect 18138 3884 18144 3896
rect 18196 3884 18202 3936
rect 19518 3884 19524 3936
rect 19576 3924 19582 3936
rect 19613 3927 19671 3933
rect 19613 3924 19625 3927
rect 19576 3896 19625 3924
rect 19576 3884 19582 3896
rect 19613 3893 19625 3896
rect 19659 3893 19671 3927
rect 19613 3887 19671 3893
rect 21818 3884 21824 3936
rect 21876 3924 21882 3936
rect 21913 3927 21971 3933
rect 21913 3924 21925 3927
rect 21876 3896 21925 3924
rect 21876 3884 21882 3896
rect 21913 3893 21925 3896
rect 21959 3893 21971 3927
rect 34698 3924 34704 3936
rect 34659 3896 34704 3924
rect 21913 3887 21971 3893
rect 34698 3884 34704 3896
rect 34756 3884 34762 3936
rect 35618 3924 35624 3936
rect 35579 3896 35624 3924
rect 35618 3884 35624 3896
rect 35676 3884 35682 3936
rect 36725 3927 36783 3933
rect 36725 3893 36737 3927
rect 36771 3924 36783 3927
rect 37458 3924 37464 3936
rect 36771 3896 37464 3924
rect 36771 3893 36783 3896
rect 36725 3887 36783 3893
rect 37458 3884 37464 3896
rect 37516 3884 37522 3936
rect 37642 3884 37648 3936
rect 37700 3924 37706 3936
rect 37921 3927 37979 3933
rect 37921 3924 37933 3927
rect 37700 3896 37933 3924
rect 37700 3884 37706 3896
rect 37921 3893 37933 3896
rect 37967 3893 37979 3927
rect 38654 3924 38660 3936
rect 38615 3896 38660 3924
rect 37921 3887 37979 3893
rect 38654 3884 38660 3896
rect 38712 3884 38718 3936
rect 1104 3834 42872 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 42872 3834
rect 1104 3760 42872 3782
rect 8110 3680 8116 3732
rect 8168 3720 8174 3732
rect 8168 3692 12296 3720
rect 8168 3680 8174 3692
rect 9858 3652 9864 3664
rect 9048 3624 9864 3652
rect 3050 3584 3056 3596
rect 3011 3556 3056 3584
rect 3050 3544 3056 3556
rect 3108 3544 3114 3596
rect 3234 3584 3240 3596
rect 3195 3556 3240 3584
rect 3234 3544 3240 3556
rect 3292 3544 3298 3596
rect 4706 3584 4712 3596
rect 4667 3556 4712 3584
rect 4706 3544 4712 3556
rect 4764 3544 4770 3596
rect 4890 3584 4896 3596
rect 4851 3556 4896 3584
rect 4890 3544 4896 3556
rect 4948 3544 4954 3596
rect 5166 3584 5172 3596
rect 5127 3556 5172 3584
rect 5166 3544 5172 3556
rect 5224 3544 5230 3596
rect 9048 3593 9076 3624
rect 9858 3612 9864 3624
rect 9916 3612 9922 3664
rect 9033 3587 9091 3593
rect 9033 3553 9045 3587
rect 9079 3553 9091 3587
rect 9214 3584 9220 3596
rect 9175 3556 9220 3584
rect 9033 3547 9091 3553
rect 9214 3544 9220 3556
rect 9272 3544 9278 3596
rect 9674 3584 9680 3596
rect 9635 3556 9680 3584
rect 9674 3544 9680 3556
rect 9732 3544 9738 3596
rect 11330 3584 11336 3596
rect 11291 3556 11336 3584
rect 11330 3544 11336 3556
rect 11388 3544 11394 3596
rect 11698 3544 11704 3596
rect 11756 3584 11762 3596
rect 11793 3587 11851 3593
rect 11793 3584 11805 3587
rect 11756 3556 11805 3584
rect 11756 3544 11762 3556
rect 11793 3553 11805 3556
rect 11839 3553 11851 3587
rect 12268 3584 12296 3692
rect 16850 3680 16856 3732
rect 16908 3720 16914 3732
rect 22462 3720 22468 3732
rect 16908 3692 22094 3720
rect 22423 3692 22468 3720
rect 16908 3680 16914 3692
rect 22066 3652 22094 3692
rect 22462 3680 22468 3692
rect 22520 3680 22526 3732
rect 22066 3624 23612 3652
rect 16666 3584 16672 3596
rect 12268 3556 16672 3584
rect 11793 3547 11851 3553
rect 16666 3544 16672 3556
rect 16724 3544 16730 3596
rect 16850 3584 16856 3596
rect 16811 3556 16856 3584
rect 16850 3544 16856 3556
rect 16908 3544 16914 3596
rect 19518 3584 19524 3596
rect 19479 3556 19524 3584
rect 19518 3544 19524 3556
rect 19576 3544 19582 3596
rect 19978 3584 19984 3596
rect 19939 3556 19984 3584
rect 19978 3544 19984 3556
rect 20036 3544 20042 3596
rect 1394 3516 1400 3528
rect 1355 3488 1400 3516
rect 1394 3476 1400 3488
rect 1452 3476 1458 3528
rect 4246 3516 4252 3528
rect 4207 3488 4252 3516
rect 4246 3476 4252 3488
rect 4304 3476 4310 3528
rect 7190 3476 7196 3528
rect 7248 3516 7254 3528
rect 7285 3519 7343 3525
rect 7285 3516 7297 3519
rect 7248 3488 7297 3516
rect 7248 3476 7254 3488
rect 7285 3485 7297 3488
rect 7331 3485 7343 3519
rect 7285 3479 7343 3485
rect 8205 3519 8263 3525
rect 8205 3485 8217 3519
rect 8251 3485 8263 3519
rect 8205 3479 8263 3485
rect 4157 3383 4215 3389
rect 4157 3349 4169 3383
rect 4203 3380 4215 3383
rect 5350 3380 5356 3392
rect 4203 3352 5356 3380
rect 4203 3349 4215 3352
rect 4157 3343 4215 3349
rect 5350 3340 5356 3352
rect 5408 3340 5414 3392
rect 7374 3340 7380 3392
rect 7432 3380 7438 3392
rect 8113 3383 8171 3389
rect 8113 3380 8125 3383
rect 7432 3352 8125 3380
rect 7432 3340 7438 3352
rect 8113 3349 8125 3352
rect 8159 3349 8171 3383
rect 8220 3380 8248 3479
rect 14274 3476 14280 3528
rect 14332 3516 14338 3528
rect 14829 3519 14887 3525
rect 14829 3516 14841 3519
rect 14332 3488 14841 3516
rect 14332 3476 14338 3488
rect 14829 3485 14841 3488
rect 14875 3485 14887 3519
rect 14829 3479 14887 3485
rect 15657 3519 15715 3525
rect 15657 3485 15669 3519
rect 15703 3516 15715 3519
rect 16117 3519 16175 3525
rect 16117 3516 16129 3519
rect 15703 3488 16129 3516
rect 15703 3485 15715 3488
rect 15657 3479 15715 3485
rect 16117 3485 16129 3488
rect 16163 3485 16175 3519
rect 18598 3516 18604 3528
rect 18559 3488 18604 3516
rect 16117 3479 16175 3485
rect 18598 3476 18604 3488
rect 18656 3516 18662 3528
rect 23109 3519 23167 3525
rect 18656 3488 19334 3516
rect 18656 3476 18662 3488
rect 11517 3451 11575 3457
rect 11517 3417 11529 3451
rect 11563 3448 11575 3451
rect 11606 3448 11612 3460
rect 11563 3420 11612 3448
rect 11563 3417 11575 3420
rect 11517 3411 11575 3417
rect 11606 3408 11612 3420
rect 11664 3408 11670 3460
rect 16301 3451 16359 3457
rect 16301 3417 16313 3451
rect 16347 3448 16359 3451
rect 16758 3448 16764 3460
rect 16347 3420 16764 3448
rect 16347 3417 16359 3420
rect 16301 3411 16359 3417
rect 16758 3408 16764 3420
rect 16816 3408 16822 3460
rect 12158 3380 12164 3392
rect 8220 3352 12164 3380
rect 8113 3343 8171 3349
rect 12158 3340 12164 3352
rect 12216 3380 12222 3392
rect 16942 3380 16948 3392
rect 12216 3352 16948 3380
rect 12216 3340 12222 3352
rect 16942 3340 16948 3352
rect 17000 3340 17006 3392
rect 18322 3340 18328 3392
rect 18380 3380 18386 3392
rect 18509 3383 18567 3389
rect 18509 3380 18521 3383
rect 18380 3352 18521 3380
rect 18380 3340 18386 3352
rect 18509 3349 18521 3352
rect 18555 3349 18567 3383
rect 19306 3380 19334 3488
rect 23109 3485 23121 3519
rect 23155 3516 23167 3519
rect 23474 3516 23480 3528
rect 23155 3488 23480 3516
rect 23155 3485 23167 3488
rect 23109 3479 23167 3485
rect 23474 3476 23480 3488
rect 23532 3476 23538 3528
rect 23584 3525 23612 3624
rect 34698 3584 34704 3596
rect 34659 3556 34704 3584
rect 34698 3544 34704 3556
rect 34756 3544 34762 3596
rect 34882 3544 34888 3596
rect 34940 3584 34946 3596
rect 35161 3587 35219 3593
rect 35161 3584 35173 3587
rect 34940 3556 35173 3584
rect 34940 3544 34946 3556
rect 35161 3553 35173 3556
rect 35207 3553 35219 3587
rect 35161 3547 35219 3553
rect 36722 3544 36728 3596
rect 36780 3584 36786 3596
rect 37001 3587 37059 3593
rect 37001 3584 37013 3587
rect 36780 3556 37013 3584
rect 36780 3544 36786 3556
rect 37001 3553 37013 3556
rect 37047 3553 37059 3587
rect 37001 3547 37059 3553
rect 37366 3544 37372 3596
rect 37424 3584 37430 3596
rect 37461 3587 37519 3593
rect 37461 3584 37473 3587
rect 37424 3556 37473 3584
rect 37424 3544 37430 3556
rect 37461 3553 37473 3556
rect 37507 3553 37519 3587
rect 37461 3547 37519 3553
rect 41782 3544 41788 3596
rect 41840 3584 41846 3596
rect 42153 3587 42211 3593
rect 42153 3584 42165 3587
rect 41840 3556 42165 3584
rect 41840 3544 41846 3556
rect 42153 3553 42165 3556
rect 42199 3553 42211 3587
rect 42153 3547 42211 3553
rect 23569 3519 23627 3525
rect 23569 3485 23581 3519
rect 23615 3516 23627 3519
rect 27614 3516 27620 3528
rect 23615 3488 27620 3516
rect 23615 3485 23627 3488
rect 23569 3479 23627 3485
rect 27614 3476 27620 3488
rect 27672 3476 27678 3528
rect 27798 3516 27804 3528
rect 27759 3488 27804 3516
rect 27798 3476 27804 3488
rect 27856 3476 27862 3528
rect 19705 3451 19763 3457
rect 19705 3417 19717 3451
rect 19751 3448 19763 3451
rect 20530 3448 20536 3460
rect 19751 3420 20536 3448
rect 19751 3417 19763 3420
rect 19705 3411 19763 3417
rect 20530 3408 20536 3420
rect 20588 3408 20594 3460
rect 34885 3451 34943 3457
rect 22066 3420 31754 3448
rect 22066 3380 22094 3420
rect 23658 3380 23664 3392
rect 19306 3352 22094 3380
rect 23619 3352 23664 3380
rect 18509 3343 18567 3349
rect 23658 3340 23664 3352
rect 23716 3340 23722 3392
rect 31726 3380 31754 3420
rect 34885 3417 34897 3451
rect 34931 3448 34943 3451
rect 35526 3448 35532 3460
rect 34931 3420 35532 3448
rect 34931 3417 34943 3420
rect 34885 3411 34943 3417
rect 35526 3408 35532 3420
rect 35584 3408 35590 3460
rect 37182 3448 37188 3460
rect 37143 3420 37188 3448
rect 37182 3408 37188 3420
rect 37240 3408 37246 3460
rect 39758 3408 39764 3460
rect 39816 3448 39822 3460
rect 40313 3451 40371 3457
rect 40313 3448 40325 3451
rect 39816 3420 40325 3448
rect 39816 3408 39822 3420
rect 40313 3417 40325 3420
rect 40359 3417 40371 3451
rect 41966 3448 41972 3460
rect 41927 3420 41972 3448
rect 40313 3411 40371 3417
rect 41966 3408 41972 3420
rect 42024 3408 42030 3460
rect 36354 3380 36360 3392
rect 31726 3352 36360 3380
rect 36354 3340 36360 3352
rect 36412 3340 36418 3392
rect 41230 3340 41236 3392
rect 41288 3380 41294 3392
rect 42150 3380 42156 3392
rect 41288 3352 42156 3380
rect 41288 3340 41294 3352
rect 42150 3340 42156 3352
rect 42208 3340 42214 3392
rect 1104 3290 42872 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 42872 3290
rect 1104 3216 42872 3238
rect 4246 3136 4252 3188
rect 4304 3176 4310 3188
rect 9582 3176 9588 3188
rect 4304 3148 9588 3176
rect 4304 3136 4310 3148
rect 658 3068 664 3120
rect 716 3108 722 3120
rect 3697 3111 3755 3117
rect 3697 3108 3709 3111
rect 716 3080 3709 3108
rect 716 3068 722 3080
rect 3697 3077 3709 3080
rect 3743 3077 3755 3111
rect 5350 3108 5356 3120
rect 5311 3080 5356 3108
rect 3697 3071 3755 3077
rect 5350 3068 5356 3080
rect 5408 3068 5414 3120
rect 1394 3040 1400 3052
rect 1355 3012 1400 3040
rect 1394 3000 1400 3012
rect 1452 3000 1458 3052
rect 5534 3000 5540 3052
rect 5592 3040 5598 3052
rect 6380 3049 6408 3148
rect 9582 3136 9588 3148
rect 9640 3136 9646 3188
rect 12066 3136 12072 3188
rect 12124 3176 12130 3188
rect 16758 3176 16764 3188
rect 12124 3148 16620 3176
rect 16719 3148 16764 3176
rect 12124 3136 12130 3148
rect 7374 3108 7380 3120
rect 7335 3080 7380 3108
rect 7374 3068 7380 3080
rect 7432 3068 7438 3120
rect 12250 3108 12256 3120
rect 10980 3080 12256 3108
rect 6365 3043 6423 3049
rect 5592 3012 5637 3040
rect 5592 3000 5598 3012
rect 6365 3009 6377 3043
rect 6411 3009 6423 3043
rect 7190 3040 7196 3052
rect 7151 3012 7196 3040
rect 6365 3003 6423 3009
rect 7190 3000 7196 3012
rect 7248 3000 7254 3052
rect 10226 3040 10232 3052
rect 10187 3012 10232 3040
rect 10226 3000 10232 3012
rect 10284 3000 10290 3052
rect 10980 3049 11008 3080
rect 12250 3068 12256 3080
rect 12308 3068 12314 3120
rect 16592 3108 16620 3148
rect 16758 3136 16764 3148
rect 16816 3136 16822 3188
rect 16942 3136 16948 3188
rect 17000 3176 17006 3188
rect 20530 3176 20536 3188
rect 17000 3148 19334 3176
rect 20491 3148 20536 3176
rect 17000 3136 17006 3148
rect 18322 3108 18328 3120
rect 16592 3080 16896 3108
rect 18283 3080 18328 3108
rect 10965 3043 11023 3049
rect 10965 3009 10977 3043
rect 11011 3009 11023 3043
rect 11514 3040 11520 3052
rect 11475 3012 11520 3040
rect 10965 3003 11023 3009
rect 11514 3000 11520 3012
rect 11572 3000 11578 3052
rect 14274 3040 14280 3052
rect 14235 3012 14280 3040
rect 14274 3000 14280 3012
rect 14332 3000 14338 3052
rect 16868 3049 16896 3080
rect 18322 3068 18328 3080
rect 18380 3068 18386 3120
rect 19306 3108 19334 3148
rect 20530 3136 20536 3148
rect 20588 3136 20594 3188
rect 22741 3179 22799 3185
rect 22741 3145 22753 3179
rect 22787 3176 22799 3179
rect 22830 3176 22836 3188
rect 22787 3148 22836 3176
rect 22787 3145 22799 3148
rect 22741 3139 22799 3145
rect 22830 3136 22836 3148
rect 22888 3136 22894 3188
rect 23658 3108 23664 3120
rect 19306 3080 22094 3108
rect 23619 3080 23664 3108
rect 16853 3043 16911 3049
rect 16853 3009 16865 3043
rect 16899 3040 16911 3043
rect 18138 3040 18144 3052
rect 16899 3012 17080 3040
rect 18099 3012 18144 3040
rect 16899 3009 16911 3012
rect 16853 3003 16911 3009
rect 1578 2972 1584 2984
rect 1539 2944 1584 2972
rect 1578 2932 1584 2944
rect 1636 2932 1642 2984
rect 2774 2932 2780 2984
rect 2832 2972 2838 2984
rect 2832 2944 2877 2972
rect 2832 2932 2838 2944
rect 7098 2932 7104 2984
rect 7156 2972 7162 2984
rect 7653 2975 7711 2981
rect 7653 2972 7665 2975
rect 7156 2944 7665 2972
rect 7156 2932 7162 2944
rect 7653 2941 7665 2944
rect 7699 2941 7711 2975
rect 7653 2935 7711 2941
rect 10873 2975 10931 2981
rect 10873 2941 10885 2975
rect 10919 2972 10931 2975
rect 11701 2975 11759 2981
rect 11701 2972 11713 2975
rect 10919 2944 11713 2972
rect 10919 2941 10931 2944
rect 10873 2935 10931 2941
rect 11701 2941 11713 2944
rect 11747 2941 11759 2975
rect 11701 2935 11759 2941
rect 11977 2975 12035 2981
rect 11977 2941 11989 2975
rect 12023 2941 12035 2975
rect 11977 2935 12035 2941
rect 14461 2975 14519 2981
rect 14461 2941 14473 2975
rect 14507 2972 14519 2975
rect 15194 2972 15200 2984
rect 14507 2944 15200 2972
rect 14507 2941 14519 2944
rect 14461 2935 14519 2941
rect 3234 2864 3240 2916
rect 3292 2904 3298 2916
rect 9122 2904 9128 2916
rect 3292 2876 9128 2904
rect 3292 2864 3298 2876
rect 9122 2864 9128 2876
rect 9180 2864 9186 2916
rect 10962 2864 10968 2916
rect 11020 2904 11026 2916
rect 11992 2904 12020 2935
rect 15194 2932 15200 2944
rect 15252 2932 15258 2984
rect 15470 2972 15476 2984
rect 15431 2944 15476 2972
rect 15470 2932 15476 2944
rect 15528 2932 15534 2984
rect 11020 2876 12020 2904
rect 17052 2904 17080 3012
rect 18138 3000 18144 3012
rect 18196 3000 18202 3052
rect 20622 3040 20628 3052
rect 20583 3012 20628 3040
rect 20622 3000 20628 3012
rect 20680 3000 20686 3052
rect 21913 3043 21971 3049
rect 21913 3009 21925 3043
rect 21959 3009 21971 3043
rect 22066 3040 22094 3080
rect 23658 3068 23664 3080
rect 23716 3068 23722 3120
rect 35618 3108 35624 3120
rect 34900 3080 35624 3108
rect 22649 3043 22707 3049
rect 22649 3040 22661 3043
rect 22066 3012 22661 3040
rect 21913 3003 21971 3009
rect 22649 3009 22661 3012
rect 22695 3009 22707 3043
rect 23474 3040 23480 3052
rect 23435 3012 23480 3040
rect 22649 3003 22707 3009
rect 18690 2972 18696 2984
rect 18651 2944 18696 2972
rect 18690 2932 18696 2944
rect 18748 2932 18754 2984
rect 21928 2904 21956 3003
rect 23474 3000 23480 3012
rect 23532 3000 23538 3052
rect 27798 3040 27804 3052
rect 27759 3012 27804 3040
rect 27798 3000 27804 3012
rect 27856 3000 27862 3052
rect 34900 3049 34928 3080
rect 35618 3068 35624 3080
rect 35676 3068 35682 3120
rect 37737 3111 37795 3117
rect 37737 3077 37749 3111
rect 37783 3108 37795 3111
rect 38654 3108 38660 3120
rect 37783 3080 38660 3108
rect 37783 3077 37795 3080
rect 37737 3071 37795 3077
rect 38654 3068 38660 3080
rect 38712 3068 38718 3120
rect 40034 3108 40040 3120
rect 39995 3080 40040 3108
rect 40034 3068 40040 3080
rect 40092 3068 40098 3120
rect 34885 3043 34943 3049
rect 34885 3009 34897 3043
rect 34931 3009 34943 3043
rect 37550 3040 37556 3052
rect 37511 3012 37556 3040
rect 34885 3003 34943 3009
rect 37550 3000 37556 3012
rect 37608 3000 37614 3052
rect 39850 3040 39856 3052
rect 39811 3012 39856 3040
rect 39850 3000 39856 3012
rect 39908 3000 39914 3052
rect 23842 2932 23848 2984
rect 23900 2972 23906 2984
rect 23937 2975 23995 2981
rect 23937 2972 23949 2975
rect 23900 2944 23949 2972
rect 23900 2932 23906 2944
rect 23937 2941 23949 2944
rect 23983 2941 23995 2975
rect 27982 2972 27988 2984
rect 27943 2944 27988 2972
rect 23937 2935 23995 2941
rect 27982 2932 27988 2944
rect 28040 2932 28046 2984
rect 28350 2972 28356 2984
rect 28311 2944 28356 2972
rect 28350 2932 28356 2944
rect 28408 2932 28414 2984
rect 35069 2975 35127 2981
rect 35069 2941 35081 2975
rect 35115 2972 35127 2975
rect 35802 2972 35808 2984
rect 35115 2944 35808 2972
rect 35115 2941 35127 2944
rect 35069 2935 35127 2941
rect 35802 2932 35808 2944
rect 35860 2932 35866 2984
rect 36078 2972 36084 2984
rect 36039 2944 36084 2972
rect 36078 2932 36084 2944
rect 36136 2932 36142 2984
rect 39298 2972 39304 2984
rect 39259 2944 39304 2972
rect 39298 2932 39304 2944
rect 39356 2932 39362 2984
rect 40586 2972 40592 2984
rect 40547 2944 40592 2972
rect 40586 2932 40592 2944
rect 40644 2932 40650 2984
rect 17052 2876 21956 2904
rect 11020 2864 11026 2876
rect 35434 2864 35440 2916
rect 35492 2904 35498 2916
rect 38930 2904 38936 2916
rect 35492 2876 38936 2904
rect 35492 2864 35498 2876
rect 38930 2864 38936 2876
rect 38988 2864 38994 2916
rect 6457 2839 6515 2845
rect 6457 2805 6469 2839
rect 6503 2836 6515 2839
rect 6546 2836 6552 2848
rect 6503 2808 6552 2836
rect 6503 2805 6515 2808
rect 6457 2799 6515 2805
rect 6546 2796 6552 2808
rect 6604 2796 6610 2848
rect 10137 2839 10195 2845
rect 10137 2805 10149 2839
rect 10183 2836 10195 2839
rect 10778 2836 10784 2848
rect 10183 2808 10784 2836
rect 10183 2805 10195 2808
rect 10137 2799 10195 2805
rect 10778 2796 10784 2808
rect 10836 2796 10842 2848
rect 22002 2836 22008 2848
rect 21963 2808 22008 2836
rect 22002 2796 22008 2808
rect 22060 2796 22066 2848
rect 1104 2746 42872 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 42872 2746
rect 1104 2672 42872 2694
rect 1578 2592 1584 2644
rect 1636 2632 1642 2644
rect 2041 2635 2099 2641
rect 2041 2632 2053 2635
rect 1636 2604 2053 2632
rect 1636 2592 1642 2604
rect 2041 2601 2053 2604
rect 2087 2601 2099 2635
rect 2041 2595 2099 2601
rect 3418 2592 3424 2644
rect 3476 2632 3482 2644
rect 11606 2632 11612 2644
rect 3476 2604 10916 2632
rect 11567 2604 11612 2632
rect 3476 2592 3482 2604
rect 4614 2564 4620 2576
rect 3804 2536 4620 2564
rect 3804 2505 3832 2536
rect 4614 2524 4620 2536
rect 4672 2524 4678 2576
rect 6822 2524 6828 2576
rect 6880 2564 6886 2576
rect 6880 2536 9628 2564
rect 6880 2524 6886 2536
rect 3789 2499 3847 2505
rect 3789 2465 3801 2499
rect 3835 2465 3847 2499
rect 3789 2459 3847 2465
rect 3970 2456 3976 2508
rect 4028 2496 4034 2508
rect 4249 2499 4307 2505
rect 4249 2496 4261 2499
rect 4028 2468 4261 2496
rect 4028 2456 4034 2468
rect 4249 2465 4261 2468
rect 4295 2465 4307 2499
rect 6362 2496 6368 2508
rect 6323 2468 6368 2496
rect 4249 2459 4307 2465
rect 6362 2456 6368 2468
rect 6420 2456 6426 2508
rect 6546 2496 6552 2508
rect 6507 2468 6552 2496
rect 6546 2456 6552 2468
rect 6604 2456 6610 2508
rect 6730 2456 6736 2508
rect 6788 2496 6794 2508
rect 6917 2499 6975 2505
rect 6917 2496 6929 2499
rect 6788 2468 6929 2496
rect 6788 2456 6794 2468
rect 6917 2465 6929 2468
rect 6963 2465 6975 2499
rect 9122 2496 9128 2508
rect 9083 2468 9128 2496
rect 6917 2459 6975 2465
rect 9122 2456 9128 2468
rect 9180 2456 9186 2508
rect 2130 2428 2136 2440
rect 2091 2400 2136 2428
rect 2130 2388 2136 2400
rect 2188 2388 2194 2440
rect 2958 2388 2964 2440
rect 3016 2428 3022 2440
rect 3053 2431 3111 2437
rect 3053 2428 3065 2431
rect 3016 2400 3065 2428
rect 3016 2388 3022 2400
rect 3053 2397 3065 2400
rect 3099 2397 3111 2431
rect 3053 2391 3111 2397
rect 3145 2363 3203 2369
rect 3145 2329 3157 2363
rect 3191 2360 3203 2363
rect 3973 2363 4031 2369
rect 3973 2360 3985 2363
rect 3191 2332 3985 2360
rect 3191 2329 3203 2332
rect 3145 2323 3203 2329
rect 3973 2329 3985 2332
rect 4019 2329 4031 2363
rect 3973 2323 4031 2329
rect 9600 2292 9628 2536
rect 10778 2496 10784 2508
rect 10739 2468 10784 2496
rect 10778 2456 10784 2468
rect 10836 2456 10842 2508
rect 10888 2496 10916 2604
rect 11606 2592 11612 2604
rect 11664 2592 11670 2644
rect 15194 2632 15200 2644
rect 15155 2604 15200 2632
rect 15194 2592 15200 2604
rect 15252 2592 15258 2644
rect 27893 2635 27951 2641
rect 27893 2601 27905 2635
rect 27939 2632 27951 2635
rect 27982 2632 27988 2644
rect 27939 2604 27988 2632
rect 27939 2601 27951 2604
rect 27893 2595 27951 2601
rect 27982 2592 27988 2604
rect 28040 2592 28046 2644
rect 35802 2632 35808 2644
rect 35763 2604 35808 2632
rect 35802 2592 35808 2604
rect 35860 2592 35866 2644
rect 36449 2635 36507 2641
rect 36449 2601 36461 2635
rect 36495 2632 36507 2635
rect 37182 2632 37188 2644
rect 36495 2604 37188 2632
rect 36495 2601 36507 2604
rect 36449 2595 36507 2601
rect 37182 2592 37188 2604
rect 37240 2592 37246 2644
rect 41414 2564 41420 2576
rect 35912 2536 41420 2564
rect 13722 2496 13728 2508
rect 10888 2468 13728 2496
rect 13722 2456 13728 2468
rect 13780 2456 13786 2508
rect 21818 2496 21824 2508
rect 15212 2468 20760 2496
rect 21779 2468 21824 2496
rect 10965 2431 11023 2437
rect 10965 2397 10977 2431
rect 11011 2397 11023 2431
rect 10965 2391 11023 2397
rect 10686 2320 10692 2372
rect 10744 2360 10750 2372
rect 10980 2360 11008 2391
rect 11422 2388 11428 2440
rect 11480 2428 11486 2440
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 11480 2400 11713 2428
rect 11480 2388 11486 2400
rect 11701 2397 11713 2400
rect 11747 2428 11759 2431
rect 15212 2428 15240 2468
rect 11747 2400 15240 2428
rect 15289 2431 15347 2437
rect 11747 2397 11759 2400
rect 11701 2391 11759 2397
rect 15289 2397 15301 2431
rect 15335 2428 15347 2431
rect 20622 2428 20628 2440
rect 15335 2400 20628 2428
rect 15335 2397 15347 2400
rect 15289 2391 15347 2397
rect 10744 2332 11008 2360
rect 10744 2320 10750 2332
rect 15304 2292 15332 2391
rect 20622 2388 20628 2400
rect 20680 2388 20686 2440
rect 20732 2360 20760 2468
rect 21818 2456 21824 2468
rect 21876 2456 21882 2508
rect 22002 2496 22008 2508
rect 21963 2468 22008 2496
rect 22002 2456 22008 2468
rect 22060 2456 22066 2508
rect 22554 2496 22560 2508
rect 22515 2468 22560 2496
rect 22554 2456 22560 2468
rect 22612 2456 22618 2508
rect 35912 2440 35940 2536
rect 41414 2524 41420 2536
rect 41472 2524 41478 2576
rect 37458 2496 37464 2508
rect 37419 2468 37464 2496
rect 37458 2456 37464 2468
rect 37516 2456 37522 2508
rect 37642 2496 37648 2508
rect 37603 2468 37648 2496
rect 37642 2456 37648 2468
rect 37700 2456 37706 2508
rect 41322 2496 41328 2508
rect 41283 2468 41328 2496
rect 41322 2456 41328 2468
rect 41380 2456 41386 2508
rect 41693 2499 41751 2505
rect 41693 2465 41705 2499
rect 41739 2496 41751 2499
rect 42058 2496 42064 2508
rect 41739 2468 42064 2496
rect 41739 2465 41751 2468
rect 41693 2459 41751 2465
rect 42058 2456 42064 2468
rect 42116 2456 42122 2508
rect 27614 2388 27620 2440
rect 27672 2428 27678 2440
rect 27801 2431 27859 2437
rect 27801 2428 27813 2431
rect 27672 2400 27813 2428
rect 27672 2388 27678 2400
rect 27801 2397 27813 2400
rect 27847 2397 27859 2431
rect 27801 2391 27859 2397
rect 35894 2388 35900 2440
rect 35952 2428 35958 2440
rect 36354 2428 36360 2440
rect 35952 2400 36045 2428
rect 36315 2400 36360 2428
rect 35952 2388 35958 2400
rect 36354 2388 36360 2400
rect 36412 2388 36418 2440
rect 41877 2431 41935 2437
rect 41877 2397 41889 2431
rect 41923 2397 41935 2431
rect 41877 2391 41935 2397
rect 37826 2360 37832 2372
rect 20732 2332 37832 2360
rect 37826 2320 37832 2332
rect 37884 2320 37890 2372
rect 39301 2363 39359 2369
rect 39301 2329 39313 2363
rect 39347 2360 39359 2363
rect 39942 2360 39948 2372
rect 39347 2332 39948 2360
rect 39347 2329 39359 2332
rect 39301 2323 39359 2329
rect 39942 2320 39948 2332
rect 40000 2320 40006 2372
rect 41690 2320 41696 2372
rect 41748 2360 41754 2372
rect 41892 2360 41920 2391
rect 41748 2332 41920 2360
rect 41748 2320 41754 2332
rect 9600 2264 15332 2292
rect 1104 2202 42872 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 42872 2202
rect 1104 2128 42872 2150
rect 10226 2048 10232 2100
rect 10284 2088 10290 2100
rect 35894 2088 35900 2100
rect 10284 2060 35900 2088
rect 10284 2048 10290 2060
rect 35894 2048 35900 2060
rect 35952 2048 35958 2100
<< via1 >>
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 5816 41148 5868 41200
rect 7932 41191 7984 41200
rect 7932 41157 7941 41191
rect 7941 41157 7975 41191
rect 7975 41157 7984 41191
rect 7932 41148 7984 41157
rect 24492 41148 24544 41200
rect 34520 41148 34572 41200
rect 42524 41148 42576 41200
rect 1860 41123 1912 41132
rect 1860 41089 1869 41123
rect 1869 41089 1903 41123
rect 1903 41089 1912 41123
rect 1860 41080 1912 41089
rect 3700 41080 3752 41132
rect 3792 41055 3844 41064
rect 3792 41021 3801 41055
rect 3801 41021 3835 41055
rect 3835 41021 3844 41055
rect 3792 41012 3844 41021
rect 4712 41012 4764 41064
rect 12900 41055 12952 41064
rect 2688 40944 2740 40996
rect 12900 41021 12909 41055
rect 12909 41021 12943 41055
rect 12943 41021 12952 41055
rect 12900 41012 12952 41021
rect 12992 41012 13044 41064
rect 13544 41055 13596 41064
rect 13544 41021 13553 41055
rect 13553 41021 13587 41055
rect 13587 41021 13596 41055
rect 13544 41012 13596 41021
rect 21824 41055 21876 41064
rect 21824 41021 21833 41055
rect 21833 41021 21867 41055
rect 21867 41021 21876 41055
rect 21824 41012 21876 41021
rect 22008 41055 22060 41064
rect 22008 41021 22017 41055
rect 22017 41021 22051 41055
rect 22051 41021 22060 41055
rect 22008 41012 22060 41021
rect 21916 40944 21968 40996
rect 34152 40944 34204 40996
rect 41144 41012 41196 41064
rect 40132 40944 40184 40996
rect 2780 40919 2832 40928
rect 2780 40885 2789 40919
rect 2789 40885 2823 40919
rect 2823 40885 2832 40919
rect 2780 40876 2832 40885
rect 8024 40919 8076 40928
rect 8024 40885 8033 40919
rect 8033 40885 8067 40919
rect 8067 40885 8076 40919
rect 8024 40876 8076 40885
rect 10968 40919 11020 40928
rect 10968 40885 10977 40919
rect 10977 40885 11011 40919
rect 11011 40885 11020 40919
rect 10968 40876 11020 40885
rect 14096 40919 14148 40928
rect 14096 40885 14105 40919
rect 14105 40885 14139 40919
rect 14139 40885 14148 40919
rect 14096 40876 14148 40885
rect 14740 40919 14792 40928
rect 14740 40885 14749 40919
rect 14749 40885 14783 40919
rect 14783 40885 14792 40919
rect 14740 40876 14792 40885
rect 20168 40919 20220 40928
rect 20168 40885 20177 40919
rect 20177 40885 20211 40919
rect 20211 40885 20220 40919
rect 20168 40876 20220 40885
rect 24952 40919 25004 40928
rect 24952 40885 24961 40919
rect 24961 40885 24995 40919
rect 24995 40885 25004 40919
rect 24952 40876 25004 40885
rect 26700 40876 26752 40928
rect 26976 40919 27028 40928
rect 26976 40885 26985 40919
rect 26985 40885 27019 40919
rect 27019 40885 27028 40919
rect 26976 40876 27028 40885
rect 29552 40919 29604 40928
rect 29552 40885 29561 40919
rect 29561 40885 29595 40919
rect 29595 40885 29604 40919
rect 29552 40876 29604 40885
rect 32128 40876 32180 40928
rect 32312 40876 32364 40928
rect 37464 40876 37516 40928
rect 40040 40876 40092 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 21824 40672 21876 40724
rect 13360 40604 13412 40656
rect 26424 40604 26476 40656
rect 2044 40579 2096 40588
rect 2044 40545 2053 40579
rect 2053 40545 2087 40579
rect 2087 40545 2096 40579
rect 2044 40536 2096 40545
rect 4896 40536 4948 40588
rect 10968 40579 11020 40588
rect 10968 40545 10977 40579
rect 10977 40545 11011 40579
rect 11011 40545 11020 40579
rect 10968 40536 11020 40545
rect 11612 40579 11664 40588
rect 11612 40545 11621 40579
rect 11621 40545 11655 40579
rect 11655 40545 11664 40579
rect 11612 40536 11664 40545
rect 14096 40579 14148 40588
rect 14096 40545 14105 40579
rect 14105 40545 14139 40579
rect 14139 40545 14148 40579
rect 14096 40536 14148 40545
rect 14280 40536 14332 40588
rect 20168 40579 20220 40588
rect 20168 40545 20177 40579
rect 20177 40545 20211 40579
rect 20211 40545 20220 40579
rect 20168 40536 20220 40545
rect 20720 40579 20772 40588
rect 20720 40545 20729 40579
rect 20729 40545 20763 40579
rect 20763 40545 20772 40579
rect 20720 40536 20772 40545
rect 23480 40536 23532 40588
rect 26700 40579 26752 40588
rect 26700 40545 26709 40579
rect 26709 40545 26743 40579
rect 26743 40545 26752 40579
rect 26700 40536 26752 40545
rect 29552 40579 29604 40588
rect 29552 40545 29561 40579
rect 29561 40545 29595 40579
rect 29595 40545 29604 40579
rect 29552 40536 29604 40545
rect 30012 40579 30064 40588
rect 30012 40545 30021 40579
rect 30021 40545 30055 40579
rect 30055 40545 30064 40579
rect 30012 40536 30064 40545
rect 32312 40579 32364 40588
rect 32312 40545 32321 40579
rect 32321 40545 32355 40579
rect 32355 40545 32364 40579
rect 32312 40536 32364 40545
rect 32864 40579 32916 40588
rect 32864 40545 32873 40579
rect 32873 40545 32907 40579
rect 32907 40545 32916 40579
rect 32864 40536 32916 40545
rect 36084 40579 36136 40588
rect 36084 40545 36093 40579
rect 36093 40545 36127 40579
rect 36127 40545 36136 40579
rect 36084 40536 36136 40545
rect 37464 40579 37516 40588
rect 37464 40545 37473 40579
rect 37473 40545 37507 40579
rect 37507 40545 37516 40579
rect 37464 40536 37516 40545
rect 39304 40579 39356 40588
rect 39304 40545 39313 40579
rect 39313 40545 39347 40579
rect 39347 40545 39356 40579
rect 39304 40536 39356 40545
rect 41880 40579 41932 40588
rect 41880 40545 41889 40579
rect 41889 40545 41923 40579
rect 41923 40545 41932 40579
rect 41880 40536 41932 40545
rect 3240 40511 3292 40520
rect 3240 40477 3249 40511
rect 3249 40477 3283 40511
rect 3283 40477 3292 40511
rect 3240 40468 3292 40477
rect 9128 40468 9180 40520
rect 3056 40443 3108 40452
rect 3056 40409 3065 40443
rect 3065 40409 3099 40443
rect 3099 40409 3108 40443
rect 3056 40400 3108 40409
rect 5632 40400 5684 40452
rect 13176 40468 13228 40520
rect 37004 40511 37056 40520
rect 37004 40477 37013 40511
rect 37013 40477 37047 40511
rect 37047 40477 37056 40511
rect 40316 40511 40368 40520
rect 37004 40468 37056 40477
rect 40316 40477 40325 40511
rect 40325 40477 40359 40511
rect 40359 40477 40368 40511
rect 40316 40468 40368 40477
rect 14280 40443 14332 40452
rect 14280 40409 14289 40443
rect 14289 40409 14323 40443
rect 14323 40409 14332 40443
rect 14280 40400 14332 40409
rect 20352 40443 20404 40452
rect 20352 40409 20361 40443
rect 20361 40409 20395 40443
rect 20395 40409 20404 40443
rect 20352 40400 20404 40409
rect 24584 40443 24636 40452
rect 24584 40409 24593 40443
rect 24593 40409 24627 40443
rect 24627 40409 24636 40443
rect 24584 40400 24636 40409
rect 26332 40400 26384 40452
rect 29736 40443 29788 40452
rect 29736 40409 29745 40443
rect 29745 40409 29779 40443
rect 29779 40409 29788 40443
rect 29736 40400 29788 40409
rect 32496 40443 32548 40452
rect 32496 40409 32505 40443
rect 32505 40409 32539 40443
rect 32539 40409 32548 40443
rect 32496 40400 32548 40409
rect 35900 40400 35952 40452
rect 37648 40443 37700 40452
rect 37648 40409 37657 40443
rect 37657 40409 37691 40443
rect 37691 40409 37700 40443
rect 37648 40400 37700 40409
rect 40500 40443 40552 40452
rect 40500 40409 40509 40443
rect 40509 40409 40543 40443
rect 40543 40409 40552 40443
rect 40500 40400 40552 40409
rect 13176 40332 13228 40384
rect 13452 40375 13504 40384
rect 13452 40341 13461 40375
rect 13461 40341 13495 40375
rect 13495 40341 13504 40375
rect 13452 40332 13504 40341
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 3056 40128 3108 40180
rect 20352 40171 20404 40180
rect 20352 40137 20361 40171
rect 20361 40137 20395 40171
rect 20395 40137 20404 40171
rect 20352 40128 20404 40137
rect 22008 40128 22060 40180
rect 29736 40128 29788 40180
rect 37648 40128 37700 40180
rect 41328 40128 41380 40180
rect 2780 40060 2832 40112
rect 3516 40103 3568 40112
rect 3516 40069 3525 40103
rect 3525 40069 3559 40103
rect 3559 40069 3568 40103
rect 3516 40060 3568 40069
rect 3700 40060 3752 40112
rect 7196 40060 7248 40112
rect 8208 40060 8260 40112
rect 13452 40060 13504 40112
rect 4712 40035 4764 40044
rect 1584 39924 1636 39976
rect 4712 40001 4721 40035
rect 4721 40001 4755 40035
rect 4755 40001 4764 40035
rect 4712 39992 4764 40001
rect 5632 40035 5684 40044
rect 4620 39924 4672 39976
rect 5632 40001 5641 40035
rect 5641 40001 5675 40035
rect 5675 40001 5684 40035
rect 5632 39992 5684 40001
rect 6736 39992 6788 40044
rect 9128 40035 9180 40044
rect 9128 40001 9137 40035
rect 9137 40001 9171 40035
rect 9171 40001 9180 40035
rect 9128 39992 9180 40001
rect 20260 40035 20312 40044
rect 20260 40001 20269 40035
rect 20269 40001 20303 40035
rect 20303 40001 20312 40035
rect 20260 39992 20312 40001
rect 21640 39992 21692 40044
rect 25964 40035 26016 40044
rect 25964 40001 25973 40035
rect 25973 40001 26007 40035
rect 26007 40001 26016 40035
rect 25964 39992 26016 40001
rect 26332 39992 26384 40044
rect 26976 40035 27028 40044
rect 26976 40001 26985 40035
rect 26985 40001 27019 40035
rect 27019 40001 27028 40035
rect 26976 39992 27028 40001
rect 29276 40035 29328 40044
rect 29276 40001 29285 40035
rect 29285 40001 29319 40035
rect 29319 40001 29328 40035
rect 29276 39992 29328 40001
rect 31392 40035 31444 40044
rect 31392 40001 31401 40035
rect 31401 40001 31435 40035
rect 31435 40001 31444 40035
rect 31392 39992 31444 40001
rect 34796 40060 34848 40112
rect 39304 40060 39356 40112
rect 32128 40035 32180 40044
rect 32128 40001 32137 40035
rect 32137 40001 32171 40035
rect 32171 40001 32180 40035
rect 32128 39992 32180 40001
rect 38200 40035 38252 40044
rect 38200 40001 38209 40035
rect 38209 40001 38243 40035
rect 38243 40001 38252 40035
rect 38200 39992 38252 40001
rect 40040 40035 40092 40044
rect 40040 40001 40049 40035
rect 40049 40001 40083 40035
rect 40083 40001 40092 40035
rect 40040 39992 40092 40001
rect 9312 39967 9364 39976
rect 9312 39933 9321 39967
rect 9321 39933 9355 39967
rect 9355 39933 9364 39967
rect 9312 39924 9364 39933
rect 9680 39967 9732 39976
rect 9680 39933 9689 39967
rect 9689 39933 9723 39967
rect 9723 39933 9732 39967
rect 9680 39924 9732 39933
rect 12256 39967 12308 39976
rect 12256 39933 12265 39967
rect 12265 39933 12299 39967
rect 12299 39933 12308 39967
rect 12256 39924 12308 39933
rect 13268 39967 13320 39976
rect 13268 39933 13277 39967
rect 13277 39933 13311 39967
rect 13311 39933 13320 39967
rect 13268 39924 13320 39933
rect 13452 39967 13504 39976
rect 13452 39933 13461 39967
rect 13461 39933 13495 39967
rect 13495 39933 13504 39967
rect 13452 39924 13504 39933
rect 14740 39924 14792 39976
rect 15936 39967 15988 39976
rect 15936 39933 15945 39967
rect 15945 39933 15979 39967
rect 15979 39933 15988 39967
rect 15936 39924 15988 39933
rect 23296 39967 23348 39976
rect 23296 39933 23305 39967
rect 23305 39933 23339 39967
rect 23339 39933 23348 39967
rect 23296 39924 23348 39933
rect 23480 39967 23532 39976
rect 23480 39933 23489 39967
rect 23489 39933 23523 39967
rect 23523 39933 23532 39967
rect 23480 39924 23532 39933
rect 23848 39967 23900 39976
rect 23848 39933 23857 39967
rect 23857 39933 23891 39967
rect 23891 39933 23900 39967
rect 23848 39924 23900 39933
rect 27160 39967 27212 39976
rect 27160 39933 27169 39967
rect 27169 39933 27203 39967
rect 27203 39933 27212 39967
rect 27160 39924 27212 39933
rect 27344 39924 27396 39976
rect 32404 39924 32456 39976
rect 35348 39924 35400 39976
rect 41972 39924 42024 39976
rect 4988 39856 5040 39908
rect 12440 39856 12492 39908
rect 20260 39856 20312 39908
rect 6460 39788 6512 39840
rect 40316 39788 40368 39840
rect 41420 39788 41472 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 3240 39584 3292 39636
rect 9312 39627 9364 39636
rect 9312 39593 9321 39627
rect 9321 39593 9355 39627
rect 9355 39593 9364 39627
rect 9312 39584 9364 39593
rect 12992 39584 13044 39636
rect 13268 39584 13320 39636
rect 14280 39584 14332 39636
rect 23296 39584 23348 39636
rect 27160 39584 27212 39636
rect 32496 39584 32548 39636
rect 34520 39584 34572 39636
rect 34796 39627 34848 39636
rect 34796 39593 34805 39627
rect 34805 39593 34839 39627
rect 34839 39593 34848 39627
rect 34796 39584 34848 39593
rect 35900 39584 35952 39636
rect 37004 39584 37056 39636
rect 40500 39584 40552 39636
rect 41144 39584 41196 39636
rect 41972 39627 42024 39636
rect 41972 39593 41981 39627
rect 41981 39593 42015 39627
rect 42015 39593 42024 39627
rect 41972 39584 42024 39593
rect 4620 39516 4672 39568
rect 14096 39516 14148 39568
rect 15936 39516 15988 39568
rect 36728 39516 36780 39568
rect 40132 39516 40184 39568
rect 2872 39491 2924 39500
rect 2872 39457 2881 39491
rect 2881 39457 2915 39491
rect 2915 39457 2924 39491
rect 2872 39448 2924 39457
rect 5264 39491 5316 39500
rect 5264 39457 5273 39491
rect 5273 39457 5307 39491
rect 5307 39457 5316 39491
rect 5264 39448 5316 39457
rect 6460 39491 6512 39500
rect 6460 39457 6469 39491
rect 6469 39457 6503 39491
rect 6503 39457 6512 39491
rect 6460 39448 6512 39457
rect 6736 39448 6788 39500
rect 1400 39423 1452 39432
rect 1400 39389 1409 39423
rect 1409 39389 1443 39423
rect 1443 39389 1452 39423
rect 1400 39380 1452 39389
rect 9220 39423 9272 39432
rect 9220 39389 9229 39423
rect 9229 39389 9263 39423
rect 9263 39389 9272 39423
rect 9220 39380 9272 39389
rect 10232 39423 10284 39432
rect 10232 39389 10241 39423
rect 10241 39389 10275 39423
rect 10275 39389 10284 39423
rect 10232 39380 10284 39389
rect 10876 39380 10928 39432
rect 12440 39423 12492 39432
rect 12440 39389 12449 39423
rect 12449 39389 12483 39423
rect 12483 39389 12492 39423
rect 13084 39423 13136 39432
rect 12440 39380 12492 39389
rect 13084 39389 13093 39423
rect 13093 39389 13127 39423
rect 13127 39389 13136 39423
rect 14096 39423 14148 39432
rect 13084 39380 13136 39389
rect 2136 39312 2188 39364
rect 4804 39312 4856 39364
rect 8944 39312 8996 39364
rect 10416 39287 10468 39296
rect 10416 39253 10425 39287
rect 10425 39253 10459 39287
rect 10459 39253 10468 39287
rect 10416 39244 10468 39253
rect 14096 39389 14105 39423
rect 14105 39389 14139 39423
rect 14139 39389 14148 39423
rect 14096 39380 14148 39389
rect 22744 39423 22796 39432
rect 22744 39389 22753 39423
rect 22753 39389 22787 39423
rect 22787 39389 22796 39423
rect 22744 39380 22796 39389
rect 24584 39380 24636 39432
rect 26608 39423 26660 39432
rect 26608 39389 26617 39423
rect 26617 39389 26651 39423
rect 26651 39389 26660 39423
rect 26608 39380 26660 39389
rect 32864 39423 32916 39432
rect 32864 39389 32873 39423
rect 32873 39389 32907 39423
rect 32907 39389 32916 39423
rect 32864 39380 32916 39389
rect 35900 39423 35952 39432
rect 35900 39389 35909 39423
rect 35909 39389 35943 39423
rect 35943 39389 35952 39423
rect 35900 39380 35952 39389
rect 39764 39380 39816 39432
rect 41236 39380 41288 39432
rect 41420 39423 41472 39432
rect 41420 39389 41429 39423
rect 41429 39389 41463 39423
rect 41463 39389 41472 39423
rect 41420 39380 41472 39389
rect 31392 39312 31444 39364
rect 21640 39244 21692 39296
rect 29276 39244 29328 39296
rect 42248 39312 42300 39364
rect 40224 39244 40276 39296
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 2136 39083 2188 39092
rect 2136 39049 2145 39083
rect 2145 39049 2179 39083
rect 2179 39049 2188 39083
rect 2136 39040 2188 39049
rect 4804 39083 4856 39092
rect 4804 39049 4813 39083
rect 4813 39049 4847 39083
rect 4847 39049 4856 39083
rect 4804 39040 4856 39049
rect 23480 39040 23532 39092
rect 25964 39040 26016 39092
rect 39764 39040 39816 39092
rect 1584 38947 1636 38956
rect 1584 38913 1593 38947
rect 1593 38913 1627 38947
rect 1627 38913 1636 38947
rect 1584 38904 1636 38913
rect 3792 38947 3844 38956
rect 3792 38913 3801 38947
rect 3801 38913 3835 38947
rect 3835 38913 3844 38947
rect 3792 38904 3844 38913
rect 4712 38947 4764 38956
rect 4712 38913 4721 38947
rect 4721 38913 4755 38947
rect 4755 38913 4764 38947
rect 8852 38947 8904 38956
rect 4712 38904 4764 38913
rect 8852 38913 8861 38947
rect 8861 38913 8895 38947
rect 8895 38913 8904 38947
rect 9588 38947 9640 38956
rect 8852 38904 8904 38913
rect 2412 38836 2464 38888
rect 8944 38836 8996 38888
rect 9588 38913 9597 38947
rect 9597 38913 9631 38947
rect 9631 38913 9640 38947
rect 9588 38904 9640 38913
rect 14096 38972 14148 39024
rect 41236 39040 41288 39092
rect 40224 39015 40276 39024
rect 40224 38981 40233 39015
rect 40233 38981 40267 39015
rect 40267 38981 40276 39015
rect 40224 38972 40276 38981
rect 41880 39015 41932 39024
rect 41880 38981 41889 39015
rect 41889 38981 41923 39015
rect 41923 38981 41932 39015
rect 41880 38972 41932 38981
rect 10416 38904 10468 38956
rect 10876 38947 10928 38956
rect 10876 38913 10885 38947
rect 10885 38913 10919 38947
rect 10919 38913 10928 38947
rect 10876 38904 10928 38913
rect 13544 38904 13596 38956
rect 22928 38904 22980 38956
rect 32680 38947 32732 38956
rect 32680 38913 32689 38947
rect 32689 38913 32723 38947
rect 32723 38913 32732 38947
rect 32680 38904 32732 38913
rect 32864 38947 32916 38956
rect 32864 38913 32873 38947
rect 32873 38913 32907 38947
rect 32907 38913 32916 38947
rect 32864 38904 32916 38913
rect 33508 38947 33560 38956
rect 33508 38913 33517 38947
rect 33517 38913 33551 38947
rect 33551 38913 33560 38947
rect 33508 38904 33560 38913
rect 35348 38904 35400 38956
rect 36084 38904 36136 38956
rect 10324 38879 10376 38888
rect 10324 38845 10333 38879
rect 10333 38845 10367 38879
rect 10367 38845 10376 38879
rect 10324 38836 10376 38845
rect 12348 38879 12400 38888
rect 12348 38845 12357 38879
rect 12357 38845 12391 38879
rect 12391 38845 12400 38879
rect 12348 38836 12400 38845
rect 36452 38904 36504 38956
rect 38108 38947 38160 38956
rect 38108 38913 38117 38947
rect 38117 38913 38151 38947
rect 38151 38913 38160 38947
rect 38108 38904 38160 38913
rect 36912 38836 36964 38888
rect 38200 38768 38252 38820
rect 9220 38700 9272 38752
rect 11980 38700 12032 38752
rect 33324 38700 33376 38752
rect 33784 38700 33836 38752
rect 35992 38743 36044 38752
rect 35992 38709 36001 38743
rect 36001 38709 36035 38743
rect 36035 38709 36044 38743
rect 35992 38700 36044 38709
rect 38660 38700 38712 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 1400 38496 1452 38548
rect 30656 38496 30708 38548
rect 36912 38539 36964 38548
rect 36912 38505 36921 38539
rect 36921 38505 36955 38539
rect 36955 38505 36964 38539
rect 36912 38496 36964 38505
rect 32680 38428 32732 38480
rect 20260 38360 20312 38412
rect 25964 38360 26016 38412
rect 8852 38292 8904 38344
rect 10876 38335 10928 38344
rect 10876 38301 10885 38335
rect 10885 38301 10919 38335
rect 10919 38301 10928 38335
rect 10876 38292 10928 38301
rect 24952 38335 25004 38344
rect 24952 38301 24961 38335
rect 24961 38301 24995 38335
rect 24995 38301 25004 38335
rect 24952 38292 25004 38301
rect 25872 38335 25924 38344
rect 4436 38224 4488 38276
rect 25872 38301 25881 38335
rect 25881 38301 25915 38335
rect 25915 38301 25924 38335
rect 25872 38292 25924 38301
rect 26056 38335 26108 38344
rect 26056 38301 26065 38335
rect 26065 38301 26099 38335
rect 26099 38301 26108 38335
rect 26056 38292 26108 38301
rect 30196 38335 30248 38344
rect 30196 38301 30205 38335
rect 30205 38301 30239 38335
rect 30239 38301 30248 38335
rect 30196 38292 30248 38301
rect 4252 38156 4304 38208
rect 11428 38156 11480 38208
rect 25228 38224 25280 38276
rect 30288 38224 30340 38276
rect 41328 38403 41380 38412
rect 41328 38369 41337 38403
rect 41337 38369 41371 38403
rect 41371 38369 41380 38403
rect 41328 38360 41380 38369
rect 32864 38292 32916 38344
rect 33784 38335 33836 38344
rect 33784 38301 33802 38335
rect 33802 38301 33836 38335
rect 33784 38292 33836 38301
rect 34796 38292 34848 38344
rect 38660 38335 38712 38344
rect 38660 38301 38678 38335
rect 38678 38301 38712 38335
rect 38936 38335 38988 38344
rect 38660 38292 38712 38301
rect 38936 38301 38945 38335
rect 38945 38301 38979 38335
rect 38979 38301 38988 38335
rect 38936 38292 38988 38301
rect 42156 38335 42208 38344
rect 42156 38301 42165 38335
rect 42165 38301 42199 38335
rect 42199 38301 42208 38335
rect 42156 38292 42208 38301
rect 31668 38224 31720 38276
rect 22744 38156 22796 38208
rect 23388 38156 23440 38208
rect 24768 38199 24820 38208
rect 24768 38165 24777 38199
rect 24777 38165 24811 38199
rect 24811 38165 24820 38199
rect 24768 38156 24820 38165
rect 26424 38156 26476 38208
rect 30104 38156 30156 38208
rect 31208 38156 31260 38208
rect 32128 38199 32180 38208
rect 32128 38165 32137 38199
rect 32137 38165 32171 38199
rect 32171 38165 32180 38199
rect 32128 38156 32180 38165
rect 35992 38224 36044 38276
rect 41696 38224 41748 38276
rect 37556 38199 37608 38208
rect 37556 38165 37565 38199
rect 37565 38165 37599 38199
rect 37599 38165 37608 38199
rect 37556 38156 37608 38165
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 24952 37952 25004 38004
rect 30288 37952 30340 38004
rect 31208 37995 31260 38004
rect 31208 37961 31217 37995
rect 31217 37961 31251 37995
rect 31251 37961 31260 37995
rect 31208 37952 31260 37961
rect 33508 37952 33560 38004
rect 36084 37952 36136 38004
rect 38108 37995 38160 38004
rect 38108 37961 38117 37995
rect 38117 37961 38151 37995
rect 38151 37961 38160 37995
rect 38108 37952 38160 37961
rect 38844 37952 38896 38004
rect 39120 37952 39172 38004
rect 41696 37995 41748 38004
rect 41696 37961 41705 37995
rect 41705 37961 41739 37995
rect 41739 37961 41748 37995
rect 41696 37952 41748 37961
rect 4252 37927 4304 37936
rect 4252 37893 4261 37927
rect 4261 37893 4295 37927
rect 4295 37893 4304 37927
rect 4252 37884 4304 37893
rect 11980 37927 12032 37936
rect 11980 37893 11989 37927
rect 11989 37893 12023 37927
rect 12023 37893 12032 37927
rect 11980 37884 12032 37893
rect 4436 37859 4488 37868
rect 4436 37825 4445 37859
rect 4445 37825 4479 37859
rect 4479 37825 4488 37859
rect 4436 37816 4488 37825
rect 10876 37816 10928 37868
rect 17500 37859 17552 37868
rect 17500 37825 17534 37859
rect 17534 37825 17552 37859
rect 21824 37859 21876 37868
rect 17500 37816 17552 37825
rect 21824 37825 21833 37859
rect 21833 37825 21867 37859
rect 21867 37825 21876 37859
rect 21824 37816 21876 37825
rect 21916 37816 21968 37868
rect 23848 37859 23900 37868
rect 23848 37825 23857 37859
rect 23857 37825 23891 37859
rect 23891 37825 23900 37859
rect 23848 37816 23900 37825
rect 24124 37859 24176 37868
rect 24124 37825 24133 37859
rect 24133 37825 24167 37859
rect 24167 37825 24176 37859
rect 24124 37816 24176 37825
rect 26332 37884 26384 37936
rect 25136 37816 25188 37868
rect 28448 37884 28500 37936
rect 28264 37859 28316 37868
rect 28264 37825 28298 37859
rect 28298 37825 28316 37859
rect 32772 37884 32824 37936
rect 28264 37816 28316 37825
rect 30104 37859 30156 37868
rect 30104 37825 30138 37859
rect 30138 37825 30156 37859
rect 30104 37816 30156 37825
rect 32680 37816 32732 37868
rect 2780 37791 2832 37800
rect 2780 37757 2789 37791
rect 2789 37757 2823 37791
rect 2823 37757 2832 37791
rect 2780 37748 2832 37757
rect 16580 37748 16632 37800
rect 34520 37859 34572 37868
rect 34520 37825 34538 37859
rect 34538 37825 34572 37859
rect 34520 37816 34572 37825
rect 36912 37816 36964 37868
rect 37556 37816 37608 37868
rect 38660 37816 38712 37868
rect 39120 37859 39172 37868
rect 39120 37825 39129 37859
rect 39129 37825 39163 37859
rect 39163 37825 39172 37859
rect 39120 37816 39172 37825
rect 40040 37859 40092 37868
rect 40040 37825 40074 37859
rect 40074 37825 40092 37859
rect 40040 37816 40092 37825
rect 42340 37816 42392 37868
rect 34796 37791 34848 37800
rect 34796 37757 34805 37791
rect 34805 37757 34839 37791
rect 34839 37757 34848 37791
rect 34796 37748 34848 37757
rect 36452 37791 36504 37800
rect 36452 37757 36461 37791
rect 36461 37757 36495 37791
rect 36495 37757 36504 37791
rect 36452 37748 36504 37757
rect 38108 37791 38160 37800
rect 38108 37757 38117 37791
rect 38117 37757 38151 37791
rect 38151 37757 38160 37791
rect 38108 37748 38160 37757
rect 1676 37655 1728 37664
rect 1676 37621 1685 37655
rect 1685 37621 1719 37655
rect 1719 37621 1728 37655
rect 1676 37612 1728 37621
rect 17868 37612 17920 37664
rect 18328 37612 18380 37664
rect 23296 37612 23348 37664
rect 24308 37655 24360 37664
rect 24308 37621 24317 37655
rect 24317 37621 24351 37655
rect 24351 37621 24360 37655
rect 24308 37612 24360 37621
rect 25964 37612 26016 37664
rect 26608 37612 26660 37664
rect 36360 37680 36412 37732
rect 31300 37612 31352 37664
rect 32864 37612 32916 37664
rect 38752 37612 38804 37664
rect 38936 37680 38988 37732
rect 39028 37612 39080 37664
rect 39120 37612 39172 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 17500 37408 17552 37460
rect 20812 37408 20864 37460
rect 25136 37451 25188 37460
rect 25136 37417 25145 37451
rect 25145 37417 25179 37451
rect 25179 37417 25188 37451
rect 25136 37408 25188 37417
rect 29736 37408 29788 37460
rect 30196 37408 30248 37460
rect 31300 37408 31352 37460
rect 31668 37451 31720 37460
rect 31668 37417 31677 37451
rect 31677 37417 31711 37451
rect 31711 37417 31720 37451
rect 31668 37408 31720 37417
rect 33324 37451 33376 37460
rect 33324 37417 33333 37451
rect 33333 37417 33367 37451
rect 33367 37417 33376 37451
rect 33324 37408 33376 37417
rect 29920 37383 29972 37392
rect 29920 37349 29929 37383
rect 29929 37349 29963 37383
rect 29963 37349 29972 37383
rect 29920 37340 29972 37349
rect 1676 37272 1728 37324
rect 17868 37272 17920 37324
rect 24308 37272 24360 37324
rect 39304 37408 39356 37460
rect 40040 37451 40092 37460
rect 40040 37417 40049 37451
rect 40049 37417 40083 37451
rect 40083 37417 40092 37451
rect 40040 37408 40092 37417
rect 42156 37408 42208 37460
rect 38752 37383 38804 37392
rect 38752 37349 38761 37383
rect 38761 37349 38795 37383
rect 38795 37349 38804 37383
rect 38752 37340 38804 37349
rect 37556 37315 37608 37324
rect 2964 37204 3016 37256
rect 4620 37204 4672 37256
rect 14096 37204 14148 37256
rect 16580 37204 16632 37256
rect 17224 37204 17276 37256
rect 18604 37204 18656 37256
rect 20720 37204 20772 37256
rect 23204 37247 23256 37256
rect 23204 37213 23213 37247
rect 23213 37213 23247 37247
rect 23247 37213 23256 37247
rect 23204 37204 23256 37213
rect 23296 37204 23348 37256
rect 25320 37247 25372 37256
rect 25320 37213 25329 37247
rect 25329 37213 25363 37247
rect 25363 37213 25372 37247
rect 25320 37204 25372 37213
rect 25964 37204 26016 37256
rect 26332 37247 26384 37256
rect 26332 37213 26341 37247
rect 26341 37213 26375 37247
rect 26375 37213 26384 37247
rect 26332 37204 26384 37213
rect 30656 37247 30708 37256
rect 30656 37213 30665 37247
rect 30665 37213 30699 37247
rect 30699 37213 30708 37247
rect 30656 37204 30708 37213
rect 31668 37204 31720 37256
rect 2044 37136 2096 37188
rect 4896 37136 4948 37188
rect 15568 37136 15620 37188
rect 16856 37111 16908 37120
rect 16856 37077 16865 37111
rect 16865 37077 16899 37111
rect 16899 37077 16908 37111
rect 16856 37068 16908 37077
rect 18052 37111 18104 37120
rect 18052 37077 18061 37111
rect 18061 37077 18095 37111
rect 18095 37077 18104 37111
rect 18052 37068 18104 37077
rect 20536 37136 20588 37188
rect 25136 37136 25188 37188
rect 25872 37136 25924 37188
rect 19248 37111 19300 37120
rect 19248 37077 19257 37111
rect 19257 37077 19291 37111
rect 19291 37077 19300 37111
rect 19248 37068 19300 37077
rect 22468 37111 22520 37120
rect 22468 37077 22477 37111
rect 22477 37077 22511 37111
rect 22511 37077 22520 37111
rect 22468 37068 22520 37077
rect 23204 37068 23256 37120
rect 24860 37068 24912 37120
rect 26056 37068 26108 37120
rect 26608 37179 26660 37188
rect 26608 37145 26642 37179
rect 26642 37145 26660 37179
rect 29000 37179 29052 37188
rect 26608 37136 26660 37145
rect 29000 37145 29009 37179
rect 29009 37145 29043 37179
rect 29043 37145 29052 37179
rect 29000 37136 29052 37145
rect 29736 37136 29788 37188
rect 28632 37111 28684 37120
rect 28632 37077 28641 37111
rect 28641 37077 28675 37111
rect 28675 37077 28684 37111
rect 28632 37068 28684 37077
rect 28908 37068 28960 37120
rect 30288 37068 30340 37120
rect 31760 37136 31812 37188
rect 32864 37204 32916 37256
rect 32956 37247 33008 37256
rect 32956 37213 32965 37247
rect 32965 37213 32999 37247
rect 32999 37213 33008 37247
rect 32956 37204 33008 37213
rect 37556 37281 37565 37315
rect 37565 37281 37599 37315
rect 37599 37281 37608 37315
rect 37556 37272 37608 37281
rect 32220 37111 32272 37120
rect 32220 37077 32229 37111
rect 32229 37077 32263 37111
rect 32263 37077 32272 37111
rect 32220 37068 32272 37077
rect 32864 37068 32916 37120
rect 36452 37204 36504 37256
rect 36544 37136 36596 37188
rect 39212 37204 39264 37256
rect 39120 37179 39172 37188
rect 39120 37145 39129 37179
rect 39129 37145 39163 37179
rect 39163 37145 39172 37179
rect 39120 37136 39172 37145
rect 34520 37068 34572 37120
rect 35900 37111 35952 37120
rect 35900 37077 35909 37111
rect 35909 37077 35943 37111
rect 35943 37077 35952 37111
rect 35900 37068 35952 37077
rect 36636 37068 36688 37120
rect 36912 37068 36964 37120
rect 37832 37111 37884 37120
rect 37832 37077 37841 37111
rect 37841 37077 37875 37111
rect 37875 37077 37884 37111
rect 37832 37068 37884 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 2044 36907 2096 36916
rect 2044 36873 2053 36907
rect 2053 36873 2087 36907
rect 2087 36873 2096 36907
rect 2044 36864 2096 36873
rect 15568 36907 15620 36916
rect 15568 36873 15577 36907
rect 15577 36873 15611 36907
rect 15611 36873 15620 36907
rect 15568 36864 15620 36873
rect 18604 36907 18656 36916
rect 18604 36873 18613 36907
rect 18613 36873 18647 36907
rect 18647 36873 18656 36907
rect 18604 36864 18656 36873
rect 20536 36864 20588 36916
rect 21088 36907 21140 36916
rect 2228 36796 2280 36848
rect 4896 36796 4948 36848
rect 14556 36796 14608 36848
rect 21088 36873 21097 36907
rect 21097 36873 21131 36907
rect 21131 36873 21140 36907
rect 21088 36864 21140 36873
rect 23204 36907 23256 36916
rect 23204 36873 23213 36907
rect 23213 36873 23247 36907
rect 23247 36873 23256 36907
rect 23204 36864 23256 36873
rect 22468 36796 22520 36848
rect 25228 36864 25280 36916
rect 25320 36864 25372 36916
rect 28264 36907 28316 36916
rect 28264 36873 28273 36907
rect 28273 36873 28307 36907
rect 28307 36873 28316 36907
rect 28264 36864 28316 36873
rect 28908 36907 28960 36916
rect 28908 36873 28917 36907
rect 28917 36873 28951 36907
rect 28951 36873 28960 36907
rect 28908 36864 28960 36873
rect 29736 36864 29788 36916
rect 23848 36796 23900 36848
rect 30656 36864 30708 36916
rect 36544 36907 36596 36916
rect 36544 36873 36553 36907
rect 36553 36873 36587 36907
rect 36587 36873 36596 36907
rect 36544 36864 36596 36873
rect 37556 36864 37608 36916
rect 38752 36864 38804 36916
rect 4620 36728 4672 36780
rect 5540 36728 5592 36780
rect 5816 36771 5868 36780
rect 5816 36737 5825 36771
rect 5825 36737 5859 36771
rect 5859 36737 5868 36771
rect 5816 36728 5868 36737
rect 10232 36728 10284 36780
rect 4528 36660 4580 36712
rect 4988 36660 5040 36712
rect 14280 36771 14332 36780
rect 14280 36737 14289 36771
rect 14289 36737 14323 36771
rect 14323 36737 14332 36771
rect 14280 36728 14332 36737
rect 15660 36728 15712 36780
rect 15936 36728 15988 36780
rect 17500 36771 17552 36780
rect 17500 36737 17509 36771
rect 17509 36737 17543 36771
rect 17543 36737 17552 36771
rect 17500 36728 17552 36737
rect 18052 36728 18104 36780
rect 14556 36660 14608 36712
rect 17132 36660 17184 36712
rect 18144 36660 18196 36712
rect 19248 36660 19300 36712
rect 20352 36728 20404 36780
rect 20812 36728 20864 36780
rect 22100 36728 22152 36780
rect 22652 36728 22704 36780
rect 23112 36728 23164 36780
rect 25320 36728 25372 36780
rect 26884 36728 26936 36780
rect 28632 36728 28684 36780
rect 36452 36796 36504 36848
rect 36820 36796 36872 36848
rect 38844 36796 38896 36848
rect 39120 36796 39172 36848
rect 39396 36839 39448 36848
rect 23296 36660 23348 36712
rect 24124 36703 24176 36712
rect 24124 36669 24133 36703
rect 24133 36669 24167 36703
rect 24167 36669 24176 36703
rect 24124 36660 24176 36669
rect 25228 36660 25280 36712
rect 25688 36660 25740 36712
rect 30288 36728 30340 36780
rect 31208 36728 31260 36780
rect 32128 36728 32180 36780
rect 35440 36771 35492 36780
rect 35440 36737 35474 36771
rect 35474 36737 35492 36771
rect 35440 36728 35492 36737
rect 38292 36728 38344 36780
rect 39212 36728 39264 36780
rect 39396 36805 39423 36839
rect 39423 36805 39448 36839
rect 39396 36796 39448 36805
rect 41604 36771 41656 36780
rect 32956 36660 33008 36712
rect 34796 36660 34848 36712
rect 41604 36737 41613 36771
rect 41613 36737 41647 36771
rect 41647 36737 41656 36771
rect 41604 36728 41656 36737
rect 5080 36524 5132 36576
rect 14372 36567 14424 36576
rect 14372 36533 14381 36567
rect 14381 36533 14415 36567
rect 14415 36533 14424 36567
rect 14372 36524 14424 36533
rect 15752 36567 15804 36576
rect 15752 36533 15761 36567
rect 15761 36533 15795 36567
rect 15795 36533 15804 36567
rect 15752 36524 15804 36533
rect 17316 36567 17368 36576
rect 17316 36533 17325 36567
rect 17325 36533 17359 36567
rect 17359 36533 17368 36567
rect 17316 36524 17368 36533
rect 17500 36524 17552 36576
rect 18512 36524 18564 36576
rect 21732 36524 21784 36576
rect 22836 36524 22888 36576
rect 23480 36567 23532 36576
rect 23480 36533 23489 36567
rect 23489 36533 23523 36567
rect 23523 36533 23532 36567
rect 23480 36524 23532 36533
rect 25596 36524 25648 36576
rect 33784 36524 33836 36576
rect 38844 36592 38896 36644
rect 39212 36524 39264 36576
rect 41972 36524 42024 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 4896 36320 4948 36372
rect 14464 36320 14516 36372
rect 15936 36363 15988 36372
rect 15936 36329 15945 36363
rect 15945 36329 15979 36363
rect 15979 36329 15988 36363
rect 15936 36320 15988 36329
rect 16948 36363 17000 36372
rect 16948 36329 16957 36363
rect 16957 36329 16991 36363
rect 16991 36329 17000 36363
rect 16948 36320 17000 36329
rect 17224 36363 17276 36372
rect 17224 36329 17233 36363
rect 17233 36329 17267 36363
rect 17267 36329 17276 36363
rect 17224 36320 17276 36329
rect 17316 36320 17368 36372
rect 21916 36363 21968 36372
rect 4528 36252 4580 36304
rect 4988 36252 5040 36304
rect 16856 36252 16908 36304
rect 1952 36116 2004 36168
rect 2780 36023 2832 36032
rect 2780 35989 2789 36023
rect 2789 35989 2823 36023
rect 2823 35989 2832 36023
rect 2780 35980 2832 35989
rect 4620 36116 4672 36168
rect 5080 36116 5132 36168
rect 14096 36159 14148 36168
rect 14096 36125 14105 36159
rect 14105 36125 14139 36159
rect 14139 36125 14148 36159
rect 14096 36116 14148 36125
rect 14372 36159 14424 36168
rect 14372 36125 14406 36159
rect 14406 36125 14424 36159
rect 14372 36116 14424 36125
rect 15660 36116 15712 36168
rect 16212 36159 16264 36168
rect 16212 36125 16221 36159
rect 16221 36125 16255 36159
rect 16255 36125 16264 36159
rect 16212 36116 16264 36125
rect 16672 36116 16724 36168
rect 17960 36116 18012 36168
rect 21916 36329 21925 36363
rect 21925 36329 21959 36363
rect 21959 36329 21968 36363
rect 21916 36320 21968 36329
rect 23848 36320 23900 36372
rect 24768 36320 24820 36372
rect 24860 36363 24912 36372
rect 24860 36329 24869 36363
rect 24869 36329 24903 36363
rect 24903 36329 24912 36363
rect 26608 36363 26660 36372
rect 24860 36320 24912 36329
rect 26608 36329 26617 36363
rect 26617 36329 26651 36363
rect 26651 36329 26660 36363
rect 26608 36320 26660 36329
rect 35900 36363 35952 36372
rect 35900 36329 35909 36363
rect 35909 36329 35943 36363
rect 35943 36329 35952 36363
rect 35900 36320 35952 36329
rect 38844 36320 38896 36372
rect 39396 36320 39448 36372
rect 18236 36252 18288 36304
rect 33784 36252 33836 36304
rect 34520 36252 34572 36304
rect 39948 36252 40000 36304
rect 18328 36184 18380 36236
rect 21732 36184 21784 36236
rect 19248 36159 19300 36168
rect 19248 36125 19257 36159
rect 19257 36125 19291 36159
rect 19291 36125 19300 36159
rect 19248 36116 19300 36125
rect 21088 36116 21140 36168
rect 24308 36184 24360 36236
rect 25872 36184 25924 36236
rect 32956 36184 33008 36236
rect 23296 36116 23348 36168
rect 5172 36048 5224 36100
rect 13084 36048 13136 36100
rect 18512 36048 18564 36100
rect 7472 35980 7524 36032
rect 15476 36023 15528 36032
rect 15476 35989 15485 36023
rect 15485 35989 15519 36023
rect 15519 35989 15528 36023
rect 15476 35980 15528 35989
rect 16212 35980 16264 36032
rect 19432 35980 19484 36032
rect 22652 36048 22704 36100
rect 25320 36116 25372 36168
rect 25688 36159 25740 36168
rect 25688 36125 25697 36159
rect 25697 36125 25731 36159
rect 25731 36125 25740 36159
rect 25688 36116 25740 36125
rect 26056 36116 26108 36168
rect 26424 36159 26476 36168
rect 26424 36125 26433 36159
rect 26433 36125 26467 36159
rect 26467 36125 26476 36159
rect 26424 36116 26476 36125
rect 29736 36159 29788 36168
rect 29736 36125 29745 36159
rect 29745 36125 29779 36159
rect 29779 36125 29788 36159
rect 29736 36116 29788 36125
rect 30656 36159 30708 36168
rect 30656 36125 30665 36159
rect 30665 36125 30699 36159
rect 30699 36125 30708 36159
rect 30656 36116 30708 36125
rect 30748 36159 30800 36168
rect 30748 36125 30757 36159
rect 30757 36125 30791 36159
rect 30791 36125 30800 36159
rect 33140 36159 33192 36168
rect 30748 36116 30800 36125
rect 33140 36125 33149 36159
rect 33149 36125 33183 36159
rect 33183 36125 33192 36159
rect 33140 36116 33192 36125
rect 35348 36184 35400 36236
rect 36544 36159 36596 36168
rect 36544 36125 36553 36159
rect 36553 36125 36587 36159
rect 36587 36125 36596 36159
rect 36544 36116 36596 36125
rect 36636 36159 36688 36168
rect 36636 36125 36645 36159
rect 36645 36125 36679 36159
rect 36679 36125 36688 36159
rect 36636 36116 36688 36125
rect 36820 36159 36872 36168
rect 36820 36125 36829 36159
rect 36829 36125 36863 36159
rect 36863 36125 36872 36159
rect 38476 36184 38528 36236
rect 39028 36184 39080 36236
rect 41328 36227 41380 36236
rect 41328 36193 41337 36227
rect 41337 36193 41371 36227
rect 41371 36193 41380 36227
rect 41328 36184 41380 36193
rect 41972 36227 42024 36236
rect 41972 36193 41981 36227
rect 41981 36193 42015 36227
rect 42015 36193 42024 36227
rect 41972 36184 42024 36193
rect 36820 36116 36872 36125
rect 38752 36116 38804 36168
rect 39120 36159 39172 36168
rect 39120 36125 39129 36159
rect 39129 36125 39163 36159
rect 39163 36125 39172 36159
rect 39120 36116 39172 36125
rect 42156 36159 42208 36168
rect 42156 36125 42165 36159
rect 42165 36125 42199 36159
rect 42199 36125 42208 36159
rect 42156 36116 42208 36125
rect 36084 36091 36136 36100
rect 36084 36057 36093 36091
rect 36093 36057 36127 36091
rect 36127 36057 36136 36091
rect 36084 36048 36136 36057
rect 25688 36023 25740 36032
rect 25688 35989 25697 36023
rect 25697 35989 25731 36023
rect 25731 35989 25740 36023
rect 25688 35980 25740 35989
rect 29552 36023 29604 36032
rect 29552 35989 29561 36023
rect 29561 35989 29595 36023
rect 29595 35989 29604 36023
rect 29552 35980 29604 35989
rect 31760 35980 31812 36032
rect 32404 35980 32456 36032
rect 33140 35980 33192 36032
rect 35716 36023 35768 36032
rect 35716 35989 35725 36023
rect 35725 35989 35759 36023
rect 35759 35989 35768 36023
rect 35716 35980 35768 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 14280 35776 14332 35828
rect 17132 35819 17184 35828
rect 17132 35785 17141 35819
rect 17141 35785 17175 35819
rect 17175 35785 17184 35819
rect 17132 35776 17184 35785
rect 24124 35776 24176 35828
rect 25504 35776 25556 35828
rect 2780 35708 2832 35760
rect 15476 35708 15528 35760
rect 1952 35683 2004 35692
rect 1952 35649 1961 35683
rect 1961 35649 1995 35683
rect 1995 35649 2004 35683
rect 1952 35640 2004 35649
rect 5080 35683 5132 35692
rect 5080 35649 5089 35683
rect 5089 35649 5123 35683
rect 5123 35649 5132 35683
rect 5080 35640 5132 35649
rect 15292 35640 15344 35692
rect 2872 35615 2924 35624
rect 2872 35581 2881 35615
rect 2881 35581 2915 35615
rect 2915 35581 2924 35615
rect 2872 35572 2924 35581
rect 4804 35615 4856 35624
rect 4804 35581 4813 35615
rect 4813 35581 4847 35615
rect 4847 35581 4856 35615
rect 4804 35572 4856 35581
rect 15292 35504 15344 35556
rect 16672 35683 16724 35692
rect 16672 35649 16681 35683
rect 16681 35649 16715 35683
rect 16715 35649 16724 35683
rect 16672 35640 16724 35649
rect 16856 35640 16908 35692
rect 17224 35640 17276 35692
rect 17960 35572 18012 35624
rect 19616 35683 19668 35692
rect 19616 35649 19625 35683
rect 19625 35649 19659 35683
rect 19659 35649 19668 35683
rect 19616 35640 19668 35649
rect 22284 35572 22336 35624
rect 22652 35615 22704 35624
rect 22652 35581 22661 35615
rect 22661 35581 22695 35615
rect 22695 35581 22704 35615
rect 22652 35572 22704 35581
rect 23480 35640 23532 35692
rect 24952 35708 25004 35760
rect 25136 35708 25188 35760
rect 23756 35572 23808 35624
rect 20168 35504 20220 35556
rect 22560 35504 22612 35556
rect 22836 35547 22888 35556
rect 22836 35513 22845 35547
rect 22845 35513 22879 35547
rect 22879 35513 22888 35547
rect 22836 35504 22888 35513
rect 14740 35479 14792 35488
rect 14740 35445 14749 35479
rect 14749 35445 14783 35479
rect 14783 35445 14792 35479
rect 14740 35436 14792 35445
rect 18328 35436 18380 35488
rect 19064 35436 19116 35488
rect 22376 35436 22428 35488
rect 24400 35683 24452 35692
rect 24400 35649 24409 35683
rect 24409 35649 24443 35683
rect 24443 35649 24452 35683
rect 24400 35640 24452 35649
rect 24768 35640 24820 35692
rect 25228 35683 25280 35692
rect 25228 35649 25237 35683
rect 25237 35649 25271 35683
rect 25271 35649 25280 35683
rect 25228 35640 25280 35649
rect 25872 35708 25924 35760
rect 26976 35640 27028 35692
rect 29736 35776 29788 35828
rect 32128 35776 32180 35828
rect 32404 35819 32456 35828
rect 32404 35785 32413 35819
rect 32413 35785 32447 35819
rect 32447 35785 32456 35819
rect 32404 35776 32456 35785
rect 35440 35776 35492 35828
rect 29552 35708 29604 35760
rect 30840 35708 30892 35760
rect 34520 35751 34572 35760
rect 34520 35717 34538 35751
rect 34538 35717 34572 35751
rect 34520 35708 34572 35717
rect 39948 35708 40000 35760
rect 28448 35683 28500 35692
rect 28448 35649 28457 35683
rect 28457 35649 28491 35683
rect 28491 35649 28500 35683
rect 28448 35640 28500 35649
rect 32036 35640 32088 35692
rect 35716 35640 35768 35692
rect 42156 35640 42208 35692
rect 25964 35572 26016 35624
rect 26056 35572 26108 35624
rect 34796 35615 34848 35624
rect 34796 35581 34805 35615
rect 34805 35581 34839 35615
rect 34839 35581 34848 35615
rect 34796 35572 34848 35581
rect 38292 35572 38344 35624
rect 38844 35615 38896 35624
rect 38844 35581 38853 35615
rect 38853 35581 38887 35615
rect 38887 35581 38896 35615
rect 38844 35572 38896 35581
rect 38936 35572 38988 35624
rect 26608 35504 26660 35556
rect 30656 35504 30708 35556
rect 31392 35504 31444 35556
rect 32772 35504 32824 35556
rect 23940 35436 23992 35488
rect 25780 35436 25832 35488
rect 26148 35436 26200 35488
rect 30932 35436 30984 35488
rect 36084 35436 36136 35488
rect 38476 35436 38528 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 15752 35232 15804 35284
rect 19616 35232 19668 35284
rect 22744 35232 22796 35284
rect 24768 35275 24820 35284
rect 24768 35241 24777 35275
rect 24777 35241 24811 35275
rect 24811 35241 24820 35275
rect 24768 35232 24820 35241
rect 25688 35232 25740 35284
rect 16672 35164 16724 35216
rect 16948 35139 17000 35148
rect 15476 34960 15528 35012
rect 16948 35105 16957 35139
rect 16957 35105 16991 35139
rect 16991 35105 17000 35139
rect 16948 35096 17000 35105
rect 18236 35096 18288 35148
rect 18420 35139 18472 35148
rect 18420 35105 18429 35139
rect 18429 35105 18463 35139
rect 18463 35105 18472 35139
rect 18420 35096 18472 35105
rect 16672 35028 16724 35080
rect 17224 35071 17276 35080
rect 17224 35037 17233 35071
rect 17233 35037 17267 35071
rect 17267 35037 17276 35071
rect 17224 35028 17276 35037
rect 19984 35096 20036 35148
rect 21824 35139 21876 35148
rect 21824 35105 21833 35139
rect 21833 35105 21867 35139
rect 21867 35105 21876 35139
rect 21824 35096 21876 35105
rect 24952 35164 25004 35216
rect 30564 35232 30616 35284
rect 30748 35232 30800 35284
rect 31208 35232 31260 35284
rect 38016 35164 38068 35216
rect 40132 35164 40184 35216
rect 16212 34960 16264 35012
rect 19708 35071 19760 35080
rect 19708 35037 19722 35071
rect 19722 35037 19756 35071
rect 19756 35037 19760 35071
rect 19708 35028 19760 35037
rect 22652 35028 22704 35080
rect 23388 35028 23440 35080
rect 25780 35096 25832 35148
rect 24952 35071 25004 35080
rect 24952 35037 24961 35071
rect 24961 35037 24995 35071
rect 24995 35037 25004 35071
rect 24952 35028 25004 35037
rect 25596 35028 25648 35080
rect 25872 35071 25924 35080
rect 25872 35037 25881 35071
rect 25881 35037 25915 35071
rect 25915 35037 25924 35071
rect 25872 35028 25924 35037
rect 25964 35071 26016 35080
rect 25964 35037 26009 35071
rect 26009 35037 26016 35071
rect 25964 35028 26016 35037
rect 26148 35071 26200 35080
rect 26148 35037 26157 35071
rect 26157 35037 26191 35071
rect 26191 35037 26200 35071
rect 26608 35071 26660 35080
rect 26148 35028 26200 35037
rect 26608 35037 26617 35071
rect 26617 35037 26651 35071
rect 26651 35037 26660 35071
rect 26608 35028 26660 35037
rect 28448 35096 28500 35148
rect 28908 35096 28960 35148
rect 32772 35139 32824 35148
rect 32772 35105 32781 35139
rect 32781 35105 32815 35139
rect 32815 35105 32824 35139
rect 32772 35096 32824 35105
rect 34796 35096 34848 35148
rect 32036 35071 32088 35080
rect 18420 34960 18472 35012
rect 20076 34960 20128 35012
rect 22192 34960 22244 35012
rect 26424 34960 26476 35012
rect 26516 34960 26568 35012
rect 32036 35037 32045 35071
rect 32045 35037 32079 35071
rect 32079 35037 32088 35071
rect 32036 35028 32088 35037
rect 32956 35028 33008 35080
rect 35532 35071 35584 35080
rect 26884 35003 26936 35012
rect 26884 34969 26893 35003
rect 26893 34969 26927 35003
rect 26927 34969 26936 35003
rect 26884 34960 26936 34969
rect 26976 35003 27028 35012
rect 26976 34969 26985 35003
rect 26985 34969 27019 35003
rect 27019 34969 27028 35003
rect 26976 34960 27028 34969
rect 29828 35003 29880 35012
rect 29828 34969 29862 35003
rect 29862 34969 29880 35003
rect 35532 35037 35541 35071
rect 35541 35037 35575 35071
rect 35575 35037 35584 35071
rect 35532 35028 35584 35037
rect 35900 35028 35952 35080
rect 38108 35096 38160 35148
rect 38936 35096 38988 35148
rect 38752 35071 38804 35080
rect 38752 35037 38761 35071
rect 38761 35037 38795 35071
rect 38795 35037 38804 35071
rect 38752 35028 38804 35037
rect 38844 35028 38896 35080
rect 40684 35071 40736 35080
rect 29828 34960 29880 34969
rect 33140 34960 33192 35012
rect 33508 34960 33560 35012
rect 37556 34960 37608 35012
rect 40684 35037 40693 35071
rect 40693 35037 40727 35071
rect 40727 35037 40736 35071
rect 40684 35028 40736 35037
rect 41972 35071 42024 35080
rect 41972 35037 41981 35071
rect 41981 35037 42015 35071
rect 42015 35037 42024 35071
rect 41972 35028 42024 35037
rect 20260 34892 20312 34944
rect 25688 34892 25740 34944
rect 27252 34935 27304 34944
rect 27252 34901 27261 34935
rect 27261 34901 27295 34935
rect 27295 34901 27304 34935
rect 27252 34892 27304 34901
rect 31852 34935 31904 34944
rect 31852 34901 31861 34935
rect 31861 34901 31895 34935
rect 31895 34901 31904 34935
rect 31852 34892 31904 34901
rect 32496 34892 32548 34944
rect 35624 34935 35676 34944
rect 35624 34901 35633 34935
rect 35633 34901 35667 34935
rect 35667 34901 35676 34935
rect 35624 34892 35676 34901
rect 36820 34892 36872 34944
rect 37280 34892 37332 34944
rect 38108 34892 38160 34944
rect 40224 34892 40276 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 4804 34688 4856 34740
rect 17224 34688 17276 34740
rect 22192 34731 22244 34740
rect 18972 34620 19024 34672
rect 19432 34663 19484 34672
rect 14648 34552 14700 34604
rect 15476 34595 15528 34604
rect 15476 34561 15485 34595
rect 15485 34561 15519 34595
rect 15519 34561 15528 34595
rect 15476 34552 15528 34561
rect 16672 34595 16724 34604
rect 16672 34561 16681 34595
rect 16681 34561 16715 34595
rect 16715 34561 16724 34595
rect 16672 34552 16724 34561
rect 18144 34595 18196 34604
rect 18144 34561 18153 34595
rect 18153 34561 18187 34595
rect 18187 34561 18196 34595
rect 18144 34552 18196 34561
rect 18236 34595 18288 34604
rect 18236 34561 18245 34595
rect 18245 34561 18279 34595
rect 18279 34561 18288 34595
rect 18420 34595 18472 34604
rect 18236 34552 18288 34561
rect 18420 34561 18429 34595
rect 18429 34561 18463 34595
rect 18463 34561 18472 34595
rect 18420 34552 18472 34561
rect 18512 34552 18564 34604
rect 19432 34629 19438 34663
rect 19438 34629 19472 34663
rect 19472 34629 19484 34663
rect 19432 34620 19484 34629
rect 22192 34697 22201 34731
rect 22201 34697 22235 34731
rect 22235 34697 22244 34731
rect 22192 34688 22244 34697
rect 30288 34731 30340 34740
rect 30288 34697 30297 34731
rect 30297 34697 30331 34731
rect 30331 34697 30340 34731
rect 30288 34688 30340 34697
rect 30564 34688 30616 34740
rect 30840 34731 30892 34740
rect 30840 34697 30849 34731
rect 30849 34697 30883 34731
rect 30883 34697 30892 34731
rect 30840 34688 30892 34697
rect 31208 34731 31260 34740
rect 31208 34697 31217 34731
rect 31217 34697 31251 34731
rect 31251 34697 31260 34731
rect 31208 34688 31260 34697
rect 22928 34620 22980 34672
rect 25044 34620 25096 34672
rect 19340 34595 19392 34604
rect 19340 34561 19349 34595
rect 19349 34561 19383 34595
rect 19383 34561 19392 34595
rect 19340 34552 19392 34561
rect 20904 34595 20956 34604
rect 15292 34527 15344 34536
rect 15292 34493 15301 34527
rect 15301 34493 15335 34527
rect 15335 34493 15344 34527
rect 15292 34484 15344 34493
rect 14372 34391 14424 34400
rect 14372 34357 14381 34391
rect 14381 34357 14415 34391
rect 14415 34357 14424 34391
rect 14372 34348 14424 34357
rect 14740 34391 14792 34400
rect 14740 34357 14749 34391
rect 14749 34357 14783 34391
rect 14783 34357 14792 34391
rect 16580 34484 16632 34536
rect 20904 34561 20913 34595
rect 20913 34561 20947 34595
rect 20947 34561 20956 34595
rect 20904 34552 20956 34561
rect 22376 34595 22428 34604
rect 22376 34561 22385 34595
rect 22385 34561 22419 34595
rect 22419 34561 22428 34595
rect 22376 34552 22428 34561
rect 22560 34595 22612 34604
rect 22560 34561 22569 34595
rect 22569 34561 22603 34595
rect 22603 34561 22612 34595
rect 22560 34552 22612 34561
rect 22744 34552 22796 34604
rect 18144 34416 18196 34468
rect 22928 34484 22980 34536
rect 25136 34552 25188 34604
rect 27252 34620 27304 34672
rect 23756 34484 23808 34536
rect 24400 34484 24452 34536
rect 25688 34595 25740 34604
rect 25688 34561 25697 34595
rect 25697 34561 25731 34595
rect 25731 34561 25740 34595
rect 25688 34552 25740 34561
rect 26424 34552 26476 34604
rect 27528 34552 27580 34604
rect 29920 34595 29972 34604
rect 29920 34561 29929 34595
rect 29929 34561 29963 34595
rect 29963 34561 29972 34595
rect 29920 34552 29972 34561
rect 30380 34595 30432 34604
rect 30380 34561 30389 34595
rect 30389 34561 30423 34595
rect 30423 34561 30432 34595
rect 30380 34552 30432 34561
rect 30656 34552 30708 34604
rect 38016 34688 38068 34740
rect 39212 34688 39264 34740
rect 32864 34620 32916 34672
rect 32956 34620 33008 34672
rect 33508 34663 33560 34672
rect 33508 34629 33517 34663
rect 33517 34629 33551 34663
rect 33551 34629 33560 34663
rect 33508 34620 33560 34629
rect 35624 34620 35676 34672
rect 36820 34620 36872 34672
rect 38476 34663 38528 34672
rect 25412 34484 25464 34536
rect 20168 34416 20220 34468
rect 25228 34416 25280 34468
rect 32036 34416 32088 34468
rect 34520 34484 34572 34536
rect 34796 34527 34848 34536
rect 34796 34493 34805 34527
rect 34805 34493 34839 34527
rect 34839 34493 34848 34527
rect 34796 34484 34848 34493
rect 38476 34629 38485 34663
rect 38485 34629 38519 34663
rect 38519 34629 38528 34663
rect 38476 34620 38528 34629
rect 40224 34663 40276 34672
rect 40224 34629 40233 34663
rect 40233 34629 40267 34663
rect 40267 34629 40276 34663
rect 40224 34620 40276 34629
rect 41880 34663 41932 34672
rect 41880 34629 41889 34663
rect 41889 34629 41923 34663
rect 41923 34629 41932 34663
rect 41880 34620 41932 34629
rect 38384 34552 38436 34604
rect 38844 34552 38896 34604
rect 38752 34527 38804 34536
rect 38752 34493 38761 34527
rect 38761 34493 38795 34527
rect 38795 34493 38804 34527
rect 38752 34484 38804 34493
rect 40684 34484 40736 34536
rect 21088 34391 21140 34400
rect 14740 34348 14792 34357
rect 21088 34357 21097 34391
rect 21097 34357 21131 34391
rect 21131 34357 21140 34391
rect 21088 34348 21140 34357
rect 26516 34348 26568 34400
rect 30012 34348 30064 34400
rect 31852 34348 31904 34400
rect 33968 34391 34020 34400
rect 33968 34357 33977 34391
rect 33977 34357 34011 34391
rect 34011 34357 34020 34391
rect 33968 34348 34020 34357
rect 36268 34348 36320 34400
rect 38660 34391 38712 34400
rect 38660 34357 38669 34391
rect 38669 34357 38703 34391
rect 38703 34357 38712 34391
rect 38660 34348 38712 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 18512 34187 18564 34196
rect 18512 34153 18521 34187
rect 18521 34153 18555 34187
rect 18555 34153 18564 34187
rect 18512 34144 18564 34153
rect 18972 34144 19024 34196
rect 20168 34187 20220 34196
rect 20168 34153 20177 34187
rect 20177 34153 20211 34187
rect 20211 34153 20220 34187
rect 20168 34144 20220 34153
rect 27160 34187 27212 34196
rect 27160 34153 27169 34187
rect 27169 34153 27203 34187
rect 27203 34153 27212 34187
rect 27160 34144 27212 34153
rect 29828 34187 29880 34196
rect 29828 34153 29837 34187
rect 29837 34153 29871 34187
rect 29871 34153 29880 34187
rect 29828 34144 29880 34153
rect 30380 34144 30432 34196
rect 32036 34144 32088 34196
rect 35532 34144 35584 34196
rect 35900 34187 35952 34196
rect 35900 34153 35909 34187
rect 35909 34153 35943 34187
rect 35943 34153 35952 34187
rect 35900 34144 35952 34153
rect 37556 34187 37608 34196
rect 37556 34153 37565 34187
rect 37565 34153 37599 34187
rect 37599 34153 37608 34187
rect 37556 34144 37608 34153
rect 38292 34187 38344 34196
rect 38292 34153 38301 34187
rect 38301 34153 38335 34187
rect 38335 34153 38344 34187
rect 38292 34144 38344 34153
rect 15292 34076 15344 34128
rect 14096 33983 14148 33992
rect 14096 33949 14105 33983
rect 14105 33949 14139 33983
rect 14139 33949 14148 33983
rect 14096 33940 14148 33949
rect 14372 33983 14424 33992
rect 14372 33949 14406 33983
rect 14406 33949 14424 33983
rect 14372 33940 14424 33949
rect 18144 34076 18196 34128
rect 20076 34076 20128 34128
rect 20628 34076 20680 34128
rect 18328 33983 18380 33992
rect 18328 33949 18337 33983
rect 18337 33949 18371 33983
rect 18371 33949 18380 33983
rect 18328 33940 18380 33949
rect 18696 33983 18748 33992
rect 18236 33872 18288 33924
rect 18696 33949 18705 33983
rect 18705 33949 18739 33983
rect 18739 33949 18748 33983
rect 18696 33940 18748 33949
rect 19432 33940 19484 33992
rect 20076 33983 20128 33992
rect 20076 33949 20085 33983
rect 20085 33949 20119 33983
rect 20119 33949 20128 33983
rect 20076 33940 20128 33949
rect 21088 33940 21140 33992
rect 22652 33940 22704 33992
rect 26148 33940 26200 33992
rect 26516 33983 26568 33992
rect 26516 33949 26525 33983
rect 26525 33949 26559 33983
rect 26559 33949 26568 33983
rect 26516 33940 26568 33949
rect 35348 34076 35400 34128
rect 38844 34119 38896 34128
rect 30288 34051 30340 34060
rect 30288 34017 30297 34051
rect 30297 34017 30331 34051
rect 30331 34017 30340 34051
rect 30288 34008 30340 34017
rect 35624 34008 35676 34060
rect 36268 34051 36320 34060
rect 30012 33983 30064 33992
rect 30012 33949 30021 33983
rect 30021 33949 30055 33983
rect 30055 33949 30064 33983
rect 30012 33940 30064 33949
rect 33876 33940 33928 33992
rect 36268 34017 36277 34051
rect 36277 34017 36311 34051
rect 36311 34017 36320 34051
rect 36268 34008 36320 34017
rect 38844 34085 38853 34119
rect 38853 34085 38887 34119
rect 38887 34085 38896 34119
rect 38844 34076 38896 34085
rect 37188 34008 37240 34060
rect 38936 34008 38988 34060
rect 39856 34051 39908 34060
rect 39856 34017 39865 34051
rect 39865 34017 39899 34051
rect 39899 34017 39908 34051
rect 39856 34008 39908 34017
rect 36820 33983 36872 33992
rect 18788 33872 18840 33924
rect 19984 33872 20036 33924
rect 22192 33872 22244 33924
rect 28448 33872 28500 33924
rect 29000 33872 29052 33924
rect 33968 33872 34020 33924
rect 36820 33949 36829 33983
rect 36829 33949 36863 33983
rect 36863 33949 36872 33983
rect 36820 33940 36872 33949
rect 38016 33940 38068 33992
rect 38660 33983 38712 33992
rect 38660 33949 38669 33983
rect 38669 33949 38703 33983
rect 38703 33949 38712 33983
rect 38660 33940 38712 33949
rect 40132 33983 40184 33992
rect 40132 33949 40166 33983
rect 40166 33949 40184 33983
rect 40132 33940 40184 33949
rect 41604 33940 41656 33992
rect 27988 33847 28040 33856
rect 27988 33813 27997 33847
rect 27997 33813 28031 33847
rect 28031 33813 28040 33847
rect 27988 33804 28040 33813
rect 38752 33872 38804 33924
rect 38476 33847 38528 33856
rect 38476 33813 38485 33847
rect 38485 33813 38519 33847
rect 38519 33813 38528 33847
rect 38476 33804 38528 33813
rect 41696 33804 41748 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 16672 33600 16724 33652
rect 19064 33600 19116 33652
rect 19156 33575 19208 33584
rect 20904 33600 20956 33652
rect 19156 33541 19191 33575
rect 19191 33541 19208 33575
rect 19156 33532 19208 33541
rect 20628 33532 20680 33584
rect 21272 33532 21324 33584
rect 22192 33575 22244 33584
rect 22192 33541 22201 33575
rect 22201 33541 22235 33575
rect 22235 33541 22244 33575
rect 22192 33532 22244 33541
rect 16856 33507 16908 33516
rect 16856 33473 16865 33507
rect 16865 33473 16899 33507
rect 16899 33473 16908 33507
rect 16856 33464 16908 33473
rect 18880 33507 18932 33516
rect 18880 33473 18889 33507
rect 18889 33473 18923 33507
rect 18923 33473 18932 33507
rect 18880 33464 18932 33473
rect 19064 33507 19116 33516
rect 19064 33473 19073 33507
rect 19073 33473 19107 33507
rect 19107 33473 19116 33507
rect 19064 33464 19116 33473
rect 20812 33464 20864 33516
rect 19984 33396 20036 33448
rect 20536 33396 20588 33448
rect 23020 33507 23072 33516
rect 23020 33473 23029 33507
rect 23029 33473 23063 33507
rect 23063 33473 23072 33507
rect 23020 33464 23072 33473
rect 23848 33507 23900 33516
rect 23848 33473 23857 33507
rect 23857 33473 23891 33507
rect 23891 33473 23900 33507
rect 23848 33464 23900 33473
rect 25044 33464 25096 33516
rect 25136 33507 25188 33516
rect 25136 33473 25145 33507
rect 25145 33473 25179 33507
rect 25179 33473 25188 33507
rect 25964 33600 26016 33652
rect 27068 33600 27120 33652
rect 27528 33643 27580 33652
rect 27528 33609 27537 33643
rect 27537 33609 27571 33643
rect 27571 33609 27580 33643
rect 27528 33600 27580 33609
rect 27988 33532 28040 33584
rect 32036 33532 32088 33584
rect 25136 33464 25188 33473
rect 17408 33328 17460 33380
rect 19156 33328 19208 33380
rect 24860 33396 24912 33448
rect 17960 33260 18012 33312
rect 20536 33260 20588 33312
rect 26148 33396 26200 33448
rect 26516 33464 26568 33516
rect 28908 33507 28960 33516
rect 28908 33473 28917 33507
rect 28917 33473 28951 33507
rect 28951 33473 28960 33507
rect 28908 33464 28960 33473
rect 32404 33464 32456 33516
rect 35348 33532 35400 33584
rect 39028 33532 39080 33584
rect 41696 33575 41748 33584
rect 41696 33541 41705 33575
rect 41705 33541 41739 33575
rect 41739 33541 41748 33575
rect 41696 33532 41748 33541
rect 32680 33464 32732 33516
rect 38936 33464 38988 33516
rect 41972 33464 42024 33516
rect 38384 33439 38436 33448
rect 38384 33405 38393 33439
rect 38393 33405 38427 33439
rect 38427 33405 38436 33439
rect 38384 33396 38436 33405
rect 41328 33439 41380 33448
rect 41328 33405 41337 33439
rect 41337 33405 41371 33439
rect 41371 33405 41380 33439
rect 41328 33396 41380 33405
rect 33232 33328 33284 33380
rect 38476 33328 38528 33380
rect 22652 33260 22704 33312
rect 23664 33303 23716 33312
rect 23664 33269 23673 33303
rect 23673 33269 23707 33303
rect 23707 33269 23716 33303
rect 23664 33260 23716 33269
rect 24768 33303 24820 33312
rect 24768 33269 24777 33303
rect 24777 33269 24811 33303
rect 24811 33269 24820 33303
rect 24768 33260 24820 33269
rect 25688 33303 25740 33312
rect 25688 33269 25697 33303
rect 25697 33269 25731 33303
rect 25731 33269 25740 33303
rect 25688 33260 25740 33269
rect 26332 33260 26384 33312
rect 38292 33260 38344 33312
rect 39304 33260 39356 33312
rect 39948 33260 40000 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 18880 33056 18932 33108
rect 20260 32988 20312 33040
rect 18420 32920 18472 32972
rect 16856 32895 16908 32904
rect 16856 32861 16865 32895
rect 16865 32861 16899 32895
rect 16899 32861 16908 32895
rect 16856 32852 16908 32861
rect 17960 32852 18012 32904
rect 18236 32852 18288 32904
rect 18512 32895 18564 32904
rect 18512 32861 18521 32895
rect 18521 32861 18555 32895
rect 18555 32861 18564 32895
rect 18512 32852 18564 32861
rect 18788 32852 18840 32904
rect 20168 32920 20220 32972
rect 20352 32920 20404 32972
rect 20076 32895 20128 32904
rect 20076 32861 20085 32895
rect 20085 32861 20119 32895
rect 20119 32861 20128 32895
rect 20076 32852 20128 32861
rect 20812 33056 20864 33108
rect 24860 33056 24912 33108
rect 26148 33056 26200 33108
rect 27160 33056 27212 33108
rect 29920 33056 29972 33108
rect 32312 33099 32364 33108
rect 25044 32988 25096 33040
rect 30932 33031 30984 33040
rect 30932 32997 30941 33031
rect 30941 32997 30975 33031
rect 30975 32997 30984 33031
rect 30932 32988 30984 32997
rect 32312 33065 32321 33099
rect 32321 33065 32355 33099
rect 32355 33065 32364 33099
rect 32312 33056 32364 33065
rect 32956 32988 33008 33040
rect 38384 33056 38436 33108
rect 39672 33056 39724 33108
rect 39488 32988 39540 33040
rect 18328 32784 18380 32836
rect 19064 32784 19116 32836
rect 20812 32784 20864 32836
rect 22560 32852 22612 32904
rect 23664 32852 23716 32904
rect 25688 32920 25740 32972
rect 24768 32895 24820 32904
rect 24768 32861 24777 32895
rect 24777 32861 24811 32895
rect 24811 32861 24820 32895
rect 24768 32852 24820 32861
rect 24860 32895 24912 32904
rect 24860 32861 24895 32895
rect 24895 32861 24912 32895
rect 25044 32895 25096 32904
rect 24860 32852 24912 32861
rect 25044 32861 25053 32895
rect 25053 32861 25087 32895
rect 25087 32861 25096 32895
rect 25044 32852 25096 32861
rect 25412 32852 25464 32904
rect 15108 32759 15160 32768
rect 15108 32725 15117 32759
rect 15117 32725 15151 32759
rect 15151 32725 15160 32759
rect 15108 32716 15160 32725
rect 18420 32716 18472 32768
rect 18696 32716 18748 32768
rect 19984 32716 20036 32768
rect 24400 32759 24452 32768
rect 24400 32725 24409 32759
rect 24409 32725 24443 32759
rect 24443 32725 24452 32759
rect 24400 32716 24452 32725
rect 26148 32852 26200 32904
rect 27068 32895 27120 32904
rect 27068 32861 27077 32895
rect 27077 32861 27111 32895
rect 27111 32861 27120 32895
rect 27068 32852 27120 32861
rect 32220 32963 32272 32972
rect 32220 32929 32229 32963
rect 32229 32929 32263 32963
rect 32263 32929 32272 32963
rect 32220 32920 32272 32929
rect 26240 32784 26292 32836
rect 26332 32716 26384 32768
rect 29920 32895 29972 32904
rect 29920 32861 29929 32895
rect 29929 32861 29963 32895
rect 29963 32861 29972 32895
rect 29920 32852 29972 32861
rect 31208 32716 31260 32768
rect 34060 32920 34112 32972
rect 35348 32920 35400 32972
rect 37832 32920 37884 32972
rect 32496 32852 32548 32904
rect 32496 32716 32548 32768
rect 33232 32895 33284 32904
rect 33232 32861 33241 32895
rect 33241 32861 33275 32895
rect 33275 32861 33284 32895
rect 33232 32852 33284 32861
rect 34704 32895 34756 32904
rect 34704 32861 34713 32895
rect 34713 32861 34747 32895
rect 34747 32861 34756 32895
rect 34704 32852 34756 32861
rect 32956 32784 33008 32836
rect 33416 32759 33468 32768
rect 33416 32725 33425 32759
rect 33425 32725 33459 32759
rect 33459 32725 33468 32759
rect 33416 32716 33468 32725
rect 34152 32784 34204 32836
rect 35808 32852 35860 32904
rect 37004 32852 37056 32904
rect 38200 32895 38252 32904
rect 38200 32861 38209 32895
rect 38209 32861 38243 32895
rect 38243 32861 38252 32895
rect 38200 32852 38252 32861
rect 38660 32852 38712 32904
rect 40316 32895 40368 32904
rect 40316 32861 40325 32895
rect 40325 32861 40359 32895
rect 40359 32861 40368 32895
rect 40316 32852 40368 32861
rect 36360 32784 36412 32836
rect 36452 32784 36504 32836
rect 36728 32827 36780 32836
rect 36728 32793 36737 32827
rect 36737 32793 36771 32827
rect 36771 32793 36780 32827
rect 36728 32784 36780 32793
rect 37924 32784 37976 32836
rect 41512 32784 41564 32836
rect 42156 32827 42208 32836
rect 42156 32793 42165 32827
rect 42165 32793 42199 32827
rect 42199 32793 42208 32827
rect 42156 32784 42208 32793
rect 35716 32716 35768 32768
rect 36636 32759 36688 32768
rect 36636 32725 36651 32759
rect 36651 32725 36685 32759
rect 36685 32725 36688 32759
rect 36636 32716 36688 32725
rect 39120 32716 39172 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 18788 32512 18840 32564
rect 19064 32555 19116 32564
rect 19064 32521 19073 32555
rect 19073 32521 19107 32555
rect 19107 32521 19116 32555
rect 19064 32512 19116 32521
rect 21272 32512 21324 32564
rect 23848 32512 23900 32564
rect 24952 32512 25004 32564
rect 26424 32512 26476 32564
rect 26976 32512 27028 32564
rect 29920 32512 29972 32564
rect 30932 32512 30984 32564
rect 34428 32512 34480 32564
rect 34704 32512 34756 32564
rect 36452 32555 36504 32564
rect 36452 32521 36461 32555
rect 36461 32521 36495 32555
rect 36495 32521 36504 32555
rect 36452 32512 36504 32521
rect 36636 32512 36688 32564
rect 38660 32555 38712 32564
rect 14096 32376 14148 32428
rect 15108 32376 15160 32428
rect 18236 32376 18288 32428
rect 18880 32444 18932 32496
rect 19340 32376 19392 32428
rect 22560 32444 22612 32496
rect 23020 32444 23072 32496
rect 20352 32419 20404 32428
rect 20352 32385 20361 32419
rect 20361 32385 20395 32419
rect 20395 32385 20404 32419
rect 20352 32376 20404 32385
rect 24400 32444 24452 32496
rect 23940 32419 23992 32428
rect 23940 32385 23949 32419
rect 23949 32385 23983 32419
rect 23983 32385 23992 32419
rect 23940 32376 23992 32385
rect 24216 32419 24268 32428
rect 24216 32385 24225 32419
rect 24225 32385 24259 32419
rect 24259 32385 24268 32419
rect 24216 32376 24268 32385
rect 24952 32419 25004 32428
rect 24952 32385 24961 32419
rect 24961 32385 24995 32419
rect 24995 32385 25004 32419
rect 24952 32376 25004 32385
rect 27160 32419 27212 32428
rect 15844 32215 15896 32224
rect 15844 32181 15853 32215
rect 15853 32181 15887 32215
rect 15887 32181 15896 32215
rect 15844 32172 15896 32181
rect 18328 32308 18380 32360
rect 23756 32308 23808 32360
rect 24768 32308 24820 32360
rect 27160 32385 27169 32419
rect 27169 32385 27203 32419
rect 27203 32385 27212 32419
rect 27160 32376 27212 32385
rect 28632 32419 28684 32428
rect 28632 32385 28641 32419
rect 28641 32385 28675 32419
rect 28675 32385 28684 32419
rect 28632 32376 28684 32385
rect 33416 32444 33468 32496
rect 34520 32444 34572 32496
rect 38660 32521 38669 32555
rect 38669 32521 38703 32555
rect 38703 32521 38712 32555
rect 38660 32512 38712 32521
rect 39488 32555 39540 32564
rect 39488 32521 39497 32555
rect 39497 32521 39531 32555
rect 39531 32521 39540 32555
rect 39488 32512 39540 32521
rect 28908 32376 28960 32428
rect 29644 32419 29696 32428
rect 29644 32385 29678 32419
rect 29678 32385 29696 32419
rect 29644 32376 29696 32385
rect 31116 32376 31168 32428
rect 32312 32376 32364 32428
rect 32680 32419 32732 32428
rect 32680 32385 32689 32419
rect 32689 32385 32723 32419
rect 32723 32385 32732 32419
rect 32680 32376 32732 32385
rect 35716 32419 35768 32428
rect 27068 32308 27120 32360
rect 31208 32351 31260 32360
rect 31208 32317 31217 32351
rect 31217 32317 31251 32351
rect 31251 32317 31260 32351
rect 31208 32308 31260 32317
rect 31576 32308 31628 32360
rect 32864 32308 32916 32360
rect 33876 32351 33928 32360
rect 33876 32317 33885 32351
rect 33885 32317 33919 32351
rect 33919 32317 33928 32351
rect 33876 32308 33928 32317
rect 35716 32385 35725 32419
rect 35725 32385 35759 32419
rect 35759 32385 35768 32419
rect 35716 32376 35768 32385
rect 35808 32376 35860 32428
rect 36728 32419 36780 32428
rect 36728 32385 36737 32419
rect 36737 32385 36771 32419
rect 36771 32385 36780 32419
rect 36728 32376 36780 32385
rect 39120 32419 39172 32428
rect 39120 32385 39129 32419
rect 39129 32385 39163 32419
rect 39163 32385 39172 32419
rect 39120 32376 39172 32385
rect 39856 32376 39908 32428
rect 40224 32419 40276 32428
rect 40224 32385 40258 32419
rect 40258 32385 40276 32419
rect 40224 32376 40276 32385
rect 20720 32240 20772 32292
rect 30380 32240 30432 32292
rect 31392 32283 31444 32292
rect 31392 32249 31401 32283
rect 31401 32249 31435 32283
rect 31435 32249 31444 32283
rect 36360 32308 36412 32360
rect 38936 32308 38988 32360
rect 39488 32308 39540 32360
rect 31392 32240 31444 32249
rect 18512 32172 18564 32224
rect 19248 32172 19300 32224
rect 25320 32215 25372 32224
rect 25320 32181 25329 32215
rect 25329 32181 25363 32215
rect 25363 32181 25372 32215
rect 25320 32172 25372 32181
rect 25504 32172 25556 32224
rect 25872 32172 25924 32224
rect 31116 32172 31168 32224
rect 34796 32172 34848 32224
rect 37004 32172 37056 32224
rect 39212 32215 39264 32224
rect 39212 32181 39221 32215
rect 39221 32181 39255 32215
rect 39255 32181 39264 32215
rect 39212 32172 39264 32181
rect 39672 32172 39724 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 16856 31968 16908 32020
rect 18236 32011 18288 32020
rect 18236 31977 18245 32011
rect 18245 31977 18279 32011
rect 18279 31977 18288 32011
rect 18236 31968 18288 31977
rect 20076 31968 20128 32020
rect 22468 31968 22520 32020
rect 24860 31968 24912 32020
rect 27160 32011 27212 32020
rect 27160 31977 27169 32011
rect 27169 31977 27203 32011
rect 27203 31977 27212 32011
rect 27160 31968 27212 31977
rect 15568 31900 15620 31952
rect 14096 31875 14148 31884
rect 14096 31841 14105 31875
rect 14105 31841 14139 31875
rect 14139 31841 14148 31875
rect 14096 31832 14148 31841
rect 20260 31900 20312 31952
rect 20628 31900 20680 31952
rect 16212 31807 16264 31816
rect 16212 31773 16221 31807
rect 16221 31773 16255 31807
rect 16255 31773 16264 31807
rect 16212 31764 16264 31773
rect 17408 31807 17460 31816
rect 17408 31773 17417 31807
rect 17417 31773 17451 31807
rect 17451 31773 17460 31807
rect 17776 31807 17828 31816
rect 17408 31764 17460 31773
rect 17776 31773 17785 31807
rect 17785 31773 17819 31807
rect 17819 31773 17828 31807
rect 17776 31764 17828 31773
rect 18420 31807 18472 31816
rect 18420 31773 18429 31807
rect 18429 31773 18463 31807
rect 18463 31773 18472 31807
rect 18420 31764 18472 31773
rect 14372 31739 14424 31748
rect 14372 31705 14406 31739
rect 14406 31705 14424 31739
rect 14372 31696 14424 31705
rect 16948 31696 17000 31748
rect 17592 31739 17644 31748
rect 17592 31705 17601 31739
rect 17601 31705 17635 31739
rect 17635 31705 17644 31739
rect 25504 31832 25556 31884
rect 20536 31807 20588 31816
rect 20536 31773 20545 31807
rect 20545 31773 20579 31807
rect 20579 31773 20588 31807
rect 20536 31764 20588 31773
rect 20812 31764 20864 31816
rect 22652 31807 22704 31816
rect 22652 31773 22661 31807
rect 22661 31773 22695 31807
rect 22695 31773 22704 31807
rect 22652 31764 22704 31773
rect 24676 31764 24728 31816
rect 24768 31764 24820 31816
rect 25964 31764 26016 31816
rect 17592 31696 17644 31705
rect 20812 31671 20864 31680
rect 20812 31637 20821 31671
rect 20821 31637 20855 31671
rect 20855 31637 20864 31671
rect 20812 31628 20864 31637
rect 22100 31696 22152 31748
rect 26424 31807 26476 31816
rect 26424 31773 26453 31807
rect 26453 31773 26476 31807
rect 28540 31875 28592 31884
rect 28540 31841 28549 31875
rect 28549 31841 28583 31875
rect 28583 31841 28592 31875
rect 28540 31832 28592 31841
rect 28908 31832 28960 31884
rect 33876 31968 33928 32020
rect 32312 31943 32364 31952
rect 32312 31909 32321 31943
rect 32321 31909 32355 31943
rect 32355 31909 32364 31943
rect 32312 31900 32364 31909
rect 33140 31832 33192 31884
rect 34152 31832 34204 31884
rect 34796 31832 34848 31884
rect 34980 31875 35032 31884
rect 34980 31841 34989 31875
rect 34989 31841 35023 31875
rect 35023 31841 35032 31875
rect 34980 31832 35032 31841
rect 37924 31832 37976 31884
rect 38660 31875 38712 31884
rect 38660 31841 38669 31875
rect 38669 31841 38703 31875
rect 38703 31841 38712 31875
rect 38660 31832 38712 31841
rect 41328 31875 41380 31884
rect 41328 31841 41337 31875
rect 41337 31841 41371 31875
rect 41371 31841 41380 31875
rect 41328 31832 41380 31841
rect 26424 31764 26476 31773
rect 31116 31807 31168 31816
rect 26976 31696 27028 31748
rect 31116 31773 31125 31807
rect 31125 31773 31159 31807
rect 31159 31773 31168 31807
rect 31116 31764 31168 31773
rect 31668 31807 31720 31816
rect 31668 31773 31677 31807
rect 31677 31773 31711 31807
rect 31711 31773 31720 31807
rect 31668 31764 31720 31773
rect 33324 31807 33376 31816
rect 33324 31773 33333 31807
rect 33333 31773 33367 31807
rect 33367 31773 33376 31807
rect 33324 31764 33376 31773
rect 37004 31807 37056 31816
rect 37004 31773 37013 31807
rect 37013 31773 37047 31807
rect 37047 31773 37056 31807
rect 37004 31764 37056 31773
rect 37280 31807 37332 31816
rect 37280 31773 37289 31807
rect 37289 31773 37323 31807
rect 37323 31773 37332 31807
rect 37280 31764 37332 31773
rect 42156 31807 42208 31816
rect 42156 31773 42165 31807
rect 42165 31773 42199 31807
rect 42199 31773 42208 31807
rect 42156 31764 42208 31773
rect 31300 31696 31352 31748
rect 31392 31696 31444 31748
rect 41972 31739 42024 31748
rect 41972 31705 41981 31739
rect 41981 31705 42015 31739
rect 42015 31705 42024 31739
rect 41972 31696 42024 31705
rect 22008 31628 22060 31680
rect 25964 31628 26016 31680
rect 29184 31628 29236 31680
rect 30840 31628 30892 31680
rect 32312 31628 32364 31680
rect 32404 31628 32456 31680
rect 33232 31628 33284 31680
rect 33324 31628 33376 31680
rect 34428 31628 34480 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 14372 31424 14424 31476
rect 15936 31467 15988 31476
rect 15936 31433 15945 31467
rect 15945 31433 15979 31467
rect 15979 31433 15988 31467
rect 15936 31424 15988 31433
rect 17776 31424 17828 31476
rect 22100 31424 22152 31476
rect 25044 31424 25096 31476
rect 25964 31424 26016 31476
rect 26240 31424 26292 31476
rect 26976 31467 27028 31476
rect 26976 31433 26985 31467
rect 26985 31433 27019 31467
rect 27019 31433 27028 31467
rect 26976 31424 27028 31433
rect 29644 31424 29696 31476
rect 15200 31356 15252 31408
rect 15568 31399 15620 31408
rect 15568 31365 15577 31399
rect 15577 31365 15611 31399
rect 15611 31365 15620 31399
rect 15568 31356 15620 31365
rect 19984 31356 20036 31408
rect 14372 31220 14424 31272
rect 14740 31331 14792 31340
rect 14740 31297 14749 31331
rect 14749 31297 14783 31331
rect 14783 31297 14792 31331
rect 14740 31288 14792 31297
rect 15844 31288 15896 31340
rect 16948 31331 17000 31340
rect 16948 31297 16957 31331
rect 16957 31297 16991 31331
rect 16991 31297 17000 31331
rect 16948 31288 17000 31297
rect 20352 31288 20404 31340
rect 20812 31331 20864 31340
rect 20812 31297 20821 31331
rect 20821 31297 20855 31331
rect 20855 31297 20864 31331
rect 20812 31288 20864 31297
rect 22008 31331 22060 31340
rect 16488 31220 16540 31272
rect 22008 31297 22017 31331
rect 22017 31297 22051 31331
rect 22051 31297 22060 31331
rect 22008 31288 22060 31297
rect 21364 31220 21416 31272
rect 21548 31220 21600 31272
rect 25688 31356 25740 31408
rect 23388 31331 23440 31340
rect 23388 31297 23397 31331
rect 23397 31297 23431 31331
rect 23431 31297 23440 31331
rect 23388 31288 23440 31297
rect 23572 31331 23624 31340
rect 23572 31297 23581 31331
rect 23581 31297 23615 31331
rect 23615 31297 23624 31331
rect 23572 31288 23624 31297
rect 24216 31288 24268 31340
rect 24768 31288 24820 31340
rect 25872 31288 25924 31340
rect 27344 31356 27396 31408
rect 28448 31399 28500 31408
rect 28448 31365 28457 31399
rect 28457 31365 28491 31399
rect 28491 31365 28500 31399
rect 28448 31356 28500 31365
rect 29000 31288 29052 31340
rect 30380 31356 30432 31408
rect 30840 31424 30892 31476
rect 32312 31467 32364 31476
rect 32312 31433 32337 31467
rect 32337 31433 32364 31467
rect 34060 31467 34112 31476
rect 32312 31424 32364 31433
rect 34060 31433 34069 31467
rect 34069 31433 34103 31467
rect 34103 31433 34112 31467
rect 34060 31424 34112 31433
rect 34428 31424 34480 31476
rect 38292 31467 38344 31476
rect 38292 31433 38301 31467
rect 38301 31433 38335 31467
rect 38335 31433 38344 31467
rect 38292 31424 38344 31433
rect 38476 31467 38528 31476
rect 38476 31433 38485 31467
rect 38485 31433 38519 31467
rect 38519 31433 38528 31467
rect 38476 31424 38528 31433
rect 39028 31424 39080 31476
rect 39488 31467 39540 31476
rect 39488 31433 39497 31467
rect 39497 31433 39531 31467
rect 39531 31433 39540 31467
rect 39488 31424 39540 31433
rect 40224 31467 40276 31476
rect 40224 31433 40233 31467
rect 40233 31433 40267 31467
rect 40267 31433 40276 31467
rect 40224 31424 40276 31433
rect 41512 31467 41564 31476
rect 41512 31433 41521 31467
rect 41521 31433 41555 31467
rect 41555 31433 41564 31467
rect 41512 31424 41564 31433
rect 26332 31220 26384 31272
rect 27160 31263 27212 31272
rect 27160 31229 27169 31263
rect 27169 31229 27203 31263
rect 27203 31229 27212 31263
rect 27160 31220 27212 31229
rect 10324 31152 10376 31204
rect 26884 31152 26936 31204
rect 20352 31084 20404 31136
rect 23296 31084 23348 31136
rect 24860 31084 24912 31136
rect 25872 31084 25924 31136
rect 25964 31084 26016 31136
rect 30840 31288 30892 31340
rect 31576 31220 31628 31272
rect 30840 31084 30892 31136
rect 32220 31356 32272 31408
rect 33140 31356 33192 31408
rect 34520 31356 34572 31408
rect 35532 31399 35584 31408
rect 32772 31152 32824 31204
rect 34428 31288 34480 31340
rect 35532 31365 35541 31399
rect 35541 31365 35575 31399
rect 35575 31365 35584 31399
rect 35532 31356 35584 31365
rect 37280 31356 37332 31408
rect 35440 31331 35492 31340
rect 35440 31297 35449 31331
rect 35449 31297 35483 31331
rect 35483 31297 35492 31331
rect 35440 31288 35492 31297
rect 37924 31331 37976 31340
rect 37924 31297 37933 31331
rect 37933 31297 37967 31331
rect 37967 31297 37976 31331
rect 37924 31288 37976 31297
rect 38292 31288 38344 31340
rect 39672 31356 39724 31408
rect 39580 31331 39632 31340
rect 39580 31297 39589 31331
rect 39589 31297 39623 31331
rect 39623 31297 39632 31331
rect 39580 31288 39632 31297
rect 39948 31288 40000 31340
rect 40316 31288 40368 31340
rect 41420 31331 41472 31340
rect 41420 31297 41429 31331
rect 41429 31297 41463 31331
rect 41463 31297 41472 31331
rect 41420 31288 41472 31297
rect 34796 31152 34848 31204
rect 34980 31152 35032 31204
rect 32404 31084 32456 31136
rect 34336 31127 34388 31136
rect 34336 31093 34345 31127
rect 34345 31093 34379 31127
rect 34379 31093 34388 31127
rect 34336 31084 34388 31093
rect 34704 31084 34756 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 14740 30880 14792 30932
rect 15200 30880 15252 30932
rect 16212 30880 16264 30932
rect 17592 30923 17644 30932
rect 17592 30889 17601 30923
rect 17601 30889 17635 30923
rect 17635 30889 17644 30923
rect 17592 30880 17644 30889
rect 21364 30923 21416 30932
rect 21364 30889 21373 30923
rect 21373 30889 21407 30923
rect 21407 30889 21416 30923
rect 21364 30880 21416 30889
rect 22560 30923 22612 30932
rect 22560 30889 22569 30923
rect 22569 30889 22603 30923
rect 22603 30889 22612 30923
rect 22560 30880 22612 30889
rect 23296 30880 23348 30932
rect 25044 30880 25096 30932
rect 25780 30923 25832 30932
rect 25780 30889 25789 30923
rect 25789 30889 25823 30923
rect 25823 30889 25832 30923
rect 25780 30880 25832 30889
rect 26884 30880 26936 30932
rect 13728 30608 13780 30660
rect 14372 30719 14424 30728
rect 14372 30685 14381 30719
rect 14381 30685 14415 30719
rect 14415 30685 14424 30719
rect 14372 30676 14424 30685
rect 16580 30812 16632 30864
rect 20996 30812 21048 30864
rect 19248 30744 19300 30796
rect 20812 30744 20864 30796
rect 15660 30608 15712 30660
rect 14188 30540 14240 30592
rect 16212 30676 16264 30728
rect 16488 30719 16540 30728
rect 16488 30685 16503 30719
rect 16503 30685 16537 30719
rect 16537 30685 16540 30719
rect 16672 30719 16724 30728
rect 16488 30676 16540 30685
rect 16672 30685 16681 30719
rect 16681 30685 16715 30719
rect 16715 30685 16724 30719
rect 16672 30676 16724 30685
rect 17224 30676 17276 30728
rect 17776 30719 17828 30728
rect 17776 30685 17785 30719
rect 17785 30685 17819 30719
rect 17819 30685 17828 30719
rect 17776 30676 17828 30685
rect 20628 30719 20680 30728
rect 20628 30685 20637 30719
rect 20637 30685 20671 30719
rect 20671 30685 20680 30719
rect 20628 30676 20680 30685
rect 20996 30676 21048 30728
rect 21548 30719 21600 30728
rect 21548 30685 21557 30719
rect 21557 30685 21591 30719
rect 21591 30685 21600 30719
rect 21548 30676 21600 30685
rect 23572 30676 23624 30728
rect 25136 30812 25188 30864
rect 29000 30812 29052 30864
rect 32404 30880 32456 30932
rect 32772 30923 32824 30932
rect 32772 30889 32781 30923
rect 32781 30889 32815 30923
rect 32815 30889 32824 30923
rect 32772 30880 32824 30889
rect 34336 30880 34388 30932
rect 34796 30812 34848 30864
rect 35348 30880 35400 30932
rect 38568 30923 38620 30932
rect 38568 30889 38577 30923
rect 38577 30889 38611 30923
rect 38611 30889 38620 30923
rect 38568 30880 38620 30889
rect 39120 30880 39172 30932
rect 39580 30880 39632 30932
rect 41972 30880 42024 30932
rect 28540 30744 28592 30796
rect 35164 30812 35216 30864
rect 24886 30719 24938 30728
rect 24886 30685 24908 30719
rect 24908 30685 24938 30719
rect 22652 30651 22704 30660
rect 22652 30617 22661 30651
rect 22661 30617 22695 30651
rect 22695 30617 22704 30651
rect 22652 30608 22704 30617
rect 24886 30676 24938 30685
rect 25044 30719 25096 30728
rect 25044 30685 25053 30719
rect 25053 30685 25087 30719
rect 25087 30685 25096 30719
rect 25044 30676 25096 30685
rect 27068 30676 27120 30728
rect 30380 30676 30432 30728
rect 30840 30676 30892 30728
rect 31576 30676 31628 30728
rect 33232 30676 33284 30728
rect 33968 30676 34020 30728
rect 34428 30676 34480 30728
rect 26240 30608 26292 30660
rect 15844 30540 15896 30592
rect 16948 30540 17000 30592
rect 18236 30540 18288 30592
rect 20536 30540 20588 30592
rect 24400 30583 24452 30592
rect 24400 30549 24409 30583
rect 24409 30549 24443 30583
rect 24443 30549 24452 30583
rect 24400 30540 24452 30549
rect 28448 30608 28500 30660
rect 28632 30651 28684 30660
rect 28632 30617 28641 30651
rect 28641 30617 28675 30651
rect 28675 30617 28684 30651
rect 28632 30608 28684 30617
rect 33416 30608 33468 30660
rect 34704 30651 34756 30660
rect 34704 30617 34713 30651
rect 34713 30617 34747 30651
rect 34747 30617 34756 30651
rect 34704 30608 34756 30617
rect 35440 30744 35492 30796
rect 35624 30744 35676 30796
rect 35532 30719 35584 30728
rect 35532 30685 35541 30719
rect 35541 30685 35575 30719
rect 35575 30685 35584 30719
rect 35532 30676 35584 30685
rect 37004 30676 37056 30728
rect 37924 30744 37976 30796
rect 38292 30676 38344 30728
rect 41880 30676 41932 30728
rect 32680 30540 32732 30592
rect 34152 30540 34204 30592
rect 36452 30540 36504 30592
rect 37924 30583 37976 30592
rect 37924 30549 37933 30583
rect 37933 30549 37967 30583
rect 37967 30549 37976 30583
rect 37924 30540 37976 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 14004 30336 14056 30388
rect 14372 30336 14424 30388
rect 16672 30379 16724 30388
rect 16672 30345 16681 30379
rect 16681 30345 16715 30379
rect 16715 30345 16724 30379
rect 16672 30336 16724 30345
rect 13728 30132 13780 30184
rect 14004 30243 14056 30252
rect 14004 30209 14013 30243
rect 14013 30209 14047 30243
rect 14047 30209 14056 30243
rect 14188 30243 14240 30252
rect 14004 30200 14056 30209
rect 14188 30209 14197 30243
rect 14197 30209 14231 30243
rect 14231 30209 14240 30243
rect 14188 30200 14240 30209
rect 14924 30268 14976 30320
rect 14464 30200 14516 30252
rect 14556 30243 14608 30252
rect 14556 30209 14565 30243
rect 14565 30209 14599 30243
rect 14599 30209 14608 30243
rect 14556 30200 14608 30209
rect 14832 30200 14884 30252
rect 21364 30336 21416 30388
rect 23572 30336 23624 30388
rect 25504 30379 25556 30388
rect 25504 30345 25513 30379
rect 25513 30345 25547 30379
rect 25547 30345 25556 30379
rect 25504 30336 25556 30345
rect 26240 30336 26292 30388
rect 15752 30132 15804 30184
rect 11980 30064 12032 30116
rect 17224 30175 17276 30184
rect 17224 30141 17233 30175
rect 17233 30141 17267 30175
rect 17267 30141 17276 30175
rect 17224 30132 17276 30141
rect 18512 30200 18564 30252
rect 19800 30200 19852 30252
rect 21548 30268 21600 30320
rect 24400 30311 24452 30320
rect 24400 30277 24418 30311
rect 24418 30277 24452 30311
rect 24400 30268 24452 30277
rect 25780 30268 25832 30320
rect 22192 30200 22244 30252
rect 22468 30200 22520 30252
rect 24676 30243 24728 30252
rect 24676 30209 24685 30243
rect 24685 30209 24719 30243
rect 24719 30209 24728 30243
rect 24676 30200 24728 30209
rect 25688 30243 25740 30252
rect 25688 30209 25697 30243
rect 25697 30209 25731 30243
rect 25731 30209 25740 30243
rect 25688 30200 25740 30209
rect 27160 30243 27212 30252
rect 17776 30064 17828 30116
rect 14464 29996 14516 30048
rect 16580 29996 16632 30048
rect 18420 30064 18472 30116
rect 18512 30039 18564 30048
rect 18512 30005 18521 30039
rect 18521 30005 18555 30039
rect 18555 30005 18564 30039
rect 18512 29996 18564 30005
rect 20720 30132 20772 30184
rect 23388 30132 23440 30184
rect 27160 30209 27169 30243
rect 27169 30209 27203 30243
rect 27203 30209 27212 30243
rect 27160 30200 27212 30209
rect 27804 30243 27856 30252
rect 27804 30209 27813 30243
rect 27813 30209 27847 30243
rect 27847 30209 27856 30243
rect 27804 30200 27856 30209
rect 28540 30200 28592 30252
rect 32680 30243 32732 30252
rect 32680 30209 32689 30243
rect 32689 30209 32723 30243
rect 32723 30209 32732 30243
rect 32680 30200 32732 30209
rect 34152 30336 34204 30388
rect 35532 30336 35584 30388
rect 33416 30311 33468 30320
rect 33416 30277 33425 30311
rect 33425 30277 33459 30311
rect 33459 30277 33468 30311
rect 33416 30268 33468 30277
rect 34520 30268 34572 30320
rect 35348 30200 35400 30252
rect 36452 30243 36504 30252
rect 36452 30209 36470 30243
rect 36470 30209 36504 30243
rect 36452 30200 36504 30209
rect 37832 30243 37884 30252
rect 37832 30209 37866 30243
rect 37866 30209 37884 30243
rect 37832 30200 37884 30209
rect 39672 30243 39724 30252
rect 39672 30209 39706 30243
rect 39706 30209 39724 30243
rect 39672 30200 39724 30209
rect 42156 30200 42208 30252
rect 34336 30132 34388 30184
rect 34152 30064 34204 30116
rect 20812 29996 20864 30048
rect 20996 29996 21048 30048
rect 22284 29996 22336 30048
rect 28632 29996 28684 30048
rect 32680 30039 32732 30048
rect 32680 30005 32689 30039
rect 32689 30005 32723 30039
rect 32723 30005 32732 30039
rect 32680 29996 32732 30005
rect 34244 30039 34296 30048
rect 34244 30005 34253 30039
rect 34253 30005 34287 30039
rect 34287 30005 34296 30039
rect 34244 29996 34296 30005
rect 38568 30064 38620 30116
rect 37740 29996 37792 30048
rect 39580 29996 39632 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 8024 29792 8076 29844
rect 22468 29792 22520 29844
rect 14924 29724 14976 29776
rect 14464 29699 14516 29708
rect 14464 29665 14473 29699
rect 14473 29665 14507 29699
rect 14507 29665 14516 29699
rect 14464 29656 14516 29665
rect 14280 29631 14332 29640
rect 14280 29597 14289 29631
rect 14289 29597 14323 29631
rect 14323 29597 14332 29631
rect 14280 29588 14332 29597
rect 14556 29631 14608 29640
rect 14556 29597 14565 29631
rect 14565 29597 14599 29631
rect 14599 29597 14608 29631
rect 14556 29588 14608 29597
rect 14740 29631 14792 29640
rect 14740 29597 14749 29631
rect 14749 29597 14783 29631
rect 14783 29597 14792 29631
rect 14740 29588 14792 29597
rect 14924 29588 14976 29640
rect 15476 29631 15528 29640
rect 15476 29597 15485 29631
rect 15485 29597 15519 29631
rect 15519 29597 15528 29631
rect 15476 29588 15528 29597
rect 16764 29724 16816 29776
rect 18512 29724 18564 29776
rect 19800 29724 19852 29776
rect 22376 29724 22428 29776
rect 22928 29792 22980 29844
rect 25872 29835 25924 29844
rect 25872 29801 25881 29835
rect 25881 29801 25915 29835
rect 25915 29801 25924 29835
rect 25872 29792 25924 29801
rect 27068 29792 27120 29844
rect 27804 29792 27856 29844
rect 29736 29835 29788 29844
rect 29736 29801 29745 29835
rect 29745 29801 29779 29835
rect 29779 29801 29788 29835
rect 29736 29792 29788 29801
rect 23388 29724 23440 29776
rect 30656 29792 30708 29844
rect 33968 29835 34020 29844
rect 33968 29801 33977 29835
rect 33977 29801 34011 29835
rect 34011 29801 34020 29835
rect 33968 29792 34020 29801
rect 35440 29792 35492 29844
rect 37740 29835 37792 29844
rect 37740 29801 37749 29835
rect 37749 29801 37783 29835
rect 37783 29801 37792 29835
rect 37740 29792 37792 29801
rect 39672 29792 39724 29844
rect 15936 29631 15988 29640
rect 15936 29597 15945 29631
rect 15945 29597 15979 29631
rect 15979 29597 15988 29631
rect 15936 29588 15988 29597
rect 16212 29588 16264 29640
rect 18512 29631 18564 29640
rect 11980 29563 12032 29572
rect 11980 29529 12014 29563
rect 12014 29529 12032 29563
rect 11980 29520 12032 29529
rect 12072 29520 12124 29572
rect 18512 29597 18521 29631
rect 18521 29597 18555 29631
rect 18555 29597 18564 29631
rect 18512 29588 18564 29597
rect 18972 29588 19024 29640
rect 19248 29631 19300 29640
rect 19248 29597 19257 29631
rect 19257 29597 19291 29631
rect 19291 29597 19300 29631
rect 19248 29588 19300 29597
rect 25136 29656 25188 29708
rect 28448 29656 28500 29708
rect 29000 29699 29052 29708
rect 29000 29665 29009 29699
rect 29009 29665 29043 29699
rect 29043 29665 29052 29699
rect 29000 29656 29052 29665
rect 39120 29724 39172 29776
rect 18236 29563 18288 29572
rect 18236 29529 18254 29563
rect 18254 29529 18288 29563
rect 18236 29520 18288 29529
rect 18420 29520 18472 29572
rect 20444 29631 20496 29640
rect 20444 29597 20453 29631
rect 20453 29597 20487 29631
rect 20487 29597 20496 29631
rect 20444 29588 20496 29597
rect 20536 29520 20588 29572
rect 20812 29520 20864 29572
rect 23848 29520 23900 29572
rect 25136 29563 25188 29572
rect 25136 29529 25145 29563
rect 25145 29529 25179 29563
rect 25179 29529 25188 29563
rect 25136 29520 25188 29529
rect 30380 29631 30432 29640
rect 25780 29520 25832 29572
rect 30380 29597 30389 29631
rect 30389 29597 30423 29631
rect 30423 29597 30432 29631
rect 30380 29588 30432 29597
rect 32680 29588 32732 29640
rect 34704 29631 34756 29640
rect 34704 29597 34713 29631
rect 34713 29597 34747 29631
rect 34747 29597 34756 29631
rect 34704 29588 34756 29597
rect 39120 29631 39172 29640
rect 39120 29597 39129 29631
rect 39129 29597 39163 29631
rect 39163 29597 39172 29631
rect 39120 29588 39172 29597
rect 30012 29520 30064 29572
rect 34796 29520 34848 29572
rect 37924 29520 37976 29572
rect 39488 29520 39540 29572
rect 42064 29563 42116 29572
rect 42064 29529 42073 29563
rect 42073 29529 42107 29563
rect 42107 29529 42116 29563
rect 42064 29520 42116 29529
rect 13084 29495 13136 29504
rect 13084 29461 13093 29495
rect 13093 29461 13127 29495
rect 13127 29461 13136 29495
rect 13084 29452 13136 29461
rect 14096 29495 14148 29504
rect 14096 29461 14105 29495
rect 14105 29461 14139 29495
rect 14139 29461 14148 29495
rect 14096 29452 14148 29461
rect 15292 29495 15344 29504
rect 15292 29461 15301 29495
rect 15301 29461 15335 29495
rect 15335 29461 15344 29495
rect 15292 29452 15344 29461
rect 17132 29452 17184 29504
rect 20628 29452 20680 29504
rect 24952 29452 25004 29504
rect 25228 29452 25280 29504
rect 25504 29452 25556 29504
rect 29000 29452 29052 29504
rect 30748 29452 30800 29504
rect 37556 29495 37608 29504
rect 37556 29461 37565 29495
rect 37565 29461 37599 29495
rect 37599 29461 37608 29495
rect 37556 29452 37608 29461
rect 41972 29495 42024 29504
rect 41972 29461 41981 29495
rect 41981 29461 42015 29495
rect 42015 29461 42024 29495
rect 41972 29452 42024 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 15752 29291 15804 29300
rect 15752 29257 15761 29291
rect 15761 29257 15795 29291
rect 15795 29257 15804 29291
rect 15752 29248 15804 29257
rect 16212 29248 16264 29300
rect 20812 29291 20864 29300
rect 20812 29257 20821 29291
rect 20821 29257 20855 29291
rect 20855 29257 20864 29291
rect 20812 29248 20864 29257
rect 14096 29180 14148 29232
rect 16488 29180 16540 29232
rect 12072 29155 12124 29164
rect 12072 29121 12081 29155
rect 12081 29121 12115 29155
rect 12115 29121 12124 29155
rect 12072 29112 12124 29121
rect 13084 29112 13136 29164
rect 15476 29112 15528 29164
rect 16764 29155 16816 29164
rect 16764 29121 16773 29155
rect 16773 29121 16807 29155
rect 16807 29121 16816 29155
rect 16764 29112 16816 29121
rect 17224 29180 17276 29232
rect 18512 29180 18564 29232
rect 18696 29180 18748 29232
rect 19432 29223 19484 29232
rect 19432 29189 19441 29223
rect 19441 29189 19475 29223
rect 19475 29189 19484 29223
rect 19432 29180 19484 29189
rect 20444 29180 20496 29232
rect 20904 29112 20956 29164
rect 20996 29155 21048 29164
rect 20996 29121 21005 29155
rect 21005 29121 21039 29155
rect 21039 29121 21048 29155
rect 23388 29180 23440 29232
rect 26608 29248 26660 29300
rect 29736 29248 29788 29300
rect 30012 29248 30064 29300
rect 34796 29248 34848 29300
rect 37832 29291 37884 29300
rect 37832 29257 37841 29291
rect 37841 29257 37875 29291
rect 37875 29257 37884 29291
rect 37832 29248 37884 29257
rect 20996 29112 21048 29121
rect 24860 29180 24912 29232
rect 25780 29180 25832 29232
rect 25964 29180 26016 29232
rect 14004 29044 14056 29096
rect 22284 29044 22336 29096
rect 14740 28976 14792 29028
rect 17224 28976 17276 29028
rect 22376 28976 22428 29028
rect 22560 28976 22612 29028
rect 24584 28976 24636 29028
rect 28356 29155 28408 29164
rect 28356 29121 28365 29155
rect 28365 29121 28399 29155
rect 28399 29121 28408 29155
rect 28356 29112 28408 29121
rect 28540 29155 28592 29164
rect 28540 29121 28549 29155
rect 28549 29121 28583 29155
rect 28583 29121 28592 29155
rect 29184 29155 29236 29164
rect 28540 29112 28592 29121
rect 29184 29121 29193 29155
rect 29193 29121 29227 29155
rect 29227 29121 29236 29155
rect 29184 29112 29236 29121
rect 29368 29155 29420 29164
rect 29368 29121 29377 29155
rect 29377 29121 29411 29155
rect 29411 29121 29420 29155
rect 29368 29112 29420 29121
rect 30748 29155 30800 29164
rect 29092 29044 29144 29096
rect 30748 29121 30757 29155
rect 30757 29121 30791 29155
rect 30791 29121 30800 29155
rect 30748 29112 30800 29121
rect 34244 29112 34296 29164
rect 37556 29112 37608 29164
rect 1676 28951 1728 28960
rect 1676 28917 1685 28951
rect 1685 28917 1719 28951
rect 1719 28917 1728 28951
rect 1676 28908 1728 28917
rect 13452 28951 13504 28960
rect 13452 28917 13461 28951
rect 13461 28917 13495 28951
rect 13495 28917 13504 28951
rect 13452 28908 13504 28917
rect 15844 28908 15896 28960
rect 24308 28951 24360 28960
rect 24308 28917 24317 28951
rect 24317 28917 24351 28951
rect 24351 28917 24360 28951
rect 24308 28908 24360 28917
rect 26332 28908 26384 28960
rect 27160 28951 27212 28960
rect 27160 28917 27169 28951
rect 27169 28917 27203 28951
rect 27203 28917 27212 28951
rect 27160 28908 27212 28917
rect 41788 28951 41840 28960
rect 41788 28917 41797 28951
rect 41797 28917 41831 28951
rect 41831 28917 41840 28951
rect 41788 28908 41840 28917
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 14556 28704 14608 28756
rect 20904 28704 20956 28756
rect 21732 28747 21784 28756
rect 21732 28713 21741 28747
rect 21741 28713 21775 28747
rect 21775 28713 21784 28747
rect 21732 28704 21784 28713
rect 1676 28568 1728 28620
rect 2780 28611 2832 28620
rect 2780 28577 2789 28611
rect 2789 28577 2823 28611
rect 2823 28577 2832 28611
rect 2780 28568 2832 28577
rect 13452 28568 13504 28620
rect 14924 28636 14976 28688
rect 14372 28611 14424 28620
rect 14372 28577 14381 28611
rect 14381 28577 14415 28611
rect 14415 28577 14424 28611
rect 14372 28568 14424 28577
rect 15752 28568 15804 28620
rect 16396 28568 16448 28620
rect 14004 28500 14056 28552
rect 15844 28500 15896 28552
rect 16948 28500 17000 28552
rect 17408 28543 17460 28552
rect 17408 28509 17417 28543
rect 17417 28509 17451 28543
rect 17451 28509 17460 28543
rect 17408 28500 17460 28509
rect 19432 28568 19484 28620
rect 2136 28432 2188 28484
rect 15936 28432 15988 28484
rect 16488 28475 16540 28484
rect 16488 28441 16497 28475
rect 16497 28441 16531 28475
rect 16531 28441 16540 28475
rect 16488 28432 16540 28441
rect 20260 28432 20312 28484
rect 22652 28704 22704 28756
rect 26884 28704 26936 28756
rect 31668 28704 31720 28756
rect 22560 28636 22612 28688
rect 22468 28611 22520 28620
rect 22468 28577 22477 28611
rect 22477 28577 22511 28611
rect 22511 28577 22520 28611
rect 22468 28568 22520 28577
rect 23664 28636 23716 28688
rect 24860 28679 24912 28688
rect 24860 28645 24869 28679
rect 24869 28645 24903 28679
rect 24903 28645 24912 28679
rect 24860 28636 24912 28645
rect 28816 28679 28868 28688
rect 25964 28568 26016 28620
rect 22376 28543 22428 28552
rect 22376 28509 22385 28543
rect 22385 28509 22419 28543
rect 22419 28509 22428 28543
rect 22376 28500 22428 28509
rect 23848 28500 23900 28552
rect 26240 28500 26292 28552
rect 27160 28500 27212 28552
rect 28816 28645 28825 28679
rect 28825 28645 28859 28679
rect 28859 28645 28868 28679
rect 28816 28636 28868 28645
rect 29368 28636 29420 28688
rect 41328 28611 41380 28620
rect 23664 28432 23716 28484
rect 27896 28543 27948 28552
rect 27896 28509 27905 28543
rect 27905 28509 27939 28543
rect 27939 28509 27948 28543
rect 27896 28500 27948 28509
rect 28356 28500 28408 28552
rect 28632 28500 28684 28552
rect 41328 28577 41337 28611
rect 41337 28577 41371 28611
rect 41371 28577 41380 28611
rect 41328 28568 41380 28577
rect 41788 28568 41840 28620
rect 29184 28500 29236 28552
rect 29644 28500 29696 28552
rect 30380 28500 30432 28552
rect 30472 28432 30524 28484
rect 41420 28432 41472 28484
rect 14280 28364 14332 28416
rect 14556 28364 14608 28416
rect 17316 28364 17368 28416
rect 18236 28364 18288 28416
rect 21180 28364 21232 28416
rect 25688 28364 25740 28416
rect 25872 28407 25924 28416
rect 25872 28373 25881 28407
rect 25881 28373 25915 28407
rect 25915 28373 25924 28407
rect 25872 28364 25924 28373
rect 29000 28364 29052 28416
rect 29276 28364 29328 28416
rect 31392 28364 31444 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 2136 28203 2188 28212
rect 2136 28169 2145 28203
rect 2145 28169 2179 28203
rect 2179 28169 2188 28203
rect 2136 28160 2188 28169
rect 17776 28203 17828 28212
rect 14004 28092 14056 28144
rect 14648 28135 14700 28144
rect 14648 28101 14657 28135
rect 14657 28101 14691 28135
rect 14691 28101 14700 28135
rect 14648 28092 14700 28101
rect 17040 28135 17092 28144
rect 17040 28101 17049 28135
rect 17049 28101 17083 28135
rect 17083 28101 17092 28135
rect 17040 28092 17092 28101
rect 2596 28024 2648 28076
rect 12716 28067 12768 28076
rect 12716 28033 12725 28067
rect 12725 28033 12759 28067
rect 12759 28033 12768 28067
rect 12716 28024 12768 28033
rect 14464 28067 14516 28076
rect 14464 28033 14473 28067
rect 14473 28033 14507 28067
rect 14507 28033 14516 28067
rect 14464 28024 14516 28033
rect 14556 28024 14608 28076
rect 15844 28067 15896 28076
rect 15844 28033 15853 28067
rect 15853 28033 15887 28067
rect 15887 28033 15896 28067
rect 15844 28024 15896 28033
rect 15936 28067 15988 28076
rect 15936 28033 15945 28067
rect 15945 28033 15979 28067
rect 15979 28033 15988 28067
rect 15936 28024 15988 28033
rect 15660 27999 15712 28008
rect 15660 27965 15669 27999
rect 15669 27965 15703 27999
rect 15703 27965 15712 27999
rect 15660 27956 15712 27965
rect 17132 28024 17184 28076
rect 17316 28067 17368 28076
rect 17316 28033 17325 28067
rect 17325 28033 17359 28067
rect 17359 28033 17368 28067
rect 17776 28169 17785 28203
rect 17785 28169 17819 28203
rect 17819 28169 17828 28203
rect 17776 28160 17828 28169
rect 20260 28203 20312 28212
rect 20260 28169 20269 28203
rect 20269 28169 20303 28203
rect 20303 28169 20312 28203
rect 20260 28160 20312 28169
rect 26332 28203 26384 28212
rect 26332 28169 26341 28203
rect 26341 28169 26375 28203
rect 26375 28169 26384 28203
rect 26332 28160 26384 28169
rect 27896 28160 27948 28212
rect 28448 28160 28500 28212
rect 29644 28160 29696 28212
rect 30472 28160 30524 28212
rect 41420 28203 41472 28212
rect 41420 28169 41429 28203
rect 41429 28169 41463 28203
rect 41463 28169 41472 28203
rect 41420 28160 41472 28169
rect 20352 28092 20404 28144
rect 21732 28092 21784 28144
rect 25872 28092 25924 28144
rect 26056 28092 26108 28144
rect 17316 28024 17368 28033
rect 18236 28067 18288 28076
rect 18236 28033 18245 28067
rect 18245 28033 18279 28067
rect 18279 28033 18288 28067
rect 18788 28067 18840 28076
rect 18236 28024 18288 28033
rect 18788 28033 18797 28067
rect 18797 28033 18831 28067
rect 18831 28033 18840 28067
rect 18788 28024 18840 28033
rect 20444 28067 20496 28076
rect 20444 28033 20453 28067
rect 20453 28033 20487 28067
rect 20487 28033 20496 28067
rect 20444 28024 20496 28033
rect 24400 28024 24452 28076
rect 25780 28024 25832 28076
rect 28448 28067 28500 28076
rect 28448 28033 28457 28067
rect 28457 28033 28491 28067
rect 28491 28033 28500 28067
rect 28448 28024 28500 28033
rect 29092 28067 29144 28076
rect 29092 28033 29101 28067
rect 29101 28033 29135 28067
rect 29135 28033 29144 28067
rect 29092 28024 29144 28033
rect 32772 28135 32824 28144
rect 17868 27956 17920 28008
rect 18052 27999 18104 28008
rect 18052 27965 18061 27999
rect 18061 27965 18095 27999
rect 18095 27965 18104 27999
rect 18052 27956 18104 27965
rect 23664 27956 23716 28008
rect 29000 27956 29052 28008
rect 31300 28024 31352 28076
rect 31484 28024 31536 28076
rect 28816 27888 28868 27940
rect 29092 27888 29144 27940
rect 29276 27888 29328 27940
rect 29368 27888 29420 27940
rect 32772 28101 32781 28135
rect 32781 28101 32815 28135
rect 32815 28101 32824 28135
rect 32772 28092 32824 28101
rect 33232 28092 33284 28144
rect 32588 28067 32640 28076
rect 32588 28033 32597 28067
rect 32597 28033 32631 28067
rect 32631 28033 32640 28067
rect 32588 28024 32640 28033
rect 32864 28024 32916 28076
rect 41236 28024 41288 28076
rect 32496 27888 32548 27940
rect 12532 27863 12584 27872
rect 12532 27829 12541 27863
rect 12541 27829 12575 27863
rect 12575 27829 12584 27863
rect 12532 27820 12584 27829
rect 15108 27820 15160 27872
rect 16764 27820 16816 27872
rect 18972 27863 19024 27872
rect 18972 27829 18981 27863
rect 18981 27829 19015 27863
rect 19015 27829 19024 27863
rect 18972 27820 19024 27829
rect 26240 27820 26292 27872
rect 27436 27820 27488 27872
rect 28172 27820 28224 27872
rect 28632 27820 28684 27872
rect 30380 27820 30432 27872
rect 31668 27820 31720 27872
rect 33416 27863 33468 27872
rect 33416 27829 33425 27863
rect 33425 27829 33459 27863
rect 33459 27829 33468 27863
rect 33416 27820 33468 27829
rect 35624 27820 35676 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 17868 27616 17920 27668
rect 18052 27548 18104 27600
rect 18604 27591 18656 27600
rect 18604 27557 18613 27591
rect 18613 27557 18647 27591
rect 18647 27557 18656 27591
rect 18604 27548 18656 27557
rect 20168 27548 20220 27600
rect 20444 27616 20496 27668
rect 21180 27616 21232 27668
rect 24400 27659 24452 27668
rect 24400 27625 24409 27659
rect 24409 27625 24443 27659
rect 24443 27625 24452 27659
rect 24400 27616 24452 27625
rect 25964 27659 26016 27668
rect 25964 27625 25973 27659
rect 25973 27625 26007 27659
rect 26007 27625 26016 27659
rect 25964 27616 26016 27625
rect 28172 27659 28224 27668
rect 28172 27625 28181 27659
rect 28181 27625 28215 27659
rect 28215 27625 28224 27659
rect 28172 27616 28224 27625
rect 28816 27659 28868 27668
rect 28816 27625 28825 27659
rect 28825 27625 28859 27659
rect 28859 27625 28868 27659
rect 28816 27616 28868 27625
rect 29092 27616 29144 27668
rect 32588 27616 32640 27668
rect 22376 27591 22428 27600
rect 22376 27557 22385 27591
rect 22385 27557 22419 27591
rect 22419 27557 22428 27591
rect 22376 27548 22428 27557
rect 11888 27523 11940 27532
rect 11888 27489 11897 27523
rect 11897 27489 11931 27523
rect 11931 27489 11940 27523
rect 11888 27480 11940 27489
rect 16396 27523 16448 27532
rect 16396 27489 16405 27523
rect 16405 27489 16439 27523
rect 16439 27489 16448 27523
rect 16396 27480 16448 27489
rect 12532 27412 12584 27464
rect 14464 27455 14516 27464
rect 14464 27421 14473 27455
rect 14473 27421 14507 27455
rect 14507 27421 14516 27455
rect 14464 27412 14516 27421
rect 14648 27455 14700 27464
rect 14648 27421 14657 27455
rect 14657 27421 14691 27455
rect 14691 27421 14700 27455
rect 14648 27412 14700 27421
rect 15108 27455 15160 27464
rect 15108 27421 15117 27455
rect 15117 27421 15151 27455
rect 15151 27421 15160 27455
rect 15108 27412 15160 27421
rect 16488 27412 16540 27464
rect 17132 27480 17184 27532
rect 17408 27480 17460 27532
rect 23296 27480 23348 27532
rect 24492 27548 24544 27600
rect 25136 27548 25188 27600
rect 30104 27548 30156 27600
rect 17040 27412 17092 27464
rect 17592 27412 17644 27464
rect 20812 27412 20864 27464
rect 21180 27455 21232 27464
rect 21180 27421 21189 27455
rect 21189 27421 21223 27455
rect 21223 27421 21232 27455
rect 21180 27412 21232 27421
rect 21456 27455 21508 27464
rect 21456 27421 21465 27455
rect 21465 27421 21499 27455
rect 21499 27421 21508 27455
rect 21456 27412 21508 27421
rect 23204 27412 23256 27464
rect 24584 27455 24636 27464
rect 24584 27421 24593 27455
rect 24593 27421 24627 27455
rect 24627 27421 24636 27455
rect 24584 27412 24636 27421
rect 25044 27412 25096 27464
rect 25780 27412 25832 27464
rect 26056 27455 26108 27464
rect 26056 27421 26065 27455
rect 26065 27421 26099 27455
rect 26099 27421 26108 27455
rect 26056 27412 26108 27421
rect 27804 27412 27856 27464
rect 28908 27480 28960 27532
rect 29000 27480 29052 27532
rect 30196 27480 30248 27532
rect 31668 27480 31720 27532
rect 28540 27412 28592 27464
rect 28632 27412 28684 27464
rect 29092 27412 29144 27464
rect 29368 27412 29420 27464
rect 33416 27412 33468 27464
rect 41512 27412 41564 27464
rect 16764 27344 16816 27396
rect 18144 27344 18196 27396
rect 18788 27344 18840 27396
rect 20996 27344 21048 27396
rect 13268 27319 13320 27328
rect 13268 27285 13277 27319
rect 13277 27285 13311 27319
rect 13311 27285 13320 27319
rect 13268 27276 13320 27285
rect 21732 27276 21784 27328
rect 22560 27319 22612 27328
rect 22560 27285 22569 27319
rect 22569 27285 22603 27319
rect 22603 27285 22612 27319
rect 22560 27276 22612 27285
rect 27896 27344 27948 27396
rect 29000 27387 29052 27396
rect 29000 27353 29009 27387
rect 29009 27353 29043 27387
rect 29043 27353 29052 27387
rect 29000 27344 29052 27353
rect 26700 27319 26752 27328
rect 26700 27285 26709 27319
rect 26709 27285 26743 27319
rect 26743 27285 26752 27319
rect 26700 27276 26752 27285
rect 28632 27319 28684 27328
rect 28632 27285 28641 27319
rect 28641 27285 28675 27319
rect 28675 27285 28684 27319
rect 28632 27276 28684 27285
rect 28908 27276 28960 27328
rect 29828 27276 29880 27328
rect 30748 27344 30800 27396
rect 30288 27276 30340 27328
rect 31392 27319 31444 27328
rect 31392 27285 31401 27319
rect 31401 27285 31435 27319
rect 31435 27285 31444 27319
rect 31392 27276 31444 27285
rect 32772 27276 32824 27328
rect 34152 27319 34204 27328
rect 34152 27285 34161 27319
rect 34161 27285 34195 27319
rect 34195 27285 34204 27319
rect 34152 27276 34204 27285
rect 41696 27276 41748 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 12716 27072 12768 27124
rect 19432 27072 19484 27124
rect 23204 27115 23256 27124
rect 23204 27081 23213 27115
rect 23213 27081 23247 27115
rect 23247 27081 23256 27115
rect 23204 27072 23256 27081
rect 23296 27072 23348 27124
rect 14740 26936 14792 26988
rect 15292 26979 15344 26988
rect 15292 26945 15301 26979
rect 15301 26945 15335 26979
rect 15335 26945 15344 26979
rect 15292 26936 15344 26945
rect 13268 26868 13320 26920
rect 14464 26868 14516 26920
rect 15384 26843 15436 26852
rect 15384 26809 15393 26843
rect 15393 26809 15427 26843
rect 15427 26809 15436 26843
rect 15384 26800 15436 26809
rect 15660 26936 15712 26988
rect 16672 26979 16724 26988
rect 16672 26945 16681 26979
rect 16681 26945 16715 26979
rect 16715 26945 16724 26979
rect 16672 26936 16724 26945
rect 19524 26936 19576 26988
rect 16948 26911 17000 26920
rect 16948 26877 16957 26911
rect 16957 26877 16991 26911
rect 16991 26877 17000 26911
rect 16948 26868 17000 26877
rect 20812 27004 20864 27056
rect 23572 27004 23624 27056
rect 27804 27072 27856 27124
rect 27896 27072 27948 27124
rect 21916 26936 21968 26988
rect 23848 27047 23900 27056
rect 23848 27013 23873 27047
rect 23873 27013 23900 27047
rect 41972 27072 42024 27124
rect 23848 27004 23900 27013
rect 25596 26936 25648 26988
rect 28356 26936 28408 26988
rect 28816 26936 28868 26988
rect 29184 26979 29236 26988
rect 29184 26945 29193 26979
rect 29193 26945 29227 26979
rect 29227 26945 29236 26979
rect 29184 26936 29236 26945
rect 30748 26936 30800 26988
rect 31392 26979 31444 26988
rect 31392 26945 31401 26979
rect 31401 26945 31435 26979
rect 31435 26945 31444 26979
rect 31392 26936 31444 26945
rect 32864 26936 32916 26988
rect 33232 27004 33284 27056
rect 20996 26911 21048 26920
rect 20996 26877 21005 26911
rect 21005 26877 21039 26911
rect 21039 26877 21048 26911
rect 28448 26911 28500 26920
rect 20996 26868 21048 26877
rect 28448 26877 28457 26911
rect 28457 26877 28491 26911
rect 28491 26877 28500 26911
rect 28448 26868 28500 26877
rect 16856 26775 16908 26784
rect 16856 26741 16865 26775
rect 16865 26741 16899 26775
rect 16899 26741 16908 26775
rect 16856 26732 16908 26741
rect 19432 26732 19484 26784
rect 19708 26732 19760 26784
rect 30840 26868 30892 26920
rect 33784 26936 33836 26988
rect 34704 27004 34756 27056
rect 41696 27047 41748 27056
rect 41696 27013 41705 27047
rect 41705 27013 41739 27047
rect 41739 27013 41748 27047
rect 41696 27004 41748 27013
rect 33324 26868 33376 26920
rect 41328 26911 41380 26920
rect 41328 26877 41337 26911
rect 41337 26877 41371 26911
rect 41371 26877 41380 26911
rect 41328 26868 41380 26877
rect 41880 26911 41932 26920
rect 41880 26877 41889 26911
rect 41889 26877 41923 26911
rect 41923 26877 41932 26911
rect 41880 26868 41932 26877
rect 26332 26732 26384 26784
rect 30012 26732 30064 26784
rect 30288 26732 30340 26784
rect 32036 26732 32088 26784
rect 35348 26732 35400 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 15476 26528 15528 26580
rect 19524 26571 19576 26580
rect 19524 26537 19533 26571
rect 19533 26537 19567 26571
rect 19567 26537 19576 26571
rect 19524 26528 19576 26537
rect 20812 26528 20864 26580
rect 21916 26528 21968 26580
rect 25596 26571 25648 26580
rect 12072 26392 12124 26444
rect 14464 26460 14516 26512
rect 14740 26435 14792 26444
rect 14740 26401 14749 26435
rect 14749 26401 14783 26435
rect 14783 26401 14792 26435
rect 14740 26392 14792 26401
rect 15384 26460 15436 26512
rect 12900 26324 12952 26376
rect 15568 26324 15620 26376
rect 16396 26392 16448 26444
rect 15292 26256 15344 26308
rect 16764 26324 16816 26376
rect 19432 26392 19484 26444
rect 22560 26460 22612 26512
rect 23020 26460 23072 26512
rect 25596 26537 25605 26571
rect 25605 26537 25639 26571
rect 25639 26537 25648 26571
rect 25596 26528 25648 26537
rect 17408 26324 17460 26376
rect 19708 26367 19760 26376
rect 19708 26333 19717 26367
rect 19717 26333 19751 26367
rect 19751 26333 19760 26367
rect 19708 26324 19760 26333
rect 16672 26256 16724 26308
rect 16948 26256 17000 26308
rect 15200 26231 15252 26240
rect 15200 26197 15209 26231
rect 15209 26197 15243 26231
rect 15243 26197 15252 26231
rect 15200 26188 15252 26197
rect 20996 26324 21048 26376
rect 23204 26392 23256 26444
rect 23664 26392 23716 26444
rect 21456 26367 21508 26376
rect 21456 26333 21468 26367
rect 21468 26333 21502 26367
rect 21502 26333 21508 26367
rect 21456 26324 21508 26333
rect 21732 26324 21784 26376
rect 23848 26324 23900 26376
rect 24584 26367 24636 26376
rect 24584 26333 24593 26367
rect 24593 26333 24627 26367
rect 24627 26333 24636 26367
rect 24584 26324 24636 26333
rect 25044 26367 25096 26376
rect 25044 26333 25053 26367
rect 25053 26333 25087 26367
rect 25087 26333 25096 26367
rect 25044 26324 25096 26333
rect 26332 26367 26384 26376
rect 26332 26333 26366 26367
rect 26366 26333 26384 26367
rect 26332 26324 26384 26333
rect 28816 26528 28868 26580
rect 30288 26528 30340 26580
rect 31852 26528 31904 26580
rect 32772 26528 32824 26580
rect 33232 26528 33284 26580
rect 34060 26571 34112 26580
rect 34060 26537 34069 26571
rect 34069 26537 34103 26571
rect 34103 26537 34112 26571
rect 34060 26528 34112 26537
rect 41880 26528 41932 26580
rect 29368 26460 29420 26512
rect 29092 26392 29144 26444
rect 29828 26435 29880 26444
rect 29828 26401 29837 26435
rect 29837 26401 29871 26435
rect 29871 26401 29880 26435
rect 29828 26392 29880 26401
rect 28448 26324 28500 26376
rect 29000 26324 29052 26376
rect 32312 26460 32364 26512
rect 34704 26460 34756 26512
rect 30196 26392 30248 26444
rect 32588 26392 32640 26444
rect 30748 26367 30800 26376
rect 28540 26256 28592 26308
rect 30748 26333 30757 26367
rect 30757 26333 30791 26367
rect 30791 26333 30800 26367
rect 30748 26324 30800 26333
rect 32036 26367 32088 26376
rect 32036 26333 32045 26367
rect 32045 26333 32079 26367
rect 32079 26333 32088 26367
rect 32036 26324 32088 26333
rect 32496 26324 32548 26376
rect 34152 26367 34204 26376
rect 34152 26333 34161 26367
rect 34161 26333 34195 26367
rect 34195 26333 34204 26367
rect 34152 26324 34204 26333
rect 35348 26324 35400 26376
rect 33876 26256 33928 26308
rect 21548 26188 21600 26240
rect 24400 26231 24452 26240
rect 24400 26197 24409 26231
rect 24409 26197 24443 26231
rect 24443 26197 24452 26231
rect 24400 26188 24452 26197
rect 25412 26231 25464 26240
rect 25412 26197 25421 26231
rect 25421 26197 25455 26231
rect 25455 26197 25464 26231
rect 25412 26188 25464 26197
rect 27528 26188 27580 26240
rect 28724 26231 28776 26240
rect 28724 26197 28733 26231
rect 28733 26197 28767 26231
rect 28767 26197 28776 26231
rect 28724 26188 28776 26197
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 14740 25984 14792 26036
rect 15568 25984 15620 26036
rect 20812 26027 20864 26036
rect 20812 25993 20821 26027
rect 20821 25993 20855 26027
rect 20855 25993 20864 26027
rect 20812 25984 20864 25993
rect 21548 25984 21600 26036
rect 17868 25916 17920 25968
rect 21180 25959 21232 25968
rect 15200 25848 15252 25900
rect 16856 25848 16908 25900
rect 17960 25848 18012 25900
rect 18696 25891 18748 25900
rect 18696 25857 18705 25891
rect 18705 25857 18739 25891
rect 18739 25857 18748 25891
rect 18696 25848 18748 25857
rect 21180 25925 21189 25959
rect 21189 25925 21223 25959
rect 21223 25925 21232 25959
rect 21180 25916 21232 25925
rect 21456 25916 21508 25968
rect 24952 25984 25004 26036
rect 25412 25984 25464 26036
rect 28816 25984 28868 26036
rect 29000 26027 29052 26036
rect 29000 25993 29009 26027
rect 29009 25993 29043 26027
rect 29043 25993 29052 26027
rect 29000 25984 29052 25993
rect 30748 25984 30800 26036
rect 32864 25984 32916 26036
rect 33324 25984 33376 26036
rect 24400 25916 24452 25968
rect 27528 25916 27580 25968
rect 23020 25891 23072 25900
rect 23020 25857 23029 25891
rect 23029 25857 23063 25891
rect 23063 25857 23072 25891
rect 23020 25848 23072 25857
rect 23664 25891 23716 25900
rect 23664 25857 23673 25891
rect 23673 25857 23707 25891
rect 23707 25857 23716 25891
rect 23664 25848 23716 25857
rect 24308 25848 24360 25900
rect 15568 25780 15620 25832
rect 25504 25848 25556 25900
rect 26332 25848 26384 25900
rect 27896 25848 27948 25900
rect 28908 25848 28960 25900
rect 29184 25848 29236 25900
rect 29552 25848 29604 25900
rect 32312 25891 32364 25900
rect 32312 25857 32321 25891
rect 32321 25857 32355 25891
rect 32355 25857 32364 25891
rect 32312 25848 32364 25857
rect 33876 25891 33928 25900
rect 33876 25857 33885 25891
rect 33885 25857 33919 25891
rect 33919 25857 33928 25891
rect 33876 25848 33928 25857
rect 34060 25891 34112 25900
rect 34060 25857 34069 25891
rect 34069 25857 34103 25891
rect 34103 25857 34112 25891
rect 34060 25848 34112 25857
rect 15200 25712 15252 25764
rect 15844 25755 15896 25764
rect 15844 25721 15853 25755
rect 15853 25721 15887 25755
rect 15887 25721 15896 25755
rect 15844 25712 15896 25721
rect 26240 25712 26292 25764
rect 17592 25644 17644 25696
rect 21732 25644 21784 25696
rect 23296 25644 23348 25696
rect 25136 25644 25188 25696
rect 27160 25687 27212 25696
rect 27160 25653 27169 25687
rect 27169 25653 27203 25687
rect 27203 25653 27212 25687
rect 27160 25644 27212 25653
rect 31576 25780 31628 25832
rect 30380 25644 30432 25696
rect 30840 25644 30892 25696
rect 41880 25644 41932 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 15292 25440 15344 25492
rect 24584 25440 24636 25492
rect 25504 25483 25556 25492
rect 25504 25449 25513 25483
rect 25513 25449 25547 25483
rect 25547 25449 25556 25483
rect 25504 25440 25556 25449
rect 28724 25440 28776 25492
rect 30104 25483 30156 25492
rect 30104 25449 30113 25483
rect 30113 25449 30147 25483
rect 30147 25449 30156 25483
rect 30104 25440 30156 25449
rect 30472 25440 30524 25492
rect 33232 25440 33284 25492
rect 15292 25304 15344 25356
rect 14556 25279 14608 25288
rect 14556 25245 14565 25279
rect 14565 25245 14599 25279
rect 14599 25245 14608 25279
rect 15384 25279 15436 25288
rect 14556 25236 14608 25245
rect 15384 25245 15393 25279
rect 15393 25245 15427 25279
rect 15427 25245 15436 25279
rect 15384 25236 15436 25245
rect 15568 25279 15620 25288
rect 15568 25245 15577 25279
rect 15577 25245 15611 25279
rect 15611 25245 15620 25279
rect 16856 25304 16908 25356
rect 17592 25347 17644 25356
rect 17592 25313 17601 25347
rect 17601 25313 17635 25347
rect 17635 25313 17644 25347
rect 17592 25304 17644 25313
rect 24308 25304 24360 25356
rect 25136 25372 25188 25424
rect 31116 25372 31168 25424
rect 26240 25304 26292 25356
rect 26608 25347 26660 25356
rect 26608 25313 26617 25347
rect 26617 25313 26651 25347
rect 26651 25313 26660 25347
rect 26608 25304 26660 25313
rect 27160 25304 27212 25356
rect 15568 25236 15620 25245
rect 16764 25236 16816 25288
rect 17040 25236 17092 25288
rect 16396 25168 16448 25220
rect 20812 25236 20864 25288
rect 25688 25279 25740 25288
rect 25688 25245 25697 25279
rect 25697 25245 25731 25279
rect 25731 25245 25740 25279
rect 25688 25236 25740 25245
rect 28540 25279 28592 25288
rect 28540 25245 28549 25279
rect 28549 25245 28583 25279
rect 28583 25245 28592 25279
rect 28540 25236 28592 25245
rect 30656 25304 30708 25356
rect 30472 25236 30524 25288
rect 31300 25279 31352 25288
rect 31300 25245 31309 25279
rect 31309 25245 31343 25279
rect 31343 25245 31352 25279
rect 31576 25279 31628 25288
rect 31300 25236 31352 25245
rect 21272 25168 21324 25220
rect 27804 25168 27856 25220
rect 31576 25245 31585 25279
rect 31585 25245 31619 25279
rect 31619 25245 31628 25279
rect 31576 25236 31628 25245
rect 32404 25279 32456 25288
rect 32404 25245 32413 25279
rect 32413 25245 32447 25279
rect 32447 25245 32456 25279
rect 32404 25236 32456 25245
rect 33048 25236 33100 25288
rect 32772 25168 32824 25220
rect 33416 25236 33468 25288
rect 40040 25236 40092 25288
rect 41512 25236 41564 25288
rect 41788 25279 41840 25288
rect 41788 25245 41797 25279
rect 41797 25245 41831 25279
rect 41831 25245 41840 25279
rect 41788 25236 41840 25245
rect 40224 25168 40276 25220
rect 20168 25100 20220 25152
rect 23480 25100 23532 25152
rect 30288 25143 30340 25152
rect 30288 25109 30297 25143
rect 30297 25109 30331 25143
rect 30331 25109 30340 25143
rect 30288 25100 30340 25109
rect 30748 25100 30800 25152
rect 31576 25100 31628 25152
rect 31760 25143 31812 25152
rect 31760 25109 31769 25143
rect 31769 25109 31803 25143
rect 31803 25109 31812 25143
rect 31760 25100 31812 25109
rect 32680 25100 32732 25152
rect 33324 25143 33376 25152
rect 33324 25109 33333 25143
rect 33333 25109 33367 25143
rect 33367 25109 33376 25143
rect 33324 25100 33376 25109
rect 40500 25100 40552 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 14556 24896 14608 24948
rect 16028 24896 16080 24948
rect 25688 24939 25740 24948
rect 25688 24905 25715 24939
rect 25715 24905 25740 24939
rect 25688 24896 25740 24905
rect 26700 24896 26752 24948
rect 28448 24896 28500 24948
rect 29552 24939 29604 24948
rect 29552 24905 29561 24939
rect 29561 24905 29595 24939
rect 29595 24905 29604 24939
rect 29552 24896 29604 24905
rect 31116 24896 31168 24948
rect 31576 24896 31628 24948
rect 33048 24896 33100 24948
rect 15844 24871 15896 24880
rect 15844 24837 15879 24871
rect 15879 24837 15896 24871
rect 15844 24828 15896 24837
rect 27528 24828 27580 24880
rect 30564 24828 30616 24880
rect 12900 24803 12952 24812
rect 12900 24769 12909 24803
rect 12909 24769 12943 24803
rect 12943 24769 12952 24803
rect 12900 24760 12952 24769
rect 13452 24760 13504 24812
rect 14924 24803 14976 24812
rect 14924 24769 14933 24803
rect 14933 24769 14967 24803
rect 14967 24769 14976 24803
rect 14924 24760 14976 24769
rect 15476 24760 15528 24812
rect 16396 24760 16448 24812
rect 17040 24803 17092 24812
rect 17040 24769 17049 24803
rect 17049 24769 17083 24803
rect 17083 24769 17092 24803
rect 17040 24760 17092 24769
rect 17224 24760 17276 24812
rect 17408 24803 17460 24812
rect 17408 24769 17417 24803
rect 17417 24769 17451 24803
rect 17451 24769 17460 24803
rect 17408 24760 17460 24769
rect 18696 24760 18748 24812
rect 19616 24760 19668 24812
rect 22008 24760 22060 24812
rect 23388 24760 23440 24812
rect 27160 24803 27212 24812
rect 27160 24769 27169 24803
rect 27169 24769 27203 24803
rect 27203 24769 27212 24803
rect 27160 24760 27212 24769
rect 29368 24803 29420 24812
rect 15936 24692 15988 24744
rect 17132 24692 17184 24744
rect 21272 24692 21324 24744
rect 22468 24692 22520 24744
rect 25320 24692 25372 24744
rect 26608 24692 26660 24744
rect 29368 24769 29377 24803
rect 29377 24769 29411 24803
rect 29411 24769 29420 24803
rect 29368 24760 29420 24769
rect 30748 24692 30800 24744
rect 33324 24828 33376 24880
rect 40224 24871 40276 24880
rect 31760 24760 31812 24812
rect 32312 24803 32364 24812
rect 32312 24769 32321 24803
rect 32321 24769 32355 24803
rect 32355 24769 32364 24803
rect 32312 24760 32364 24769
rect 31576 24692 31628 24744
rect 32404 24692 32456 24744
rect 32772 24692 32824 24744
rect 34704 24760 34756 24812
rect 36360 24803 36412 24812
rect 36360 24769 36378 24803
rect 36378 24769 36412 24803
rect 40224 24837 40233 24871
rect 40233 24837 40267 24871
rect 40267 24837 40276 24871
rect 40224 24828 40276 24837
rect 36360 24760 36412 24769
rect 39304 24803 39356 24812
rect 39304 24769 39313 24803
rect 39313 24769 39347 24803
rect 39347 24769 39356 24803
rect 39304 24760 39356 24769
rect 40040 24803 40092 24812
rect 40040 24769 40049 24803
rect 40049 24769 40083 24803
rect 40083 24769 40092 24803
rect 40040 24760 40092 24769
rect 33048 24692 33100 24744
rect 41236 24735 41288 24744
rect 13912 24624 13964 24676
rect 13820 24556 13872 24608
rect 14188 24556 14240 24608
rect 16764 24556 16816 24608
rect 17960 24624 18012 24676
rect 25044 24624 25096 24676
rect 27436 24624 27488 24676
rect 18604 24556 18656 24608
rect 20904 24599 20956 24608
rect 20904 24565 20913 24599
rect 20913 24565 20947 24599
rect 20947 24565 20956 24599
rect 20904 24556 20956 24565
rect 22560 24599 22612 24608
rect 22560 24565 22569 24599
rect 22569 24565 22603 24599
rect 22603 24565 22612 24599
rect 22560 24556 22612 24565
rect 23204 24599 23256 24608
rect 23204 24565 23213 24599
rect 23213 24565 23247 24599
rect 23247 24565 23256 24599
rect 23204 24556 23256 24565
rect 26240 24556 26292 24608
rect 31300 24556 31352 24608
rect 31484 24556 31536 24608
rect 33232 24556 33284 24608
rect 41236 24701 41245 24735
rect 41245 24701 41279 24735
rect 41279 24701 41288 24735
rect 41236 24692 41288 24701
rect 40040 24556 40092 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 13452 24395 13504 24404
rect 13452 24361 13461 24395
rect 13461 24361 13495 24395
rect 13495 24361 13504 24395
rect 13452 24352 13504 24361
rect 14832 24352 14884 24404
rect 15292 24352 15344 24404
rect 15568 24395 15620 24404
rect 15568 24361 15577 24395
rect 15577 24361 15611 24395
rect 15611 24361 15620 24395
rect 15568 24352 15620 24361
rect 17132 24395 17184 24404
rect 17132 24361 17141 24395
rect 17141 24361 17175 24395
rect 17175 24361 17184 24395
rect 17132 24352 17184 24361
rect 19616 24395 19668 24404
rect 19616 24361 19625 24395
rect 19625 24361 19659 24395
rect 19659 24361 19668 24395
rect 19616 24352 19668 24361
rect 20812 24395 20864 24404
rect 20812 24361 20821 24395
rect 20821 24361 20855 24395
rect 20855 24361 20864 24395
rect 20812 24352 20864 24361
rect 23388 24395 23440 24404
rect 23388 24361 23397 24395
rect 23397 24361 23431 24395
rect 23431 24361 23440 24395
rect 23388 24352 23440 24361
rect 29644 24352 29696 24404
rect 30656 24352 30708 24404
rect 31484 24395 31536 24404
rect 31484 24361 31493 24395
rect 31493 24361 31527 24395
rect 31527 24361 31536 24395
rect 32680 24395 32732 24404
rect 31484 24352 31536 24361
rect 3608 24216 3660 24268
rect 5632 24259 5684 24268
rect 5632 24225 5641 24259
rect 5641 24225 5675 24259
rect 5675 24225 5684 24259
rect 5632 24216 5684 24225
rect 13820 24216 13872 24268
rect 13912 24148 13964 24200
rect 14924 24216 14976 24268
rect 3424 24080 3476 24132
rect 14464 24012 14516 24064
rect 15200 24012 15252 24064
rect 17132 24216 17184 24268
rect 18144 24216 18196 24268
rect 16948 24191 17000 24200
rect 15752 24123 15804 24132
rect 15752 24089 15761 24123
rect 15761 24089 15795 24123
rect 15795 24089 15804 24123
rect 15752 24080 15804 24089
rect 16948 24157 16957 24191
rect 16957 24157 16991 24191
rect 16991 24157 17000 24191
rect 16948 24148 17000 24157
rect 20168 24216 20220 24268
rect 16764 24080 16816 24132
rect 19432 24080 19484 24132
rect 20076 24191 20128 24200
rect 20076 24157 20085 24191
rect 20085 24157 20119 24191
rect 20119 24157 20128 24191
rect 20904 24284 20956 24336
rect 21180 24284 21232 24336
rect 26332 24284 26384 24336
rect 29276 24284 29328 24336
rect 32680 24361 32689 24395
rect 32689 24361 32723 24395
rect 32723 24361 32732 24395
rect 32680 24352 32732 24361
rect 33416 24352 33468 24404
rect 36360 24352 36412 24404
rect 37556 24327 37608 24336
rect 20628 24216 20680 24268
rect 23756 24259 23808 24268
rect 23756 24225 23765 24259
rect 23765 24225 23799 24259
rect 23799 24225 23808 24259
rect 23756 24216 23808 24225
rect 24032 24216 24084 24268
rect 25596 24216 25648 24268
rect 27160 24216 27212 24268
rect 28540 24216 28592 24268
rect 20076 24148 20128 24157
rect 20812 24148 20864 24200
rect 22376 24191 22428 24200
rect 22376 24157 22385 24191
rect 22385 24157 22419 24191
rect 22419 24157 22428 24191
rect 22376 24148 22428 24157
rect 22560 24148 22612 24200
rect 24400 24191 24452 24200
rect 24400 24157 24409 24191
rect 24409 24157 24443 24191
rect 24443 24157 24452 24191
rect 24400 24148 24452 24157
rect 24492 24191 24544 24200
rect 24492 24157 24501 24191
rect 24501 24157 24535 24191
rect 24535 24157 24544 24191
rect 24492 24148 24544 24157
rect 25688 24148 25740 24200
rect 26240 24148 26292 24200
rect 28264 24148 28316 24200
rect 28724 24191 28776 24200
rect 28724 24157 28733 24191
rect 28733 24157 28767 24191
rect 28767 24157 28776 24191
rect 28724 24148 28776 24157
rect 30380 24148 30432 24200
rect 30564 24148 30616 24200
rect 37556 24293 37565 24327
rect 37565 24293 37599 24327
rect 37599 24293 37608 24327
rect 37556 24284 37608 24293
rect 40040 24259 40092 24268
rect 31300 24191 31352 24200
rect 31300 24157 31309 24191
rect 31309 24157 31343 24191
rect 31343 24157 31352 24191
rect 31300 24148 31352 24157
rect 31760 24148 31812 24200
rect 33232 24148 33284 24200
rect 40040 24225 40049 24259
rect 40049 24225 40083 24259
rect 40083 24225 40092 24259
rect 40040 24216 40092 24225
rect 40408 24216 40460 24268
rect 38660 24148 38712 24200
rect 39120 24191 39172 24200
rect 39120 24157 39129 24191
rect 39129 24157 39163 24191
rect 39163 24157 39172 24191
rect 39120 24148 39172 24157
rect 22008 24080 22060 24132
rect 26976 24080 27028 24132
rect 28172 24080 28224 24132
rect 28908 24080 28960 24132
rect 29184 24080 29236 24132
rect 32312 24080 32364 24132
rect 18052 24055 18104 24064
rect 18052 24021 18061 24055
rect 18061 24021 18095 24055
rect 18095 24021 18104 24055
rect 18052 24012 18104 24021
rect 20812 24012 20864 24064
rect 21088 24055 21140 24064
rect 21088 24021 21097 24055
rect 21097 24021 21131 24055
rect 21131 24021 21140 24055
rect 24676 24055 24728 24064
rect 21088 24012 21140 24021
rect 24676 24021 24685 24055
rect 24685 24021 24719 24055
rect 24719 24021 24728 24055
rect 24676 24012 24728 24021
rect 28356 24012 28408 24064
rect 29368 24012 29420 24064
rect 29460 24012 29512 24064
rect 30932 24012 30984 24064
rect 31116 24055 31168 24064
rect 31116 24021 31125 24055
rect 31125 24021 31159 24055
rect 31159 24021 31168 24055
rect 31116 24012 31168 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 3424 23851 3476 23860
rect 3424 23817 3433 23851
rect 3433 23817 3467 23851
rect 3467 23817 3476 23851
rect 3424 23808 3476 23817
rect 16028 23808 16080 23860
rect 20076 23808 20128 23860
rect 21548 23808 21600 23860
rect 22376 23808 22428 23860
rect 24400 23808 24452 23860
rect 25596 23851 25648 23860
rect 25596 23817 25605 23851
rect 25605 23817 25639 23851
rect 25639 23817 25648 23851
rect 25596 23808 25648 23817
rect 27344 23808 27396 23860
rect 3332 23715 3384 23724
rect 3332 23681 3341 23715
rect 3341 23681 3375 23715
rect 3375 23681 3384 23715
rect 3332 23672 3384 23681
rect 14464 23672 14516 23724
rect 17040 23672 17092 23724
rect 17684 23715 17736 23724
rect 17684 23681 17718 23715
rect 17718 23681 17736 23715
rect 17684 23672 17736 23681
rect 14372 23647 14424 23656
rect 14372 23613 14381 23647
rect 14381 23613 14415 23647
rect 14415 23613 14424 23647
rect 14372 23604 14424 23613
rect 16672 23604 16724 23656
rect 15752 23579 15804 23588
rect 15752 23545 15761 23579
rect 15761 23545 15795 23579
rect 15795 23545 15804 23579
rect 15752 23536 15804 23545
rect 20628 23672 20680 23724
rect 20720 23672 20772 23724
rect 21272 23740 21324 23792
rect 23204 23740 23256 23792
rect 24676 23740 24728 23792
rect 23848 23672 23900 23724
rect 25136 23715 25188 23724
rect 25136 23681 25145 23715
rect 25145 23681 25179 23715
rect 25179 23681 25188 23715
rect 25136 23672 25188 23681
rect 20812 23604 20864 23656
rect 21088 23647 21140 23656
rect 21088 23613 21097 23647
rect 21097 23613 21131 23647
rect 21131 23613 21140 23647
rect 21088 23604 21140 23613
rect 21180 23647 21232 23656
rect 21180 23613 21189 23647
rect 21189 23613 21223 23647
rect 21223 23613 21232 23647
rect 21180 23604 21232 23613
rect 22008 23604 22060 23656
rect 22468 23647 22520 23656
rect 22468 23613 22477 23647
rect 22477 23613 22511 23647
rect 22511 23613 22520 23647
rect 22468 23604 22520 23613
rect 19800 23579 19852 23588
rect 19800 23545 19809 23579
rect 19809 23545 19843 23579
rect 19843 23545 19852 23579
rect 19800 23536 19852 23545
rect 21364 23536 21416 23588
rect 24860 23604 24912 23656
rect 26700 23672 26752 23724
rect 26976 23715 27028 23724
rect 26976 23681 26985 23715
rect 26985 23681 27019 23715
rect 27019 23681 27028 23715
rect 26976 23672 27028 23681
rect 27160 23715 27212 23724
rect 27160 23681 27169 23715
rect 27169 23681 27203 23715
rect 27203 23681 27212 23715
rect 27160 23672 27212 23681
rect 27436 23672 27488 23724
rect 28172 23715 28224 23724
rect 28172 23681 28181 23715
rect 28181 23681 28215 23715
rect 28215 23681 28224 23715
rect 28172 23672 28224 23681
rect 29460 23808 29512 23860
rect 31300 23808 31352 23860
rect 28724 23740 28776 23792
rect 28540 23715 28592 23724
rect 28540 23681 28549 23715
rect 28549 23681 28583 23715
rect 28583 23681 28592 23715
rect 29276 23715 29328 23724
rect 28540 23672 28592 23681
rect 29276 23681 29285 23715
rect 29285 23681 29319 23715
rect 29319 23681 29328 23715
rect 29276 23672 29328 23681
rect 29368 23672 29420 23724
rect 27252 23647 27304 23656
rect 27252 23613 27261 23647
rect 27261 23613 27295 23647
rect 27295 23613 27304 23647
rect 27252 23604 27304 23613
rect 27344 23647 27396 23656
rect 27344 23613 27353 23647
rect 27353 23613 27387 23647
rect 27387 23613 27396 23647
rect 27344 23604 27396 23613
rect 29184 23604 29236 23656
rect 30564 23647 30616 23656
rect 30564 23613 30573 23647
rect 30573 23613 30607 23647
rect 30607 23613 30616 23647
rect 30564 23604 30616 23613
rect 30932 23604 30984 23656
rect 31484 23672 31536 23724
rect 32220 23715 32272 23724
rect 32220 23681 32229 23715
rect 32229 23681 32263 23715
rect 32263 23681 32272 23715
rect 32220 23672 32272 23681
rect 34704 23672 34756 23724
rect 35348 23672 35400 23724
rect 38016 23715 38068 23724
rect 38016 23681 38050 23715
rect 38050 23681 38068 23715
rect 38016 23672 38068 23681
rect 41880 23715 41932 23724
rect 41880 23681 41889 23715
rect 41889 23681 41923 23715
rect 41923 23681 41932 23715
rect 41880 23672 41932 23681
rect 31760 23604 31812 23656
rect 32312 23604 32364 23656
rect 41328 23647 41380 23656
rect 20904 23468 20956 23520
rect 21916 23468 21968 23520
rect 29552 23536 29604 23588
rect 29644 23536 29696 23588
rect 41328 23613 41337 23647
rect 41337 23613 41371 23647
rect 41371 23613 41380 23647
rect 41328 23604 41380 23613
rect 41696 23647 41748 23656
rect 41696 23613 41705 23647
rect 41705 23613 41739 23647
rect 41739 23613 41748 23647
rect 41696 23604 41748 23613
rect 27344 23468 27396 23520
rect 30104 23468 30156 23520
rect 30380 23511 30432 23520
rect 30380 23477 30389 23511
rect 30389 23477 30423 23511
rect 30423 23477 30432 23511
rect 30380 23468 30432 23477
rect 39028 23468 39080 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 19432 23307 19484 23316
rect 19432 23273 19441 23307
rect 19441 23273 19475 23307
rect 19475 23273 19484 23307
rect 19432 23264 19484 23273
rect 20812 23307 20864 23316
rect 20812 23273 20821 23307
rect 20821 23273 20855 23307
rect 20855 23273 20864 23307
rect 20812 23264 20864 23273
rect 24860 23264 24912 23316
rect 26240 23264 26292 23316
rect 26884 23307 26936 23316
rect 26884 23273 26893 23307
rect 26893 23273 26927 23307
rect 26927 23273 26936 23307
rect 26884 23264 26936 23273
rect 32220 23307 32272 23316
rect 22008 23196 22060 23248
rect 17868 23171 17920 23180
rect 17868 23137 17877 23171
rect 17877 23137 17911 23171
rect 17911 23137 17920 23171
rect 17868 23128 17920 23137
rect 1400 23060 1452 23112
rect 18144 23103 18196 23112
rect 18144 23069 18153 23103
rect 18153 23069 18187 23103
rect 18187 23069 18196 23103
rect 18144 23060 18196 23069
rect 20168 23128 20220 23180
rect 23388 23171 23440 23180
rect 19800 23103 19852 23112
rect 19800 23069 19809 23103
rect 19809 23069 19843 23103
rect 19843 23069 19852 23103
rect 19800 23060 19852 23069
rect 20720 23060 20772 23112
rect 23388 23137 23397 23171
rect 23397 23137 23431 23171
rect 23431 23137 23440 23171
rect 23388 23128 23440 23137
rect 24400 23171 24452 23180
rect 24400 23137 24409 23171
rect 24409 23137 24443 23171
rect 24443 23137 24452 23171
rect 24400 23128 24452 23137
rect 26332 23196 26384 23248
rect 32220 23273 32229 23307
rect 32229 23273 32263 23307
rect 32263 23273 32272 23307
rect 32220 23264 32272 23273
rect 38660 23307 38712 23316
rect 38660 23273 38669 23307
rect 38669 23273 38703 23307
rect 38703 23273 38712 23307
rect 38660 23264 38712 23273
rect 28816 23128 28868 23180
rect 29552 23171 29604 23180
rect 29552 23137 29561 23171
rect 29561 23137 29595 23171
rect 29595 23137 29604 23171
rect 29552 23128 29604 23137
rect 20628 22992 20680 23044
rect 20904 23035 20956 23044
rect 20904 23001 20913 23035
rect 20913 23001 20947 23035
rect 20947 23001 20956 23035
rect 20904 22992 20956 23001
rect 21180 22992 21232 23044
rect 23296 23103 23348 23112
rect 23296 23069 23305 23103
rect 23305 23069 23339 23103
rect 23339 23069 23348 23103
rect 23296 23060 23348 23069
rect 23848 23060 23900 23112
rect 24492 23060 24544 23112
rect 32404 23196 32456 23248
rect 30380 23128 30432 23180
rect 30840 23171 30892 23180
rect 30840 23137 30849 23171
rect 30849 23137 30883 23171
rect 30883 23137 30892 23171
rect 30840 23128 30892 23137
rect 34704 23128 34756 23180
rect 39396 23196 39448 23248
rect 40500 23171 40552 23180
rect 24216 22992 24268 23044
rect 24400 22992 24452 23044
rect 26976 22992 27028 23044
rect 31116 23103 31168 23112
rect 31116 23069 31150 23103
rect 31150 23069 31168 23103
rect 31116 23060 31168 23069
rect 40500 23137 40509 23171
rect 40509 23137 40543 23171
rect 40543 23137 40552 23171
rect 40500 23128 40552 23137
rect 38936 23060 38988 23112
rect 39948 23060 40000 23112
rect 40316 23103 40368 23112
rect 40316 23069 40325 23103
rect 40325 23069 40359 23103
rect 40359 23069 40368 23103
rect 40316 23060 40368 23069
rect 28816 22967 28868 22976
rect 28816 22933 28825 22967
rect 28825 22933 28859 22967
rect 28859 22933 28868 22967
rect 28816 22924 28868 22933
rect 30472 22992 30524 23044
rect 34888 22992 34940 23044
rect 37096 23035 37148 23044
rect 37096 23001 37130 23035
rect 37130 23001 37148 23035
rect 37096 22992 37148 23001
rect 39580 22924 39632 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 17684 22720 17736 22772
rect 20628 22720 20680 22772
rect 21456 22652 21508 22704
rect 2136 22627 2188 22636
rect 2136 22593 2145 22627
rect 2145 22593 2179 22627
rect 2179 22593 2188 22627
rect 2136 22584 2188 22593
rect 9220 22584 9272 22636
rect 18052 22627 18104 22636
rect 18052 22593 18061 22627
rect 18061 22593 18095 22627
rect 18095 22593 18104 22627
rect 18052 22584 18104 22593
rect 18604 22627 18656 22636
rect 18604 22593 18613 22627
rect 18613 22593 18647 22627
rect 18647 22593 18656 22627
rect 18604 22584 18656 22593
rect 20904 22584 20956 22636
rect 22744 22516 22796 22568
rect 23848 22627 23900 22636
rect 23848 22593 23857 22627
rect 23857 22593 23891 22627
rect 23891 22593 23900 22627
rect 27252 22720 27304 22772
rect 40316 22720 40368 22772
rect 26332 22652 26384 22704
rect 34704 22652 34756 22704
rect 23848 22584 23900 22593
rect 26976 22627 27028 22636
rect 25136 22516 25188 22568
rect 26976 22593 26985 22627
rect 26985 22593 27019 22627
rect 27019 22593 27028 22627
rect 26976 22584 27028 22593
rect 27160 22627 27212 22636
rect 27160 22593 27169 22627
rect 27169 22593 27203 22627
rect 27203 22593 27212 22627
rect 27160 22584 27212 22593
rect 27528 22627 27580 22636
rect 27528 22593 27537 22627
rect 27537 22593 27571 22627
rect 27571 22593 27580 22627
rect 28356 22627 28408 22636
rect 27528 22584 27580 22593
rect 28356 22593 28365 22627
rect 28365 22593 28399 22627
rect 28399 22593 28408 22627
rect 28356 22584 28408 22593
rect 28448 22627 28500 22636
rect 28448 22593 28457 22627
rect 28457 22593 28491 22627
rect 28491 22593 28500 22627
rect 29092 22627 29144 22636
rect 28448 22584 28500 22593
rect 29092 22593 29101 22627
rect 29101 22593 29135 22627
rect 29135 22593 29144 22627
rect 29092 22584 29144 22593
rect 29184 22627 29236 22636
rect 29184 22593 29193 22627
rect 29193 22593 29227 22627
rect 29227 22593 29236 22627
rect 29184 22584 29236 22593
rect 29828 22584 29880 22636
rect 23388 22448 23440 22500
rect 27344 22559 27396 22568
rect 27344 22525 27353 22559
rect 27353 22525 27387 22559
rect 27387 22525 27396 22559
rect 27344 22516 27396 22525
rect 29552 22516 29604 22568
rect 31392 22584 31444 22636
rect 32128 22627 32180 22636
rect 32128 22593 32137 22627
rect 32137 22593 32171 22627
rect 32171 22593 32180 22627
rect 32128 22584 32180 22593
rect 32220 22584 32272 22636
rect 32404 22627 32456 22636
rect 32404 22593 32413 22627
rect 32413 22593 32447 22627
rect 32447 22593 32456 22627
rect 32404 22584 32456 22593
rect 34520 22584 34572 22636
rect 29736 22448 29788 22500
rect 1584 22380 1636 22432
rect 19064 22380 19116 22432
rect 27160 22380 27212 22432
rect 28724 22380 28776 22432
rect 32864 22380 32916 22432
rect 38844 22584 38896 22636
rect 39948 22584 40000 22636
rect 41972 22584 42024 22636
rect 40684 22380 40736 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 18604 22176 18656 22228
rect 21732 22176 21784 22228
rect 22744 22219 22796 22228
rect 22744 22185 22753 22219
rect 22753 22185 22787 22219
rect 22787 22185 22796 22219
rect 22744 22176 22796 22185
rect 24492 22219 24544 22228
rect 24492 22185 24501 22219
rect 24501 22185 24535 22219
rect 24535 22185 24544 22219
rect 24492 22176 24544 22185
rect 26976 22176 27028 22228
rect 29644 22176 29696 22228
rect 29828 22219 29880 22228
rect 29828 22185 29837 22219
rect 29837 22185 29871 22219
rect 29871 22185 29880 22219
rect 29828 22176 29880 22185
rect 32128 22176 32180 22228
rect 1400 22083 1452 22092
rect 1400 22049 1409 22083
rect 1409 22049 1443 22083
rect 1443 22049 1452 22083
rect 1400 22040 1452 22049
rect 1584 22083 1636 22092
rect 1584 22049 1593 22083
rect 1593 22049 1627 22083
rect 1627 22049 1636 22083
rect 1584 22040 1636 22049
rect 1860 22083 1912 22092
rect 1860 22049 1869 22083
rect 1869 22049 1903 22083
rect 1903 22049 1912 22083
rect 1860 22040 1912 22049
rect 15660 22040 15712 22092
rect 16212 22083 16264 22092
rect 16212 22049 16221 22083
rect 16221 22049 16255 22083
rect 16255 22049 16264 22083
rect 16212 22040 16264 22049
rect 17868 22108 17920 22160
rect 20720 22151 20772 22160
rect 20720 22117 20729 22151
rect 20729 22117 20763 22151
rect 20763 22117 20772 22151
rect 20720 22108 20772 22117
rect 23388 22108 23440 22160
rect 12900 21972 12952 22024
rect 14372 21972 14424 22024
rect 15476 22015 15528 22024
rect 15476 21981 15485 22015
rect 15485 21981 15519 22015
rect 15519 21981 15528 22015
rect 15476 21972 15528 21981
rect 15844 21972 15896 22024
rect 17960 22015 18012 22024
rect 17960 21981 17969 22015
rect 17969 21981 18003 22015
rect 18003 21981 18012 22015
rect 17960 21972 18012 21981
rect 18144 21972 18196 22024
rect 15384 21904 15436 21956
rect 20904 22015 20956 22024
rect 20904 21981 20913 22015
rect 20913 21981 20947 22015
rect 20947 21981 20956 22015
rect 20904 21972 20956 21981
rect 21364 22015 21416 22024
rect 21364 21981 21373 22015
rect 21373 21981 21407 22015
rect 21407 21981 21416 22015
rect 21364 21972 21416 21981
rect 22008 21972 22060 22024
rect 24216 21972 24268 22024
rect 25136 22108 25188 22160
rect 26056 21972 26108 22024
rect 21824 21904 21876 21956
rect 25964 21947 26016 21956
rect 25964 21913 25973 21947
rect 25973 21913 26007 21947
rect 26007 21913 26016 21947
rect 25964 21904 26016 21913
rect 28356 22108 28408 22160
rect 27804 22083 27856 22092
rect 27804 22049 27813 22083
rect 27813 22049 27847 22083
rect 27847 22049 27856 22083
rect 27804 22040 27856 22049
rect 28172 22040 28224 22092
rect 28954 22108 29006 22160
rect 29552 22108 29604 22160
rect 29736 22083 29788 22092
rect 29736 22049 29745 22083
rect 29745 22049 29779 22083
rect 29779 22049 29788 22083
rect 29736 22040 29788 22049
rect 32404 22108 32456 22160
rect 28448 21972 28500 22024
rect 28908 21981 28917 22002
rect 28917 21981 28951 22002
rect 28951 21981 28960 22002
rect 28908 21950 28960 21981
rect 29000 21972 29052 22024
rect 15108 21836 15160 21888
rect 19984 21836 20036 21888
rect 20628 21836 20680 21888
rect 22928 21836 22980 21888
rect 29736 21904 29788 21956
rect 30196 21972 30248 22024
rect 30288 21972 30340 22024
rect 32220 21972 32272 22024
rect 32312 21972 32364 22024
rect 32864 21972 32916 22024
rect 28172 21836 28224 21888
rect 29460 21836 29512 21888
rect 30288 21836 30340 21888
rect 38936 22040 38988 22092
rect 39304 22083 39356 22092
rect 34796 21972 34848 22024
rect 35532 21972 35584 22024
rect 39028 22015 39080 22024
rect 35348 21904 35400 21956
rect 35716 21904 35768 21956
rect 39028 21981 39037 22015
rect 39037 21981 39071 22015
rect 39071 21981 39080 22015
rect 39028 21972 39080 21981
rect 39304 22049 39313 22083
rect 39313 22049 39347 22083
rect 39347 22049 39356 22083
rect 39304 22040 39356 22049
rect 40684 22040 40736 22092
rect 42156 22083 42208 22092
rect 42156 22049 42165 22083
rect 42165 22049 42199 22083
rect 42199 22049 42208 22083
rect 42156 22040 42208 22049
rect 39672 21972 39724 22024
rect 36360 21879 36412 21888
rect 36360 21845 36369 21879
rect 36369 21845 36403 21879
rect 36403 21845 36412 21879
rect 36360 21836 36412 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 14372 21632 14424 21684
rect 16212 21632 16264 21684
rect 20904 21632 20956 21684
rect 22928 21675 22980 21684
rect 22928 21641 22937 21675
rect 22937 21641 22971 21675
rect 22971 21641 22980 21675
rect 22928 21632 22980 21641
rect 24124 21632 24176 21684
rect 24400 21632 24452 21684
rect 26056 21675 26108 21684
rect 26056 21641 26065 21675
rect 26065 21641 26099 21675
rect 26099 21641 26108 21675
rect 26056 21632 26108 21641
rect 19064 21564 19116 21616
rect 20720 21564 20772 21616
rect 21916 21564 21968 21616
rect 29000 21632 29052 21684
rect 29736 21675 29788 21684
rect 29736 21641 29745 21675
rect 29745 21641 29779 21675
rect 29779 21641 29788 21675
rect 29736 21632 29788 21641
rect 32404 21632 32456 21684
rect 32588 21632 32640 21684
rect 38844 21632 38896 21684
rect 6368 21539 6420 21548
rect 6368 21505 6377 21539
rect 6377 21505 6411 21539
rect 6411 21505 6420 21539
rect 6368 21496 6420 21505
rect 14740 21539 14792 21548
rect 14740 21505 14749 21539
rect 14749 21505 14783 21539
rect 14783 21505 14792 21539
rect 14740 21496 14792 21505
rect 15108 21496 15160 21548
rect 15476 21496 15528 21548
rect 16672 21539 16724 21548
rect 16672 21505 16681 21539
rect 16681 21505 16715 21539
rect 16715 21505 16724 21539
rect 16672 21496 16724 21505
rect 17224 21496 17276 21548
rect 18788 21496 18840 21548
rect 23480 21496 23532 21548
rect 24400 21496 24452 21548
rect 1860 21471 1912 21480
rect 1860 21437 1869 21471
rect 1869 21437 1903 21471
rect 1903 21437 1912 21471
rect 1860 21428 1912 21437
rect 2688 21428 2740 21480
rect 2780 21471 2832 21480
rect 2780 21437 2789 21471
rect 2789 21437 2823 21471
rect 2823 21437 2832 21471
rect 7104 21471 7156 21480
rect 2780 21428 2832 21437
rect 7104 21437 7113 21471
rect 7113 21437 7147 21471
rect 7147 21437 7156 21471
rect 7104 21428 7156 21437
rect 15844 21428 15896 21480
rect 24676 21496 24728 21548
rect 27620 21564 27672 21616
rect 28356 21564 28408 21616
rect 27528 21539 27580 21548
rect 21824 21403 21876 21412
rect 21824 21369 21833 21403
rect 21833 21369 21867 21403
rect 21867 21369 21876 21403
rect 21824 21360 21876 21369
rect 17592 21292 17644 21344
rect 20812 21292 20864 21344
rect 24768 21428 24820 21480
rect 24584 21360 24636 21412
rect 27528 21505 27537 21539
rect 27537 21505 27571 21539
rect 27571 21505 27580 21539
rect 27528 21496 27580 21505
rect 28172 21496 28224 21548
rect 28540 21539 28592 21548
rect 28540 21505 28549 21539
rect 28549 21505 28583 21539
rect 28583 21505 28592 21539
rect 28540 21496 28592 21505
rect 30564 21564 30616 21616
rect 33048 21564 33100 21616
rect 41880 21607 41932 21616
rect 29276 21539 29328 21548
rect 29276 21505 29285 21539
rect 29285 21505 29319 21539
rect 29319 21505 29328 21539
rect 29276 21496 29328 21505
rect 30656 21496 30708 21548
rect 35532 21539 35584 21548
rect 35532 21505 35541 21539
rect 35541 21505 35575 21539
rect 35575 21505 35584 21539
rect 35532 21496 35584 21505
rect 35716 21539 35768 21548
rect 35716 21505 35725 21539
rect 35725 21505 35759 21539
rect 35759 21505 35768 21539
rect 35716 21496 35768 21505
rect 41880 21573 41889 21607
rect 41889 21573 41923 21607
rect 41923 21573 41932 21607
rect 41880 21564 41932 21573
rect 36360 21539 36412 21548
rect 36360 21505 36369 21539
rect 36369 21505 36403 21539
rect 36403 21505 36412 21539
rect 36360 21496 36412 21505
rect 28448 21428 28500 21480
rect 33692 21428 33744 21480
rect 37280 21428 37332 21480
rect 39672 21496 39724 21548
rect 39304 21428 39356 21480
rect 40960 21428 41012 21480
rect 27896 21360 27948 21412
rect 30288 21360 30340 21412
rect 32496 21360 32548 21412
rect 38476 21360 38528 21412
rect 24676 21292 24728 21344
rect 25136 21335 25188 21344
rect 25136 21301 25145 21335
rect 25145 21301 25179 21335
rect 25179 21301 25188 21335
rect 25136 21292 25188 21301
rect 29276 21292 29328 21344
rect 32220 21292 32272 21344
rect 34796 21292 34848 21344
rect 36176 21335 36228 21344
rect 36176 21301 36185 21335
rect 36185 21301 36219 21335
rect 36219 21301 36228 21335
rect 36176 21292 36228 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 1860 21088 1912 21140
rect 2688 21131 2740 21140
rect 2688 21097 2697 21131
rect 2697 21097 2731 21131
rect 2731 21097 2740 21131
rect 2688 21088 2740 21097
rect 7472 21131 7524 21140
rect 7472 21097 7481 21131
rect 7481 21097 7515 21131
rect 7515 21097 7524 21131
rect 7472 21088 7524 21097
rect 8116 21088 8168 21140
rect 15384 21088 15436 21140
rect 17224 21131 17276 21140
rect 17224 21097 17233 21131
rect 17233 21097 17267 21131
rect 17267 21097 17276 21131
rect 17224 21088 17276 21097
rect 20812 21131 20864 21140
rect 3332 20884 3384 20936
rect 5724 20927 5776 20936
rect 5724 20893 5733 20927
rect 5733 20893 5767 20927
rect 5767 20893 5776 20927
rect 5724 20884 5776 20893
rect 6368 20884 6420 20936
rect 14372 20927 14424 20936
rect 5448 20859 5500 20868
rect 5448 20825 5457 20859
rect 5457 20825 5491 20859
rect 5491 20825 5500 20859
rect 5448 20816 5500 20825
rect 14372 20893 14381 20927
rect 14381 20893 14415 20927
rect 14415 20893 14424 20927
rect 14372 20884 14424 20893
rect 14648 20884 14700 20936
rect 15660 20927 15712 20936
rect 15660 20893 15669 20927
rect 15669 20893 15703 20927
rect 15703 20893 15712 20927
rect 15660 20884 15712 20893
rect 16212 21020 16264 21072
rect 16856 21020 16908 21072
rect 17684 21063 17736 21072
rect 17684 21029 17693 21063
rect 17693 21029 17727 21063
rect 17727 21029 17736 21063
rect 17684 21020 17736 21029
rect 20812 21097 20821 21131
rect 20821 21097 20855 21131
rect 20855 21097 20864 21131
rect 20812 21088 20864 21097
rect 24400 21088 24452 21140
rect 25136 21088 25188 21140
rect 28632 21088 28684 21140
rect 29092 21088 29144 21140
rect 21824 21020 21876 21072
rect 27344 21020 27396 21072
rect 28448 21020 28500 21072
rect 32404 21088 32456 21140
rect 33692 21088 33744 21140
rect 34520 21088 34572 21140
rect 37188 21131 37240 21140
rect 33048 21063 33100 21072
rect 33048 21029 33057 21063
rect 33057 21029 33091 21063
rect 33091 21029 33100 21063
rect 37188 21097 37197 21131
rect 37197 21097 37231 21131
rect 37231 21097 37240 21131
rect 37188 21088 37240 21097
rect 38016 21088 38068 21140
rect 39304 21131 39356 21140
rect 39304 21097 39313 21131
rect 39313 21097 39347 21131
rect 39347 21097 39356 21131
rect 39304 21088 39356 21097
rect 40960 21131 41012 21140
rect 40960 21097 40969 21131
rect 40969 21097 41003 21131
rect 41003 21097 41012 21131
rect 40960 21088 41012 21097
rect 41696 21088 41748 21140
rect 33048 21020 33100 21029
rect 15844 20952 15896 21004
rect 16580 20927 16632 20936
rect 14096 20791 14148 20800
rect 14096 20757 14105 20791
rect 14105 20757 14139 20791
rect 14139 20757 14148 20791
rect 14096 20748 14148 20757
rect 15016 20816 15068 20868
rect 16580 20893 16589 20927
rect 16589 20893 16623 20927
rect 16623 20893 16632 20927
rect 16580 20884 16632 20893
rect 16856 20927 16908 20936
rect 16856 20893 16864 20927
rect 16864 20893 16898 20927
rect 16898 20893 16908 20927
rect 16856 20884 16908 20893
rect 17132 20884 17184 20936
rect 15568 20748 15620 20800
rect 16304 20816 16356 20868
rect 17592 20816 17644 20868
rect 20720 20952 20772 21004
rect 25964 20952 26016 21004
rect 33692 20995 33744 21004
rect 33692 20961 33701 20995
rect 33701 20961 33735 20995
rect 33735 20961 33744 20995
rect 33692 20952 33744 20961
rect 17960 20927 18012 20936
rect 17960 20893 17969 20927
rect 17969 20893 18003 20927
rect 18003 20893 18012 20927
rect 17960 20884 18012 20893
rect 21088 20927 21140 20936
rect 21088 20893 21097 20927
rect 21097 20893 21131 20927
rect 21131 20893 21140 20927
rect 21088 20884 21140 20893
rect 23480 20884 23532 20936
rect 24584 20927 24636 20936
rect 24584 20893 24593 20927
rect 24593 20893 24627 20927
rect 24627 20893 24636 20927
rect 24584 20884 24636 20893
rect 25044 20884 25096 20936
rect 27068 20927 27120 20936
rect 27068 20893 27077 20927
rect 27077 20893 27111 20927
rect 27111 20893 27120 20927
rect 27068 20884 27120 20893
rect 27620 20884 27672 20936
rect 19984 20816 20036 20868
rect 20812 20859 20864 20868
rect 20812 20825 20821 20859
rect 20821 20825 20855 20859
rect 20855 20825 20864 20859
rect 20812 20816 20864 20825
rect 24860 20816 24912 20868
rect 26700 20859 26752 20868
rect 26700 20825 26709 20859
rect 26709 20825 26743 20859
rect 26743 20825 26752 20859
rect 26700 20816 26752 20825
rect 27896 20927 27948 20936
rect 27896 20893 27905 20927
rect 27905 20893 27939 20927
rect 27939 20893 27948 20927
rect 28724 20927 28776 20936
rect 27896 20884 27948 20893
rect 28724 20893 28733 20927
rect 28733 20893 28767 20927
rect 28767 20893 28776 20927
rect 28724 20884 28776 20893
rect 28816 20884 28868 20936
rect 32312 20884 32364 20936
rect 34796 20884 34848 20936
rect 36360 20952 36412 21004
rect 28172 20816 28224 20868
rect 20076 20791 20128 20800
rect 20076 20757 20085 20791
rect 20085 20757 20119 20791
rect 20119 20757 20128 20791
rect 20076 20748 20128 20757
rect 21272 20791 21324 20800
rect 21272 20757 21281 20791
rect 21281 20757 21315 20791
rect 21315 20757 21324 20791
rect 21272 20748 21324 20757
rect 21824 20791 21876 20800
rect 21824 20757 21833 20791
rect 21833 20757 21867 20791
rect 21867 20757 21876 20791
rect 21824 20748 21876 20757
rect 27620 20748 27672 20800
rect 30288 20748 30340 20800
rect 31392 20748 31444 20800
rect 31576 20816 31628 20868
rect 34888 20859 34940 20868
rect 34888 20825 34897 20859
rect 34897 20825 34931 20859
rect 34931 20825 34940 20859
rect 34888 20816 34940 20825
rect 32128 20748 32180 20800
rect 34060 20748 34112 20800
rect 36268 20884 36320 20936
rect 37188 20952 37240 21004
rect 36912 20927 36964 20936
rect 36912 20893 36921 20927
rect 36921 20893 36955 20927
rect 36955 20893 36964 20927
rect 38752 20952 38804 21004
rect 36912 20884 36964 20893
rect 37924 20927 37976 20936
rect 36820 20816 36872 20868
rect 37924 20893 37933 20927
rect 37933 20893 37967 20927
rect 37967 20893 37976 20927
rect 37924 20884 37976 20893
rect 40316 20927 40368 20936
rect 40316 20893 40325 20927
rect 40325 20893 40359 20927
rect 40359 20893 40368 20927
rect 40868 20927 40920 20936
rect 40316 20884 40368 20893
rect 40868 20893 40877 20927
rect 40877 20893 40911 20927
rect 40911 20893 40920 20927
rect 40868 20884 40920 20893
rect 41512 20927 41564 20936
rect 41512 20893 41521 20927
rect 41521 20893 41555 20927
rect 41555 20893 41564 20927
rect 41512 20884 41564 20893
rect 37832 20816 37884 20868
rect 35348 20748 35400 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 5724 20587 5776 20596
rect 5724 20553 5733 20587
rect 5733 20553 5767 20587
rect 5767 20553 5776 20587
rect 5724 20544 5776 20553
rect 10324 20476 10376 20528
rect 14096 20476 14148 20528
rect 5540 20451 5592 20460
rect 5540 20417 5549 20451
rect 5549 20417 5583 20451
rect 5583 20417 5592 20451
rect 5540 20408 5592 20417
rect 6368 20451 6420 20460
rect 6368 20417 6377 20451
rect 6377 20417 6411 20451
rect 6411 20417 6420 20451
rect 6368 20408 6420 20417
rect 8116 20408 8168 20460
rect 14832 20519 14884 20528
rect 14832 20485 14841 20519
rect 14841 20485 14875 20519
rect 14875 20485 14884 20519
rect 14832 20476 14884 20485
rect 17132 20544 17184 20596
rect 21088 20544 21140 20596
rect 24216 20587 24268 20596
rect 24216 20553 24225 20587
rect 24225 20553 24259 20587
rect 24259 20553 24268 20587
rect 24216 20544 24268 20553
rect 24768 20587 24820 20596
rect 24768 20553 24777 20587
rect 24777 20553 24811 20587
rect 24811 20553 24820 20587
rect 24768 20544 24820 20553
rect 27528 20587 27580 20596
rect 7656 20340 7708 20392
rect 12900 20383 12952 20392
rect 12900 20349 12909 20383
rect 12909 20349 12943 20383
rect 12943 20349 12952 20383
rect 12900 20340 12952 20349
rect 16028 20408 16080 20460
rect 17684 20408 17736 20460
rect 20076 20476 20128 20528
rect 25044 20476 25096 20528
rect 16120 20340 16172 20392
rect 17592 20340 17644 20392
rect 17960 20340 18012 20392
rect 23940 20408 23992 20460
rect 24124 20451 24176 20460
rect 24124 20417 24133 20451
rect 24133 20417 24167 20451
rect 24167 20417 24176 20451
rect 24124 20408 24176 20417
rect 24308 20451 24360 20460
rect 24308 20417 24317 20451
rect 24317 20417 24351 20451
rect 24351 20417 24360 20451
rect 24308 20408 24360 20417
rect 24860 20408 24912 20460
rect 27528 20553 27537 20587
rect 27537 20553 27571 20587
rect 27571 20553 27580 20587
rect 27528 20544 27580 20553
rect 14740 20272 14792 20324
rect 16580 20272 16632 20324
rect 1400 20204 1452 20256
rect 15108 20204 15160 20256
rect 15844 20247 15896 20256
rect 15844 20213 15853 20247
rect 15853 20213 15887 20247
rect 15887 20213 15896 20247
rect 15844 20204 15896 20213
rect 17224 20204 17276 20256
rect 18880 20247 18932 20256
rect 18880 20213 18889 20247
rect 18889 20213 18923 20247
rect 18923 20213 18932 20247
rect 18880 20204 18932 20213
rect 19340 20340 19392 20392
rect 26700 20408 26752 20460
rect 27620 20476 27672 20528
rect 29644 20544 29696 20596
rect 30012 20587 30064 20596
rect 30012 20553 30021 20587
rect 30021 20553 30055 20587
rect 30055 20553 30064 20587
rect 30012 20544 30064 20553
rect 31576 20587 31628 20596
rect 31576 20553 31585 20587
rect 31585 20553 31619 20587
rect 31619 20553 31628 20587
rect 31576 20544 31628 20553
rect 32128 20587 32180 20596
rect 32128 20553 32137 20587
rect 32137 20553 32171 20587
rect 32171 20553 32180 20587
rect 32128 20544 32180 20553
rect 32220 20544 32272 20596
rect 34888 20544 34940 20596
rect 28172 20451 28224 20460
rect 28172 20417 28181 20451
rect 28181 20417 28215 20451
rect 28215 20417 28224 20451
rect 28172 20408 28224 20417
rect 24860 20272 24912 20324
rect 27252 20340 27304 20392
rect 28724 20408 28776 20460
rect 31852 20476 31904 20528
rect 25780 20272 25832 20324
rect 27896 20272 27948 20324
rect 31392 20451 31444 20460
rect 31392 20417 31401 20451
rect 31401 20417 31435 20451
rect 31435 20417 31444 20451
rect 31392 20408 31444 20417
rect 33048 20476 33100 20528
rect 32588 20451 32640 20460
rect 32588 20417 32597 20451
rect 32597 20417 32631 20451
rect 32631 20417 32640 20451
rect 32588 20408 32640 20417
rect 34060 20451 34112 20460
rect 30196 20340 30248 20392
rect 30288 20340 30340 20392
rect 34060 20417 34069 20451
rect 34069 20417 34103 20451
rect 34103 20417 34112 20451
rect 34060 20408 34112 20417
rect 33876 20272 33928 20324
rect 19984 20204 20036 20256
rect 25228 20247 25280 20256
rect 25228 20213 25237 20247
rect 25237 20213 25271 20247
rect 25271 20213 25280 20247
rect 25228 20204 25280 20213
rect 26332 20204 26384 20256
rect 27160 20204 27212 20256
rect 28540 20247 28592 20256
rect 28540 20213 28549 20247
rect 28549 20213 28583 20247
rect 28583 20213 28592 20247
rect 28540 20204 28592 20213
rect 29552 20247 29604 20256
rect 29552 20213 29561 20247
rect 29561 20213 29595 20247
rect 29595 20213 29604 20247
rect 29552 20204 29604 20213
rect 30380 20204 30432 20256
rect 32220 20204 32272 20256
rect 36268 20519 36320 20528
rect 36268 20485 36277 20519
rect 36277 20485 36311 20519
rect 36311 20485 36320 20519
rect 36268 20476 36320 20485
rect 37188 20476 37240 20528
rect 36176 20408 36228 20460
rect 36912 20408 36964 20460
rect 37096 20408 37148 20460
rect 37832 20408 37884 20460
rect 40316 20544 40368 20596
rect 35900 20340 35952 20392
rect 36176 20272 36228 20324
rect 37280 20204 37332 20256
rect 37556 20340 37608 20392
rect 40224 20204 40276 20256
rect 41696 20247 41748 20256
rect 41696 20213 41705 20247
rect 41705 20213 41739 20247
rect 41739 20213 41748 20247
rect 41696 20204 41748 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 5448 20000 5500 20052
rect 39120 20000 39172 20052
rect 40868 20000 40920 20052
rect 16672 19932 16724 19984
rect 17776 19932 17828 19984
rect 18788 19932 18840 19984
rect 20720 19975 20772 19984
rect 1400 19907 1452 19916
rect 1400 19873 1409 19907
rect 1409 19873 1443 19907
rect 1443 19873 1452 19907
rect 1400 19864 1452 19873
rect 1860 19907 1912 19916
rect 1860 19873 1869 19907
rect 1869 19873 1903 19907
rect 1903 19873 1912 19907
rect 1860 19864 1912 19873
rect 6736 19907 6788 19916
rect 6736 19873 6745 19907
rect 6745 19873 6779 19907
rect 6779 19873 6788 19907
rect 6736 19864 6788 19873
rect 11612 19907 11664 19916
rect 11612 19873 11621 19907
rect 11621 19873 11655 19907
rect 11655 19873 11664 19907
rect 11612 19864 11664 19873
rect 13360 19864 13412 19916
rect 16580 19864 16632 19916
rect 20720 19941 20729 19975
rect 20729 19941 20763 19975
rect 20763 19941 20772 19975
rect 20720 19932 20772 19941
rect 24124 19932 24176 19984
rect 26884 19932 26936 19984
rect 6368 19796 6420 19848
rect 10324 19839 10376 19848
rect 10324 19805 10333 19839
rect 10333 19805 10367 19839
rect 10367 19805 10376 19839
rect 10324 19796 10376 19805
rect 11244 19796 11296 19848
rect 15844 19796 15896 19848
rect 16028 19839 16080 19848
rect 16028 19805 16037 19839
rect 16037 19805 16071 19839
rect 16071 19805 16080 19839
rect 16028 19796 16080 19805
rect 19340 19839 19392 19848
rect 19340 19805 19349 19839
rect 19349 19805 19383 19839
rect 19383 19805 19392 19839
rect 19340 19796 19392 19805
rect 2044 19728 2096 19780
rect 19432 19728 19484 19780
rect 2596 19660 2648 19712
rect 11612 19660 11664 19712
rect 19340 19660 19392 19712
rect 22008 19728 22060 19780
rect 22744 19728 22796 19780
rect 21640 19660 21692 19712
rect 25504 19907 25556 19916
rect 25504 19873 25513 19907
rect 25513 19873 25547 19907
rect 25547 19873 25556 19907
rect 25504 19864 25556 19873
rect 25780 19907 25832 19916
rect 25780 19873 25789 19907
rect 25789 19873 25823 19907
rect 25823 19873 25832 19907
rect 25780 19864 25832 19873
rect 26332 19864 26384 19916
rect 28264 19932 28316 19984
rect 30656 19932 30708 19984
rect 32588 19932 32640 19984
rect 37280 19932 37332 19984
rect 27344 19907 27396 19916
rect 27344 19873 27353 19907
rect 27353 19873 27387 19907
rect 27387 19873 27396 19907
rect 27344 19864 27396 19873
rect 24584 19796 24636 19848
rect 24768 19839 24820 19848
rect 24768 19805 24777 19839
rect 24777 19805 24811 19839
rect 24811 19805 24820 19839
rect 24768 19796 24820 19805
rect 24952 19839 25004 19848
rect 24952 19805 24961 19839
rect 24961 19805 24995 19839
rect 24995 19805 25004 19839
rect 24952 19796 25004 19805
rect 25228 19796 25280 19848
rect 27252 19796 27304 19848
rect 28356 19864 28408 19916
rect 34704 19864 34756 19916
rect 37096 19864 37148 19916
rect 30104 19839 30156 19848
rect 30104 19805 30113 19839
rect 30113 19805 30147 19839
rect 30147 19805 30156 19839
rect 30104 19796 30156 19805
rect 30196 19839 30248 19848
rect 30196 19805 30205 19839
rect 30205 19805 30239 19839
rect 30239 19805 30248 19839
rect 30380 19839 30432 19848
rect 30196 19796 30248 19805
rect 30380 19805 30389 19839
rect 30389 19805 30423 19839
rect 30423 19805 30432 19839
rect 30380 19796 30432 19805
rect 32404 19796 32456 19848
rect 33600 19796 33652 19848
rect 36820 19839 36872 19848
rect 36820 19805 36829 19839
rect 36829 19805 36863 19839
rect 36863 19805 36872 19839
rect 36820 19796 36872 19805
rect 37188 19796 37240 19848
rect 37924 19796 37976 19848
rect 38476 19839 38528 19848
rect 38476 19805 38485 19839
rect 38485 19805 38519 19839
rect 38519 19805 38528 19839
rect 38476 19796 38528 19805
rect 41696 19864 41748 19916
rect 40316 19839 40368 19848
rect 40316 19805 40325 19839
rect 40325 19805 40359 19839
rect 40359 19805 40368 19839
rect 40316 19796 40368 19805
rect 23940 19728 23992 19780
rect 35900 19728 35952 19780
rect 37096 19728 37148 19780
rect 42156 19771 42208 19780
rect 42156 19737 42165 19771
rect 42165 19737 42199 19771
rect 42199 19737 42208 19771
rect 42156 19728 42208 19737
rect 24584 19660 24636 19712
rect 32496 19660 32548 19712
rect 34980 19660 35032 19712
rect 36636 19703 36688 19712
rect 36636 19669 36645 19703
rect 36645 19669 36679 19703
rect 36679 19669 36688 19703
rect 36636 19660 36688 19669
rect 38016 19703 38068 19712
rect 38016 19669 38025 19703
rect 38025 19669 38059 19703
rect 38059 19669 38068 19703
rect 38016 19660 38068 19669
rect 40408 19660 40460 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 2044 19499 2096 19508
rect 2044 19465 2053 19499
rect 2053 19465 2087 19499
rect 2087 19465 2096 19499
rect 2044 19456 2096 19465
rect 8944 19456 8996 19508
rect 2136 19363 2188 19372
rect 2136 19329 2145 19363
rect 2145 19329 2179 19363
rect 2179 19329 2188 19363
rect 2136 19320 2188 19329
rect 12164 19388 12216 19440
rect 15016 19388 15068 19440
rect 16212 19456 16264 19508
rect 19340 19456 19392 19508
rect 24308 19499 24360 19508
rect 16304 19388 16356 19440
rect 10692 19320 10744 19372
rect 11244 19320 11296 19372
rect 12900 19363 12952 19372
rect 12900 19329 12909 19363
rect 12909 19329 12943 19363
rect 12943 19329 12952 19363
rect 12900 19320 12952 19329
rect 15660 19363 15712 19372
rect 15660 19329 15669 19363
rect 15669 19329 15703 19363
rect 15703 19329 15712 19363
rect 15660 19320 15712 19329
rect 16120 19363 16172 19372
rect 16120 19329 16129 19363
rect 16129 19329 16163 19363
rect 16163 19329 16172 19363
rect 16120 19320 16172 19329
rect 15844 19252 15896 19304
rect 17776 19363 17828 19372
rect 17776 19329 17792 19363
rect 17792 19329 17826 19363
rect 17826 19329 17828 19363
rect 17776 19320 17828 19329
rect 18052 19363 18104 19372
rect 18052 19329 18086 19363
rect 18086 19329 18104 19363
rect 18052 19320 18104 19329
rect 18880 19320 18932 19372
rect 22008 19320 22060 19372
rect 22468 19320 22520 19372
rect 24308 19465 24317 19499
rect 24317 19465 24351 19499
rect 24351 19465 24360 19499
rect 24308 19456 24360 19465
rect 24952 19456 25004 19508
rect 25228 19499 25280 19508
rect 25228 19465 25237 19499
rect 25237 19465 25271 19499
rect 25271 19465 25280 19499
rect 25228 19456 25280 19465
rect 27068 19499 27120 19508
rect 27068 19465 27077 19499
rect 27077 19465 27111 19499
rect 27111 19465 27120 19499
rect 27068 19456 27120 19465
rect 32404 19499 32456 19508
rect 32404 19465 32413 19499
rect 32413 19465 32447 19499
rect 32447 19465 32456 19499
rect 32404 19456 32456 19465
rect 37188 19456 37240 19508
rect 26884 19388 26936 19440
rect 32220 19388 32272 19440
rect 33600 19388 33652 19440
rect 40224 19431 40276 19440
rect 40224 19397 40233 19431
rect 40233 19397 40267 19431
rect 40267 19397 40276 19431
rect 40224 19388 40276 19397
rect 24492 19363 24544 19372
rect 24492 19329 24501 19363
rect 24501 19329 24535 19363
rect 24535 19329 24544 19363
rect 24492 19320 24544 19329
rect 24768 19320 24820 19372
rect 25504 19320 25556 19372
rect 24584 19295 24636 19304
rect 14280 19159 14332 19168
rect 14280 19125 14289 19159
rect 14289 19125 14323 19159
rect 14323 19125 14332 19159
rect 14280 19116 14332 19125
rect 16948 19116 17000 19168
rect 24584 19261 24593 19295
rect 24593 19261 24627 19295
rect 24627 19261 24636 19295
rect 27344 19320 27396 19372
rect 28724 19363 28776 19372
rect 28724 19329 28733 19363
rect 28733 19329 28767 19363
rect 28767 19329 28776 19363
rect 28724 19320 28776 19329
rect 29552 19320 29604 19372
rect 29920 19320 29972 19372
rect 24584 19252 24636 19261
rect 30472 19320 30524 19372
rect 32588 19363 32640 19372
rect 32588 19329 32597 19363
rect 32597 19329 32631 19363
rect 32631 19329 32640 19363
rect 32588 19320 32640 19329
rect 35348 19320 35400 19372
rect 30104 19295 30156 19304
rect 30104 19261 30113 19295
rect 30113 19261 30147 19295
rect 30147 19261 30156 19295
rect 32128 19295 32180 19304
rect 30104 19252 30156 19261
rect 32128 19261 32137 19295
rect 32137 19261 32171 19295
rect 32171 19261 32180 19295
rect 32128 19252 32180 19261
rect 34980 19295 35032 19304
rect 34980 19261 34989 19295
rect 34989 19261 35023 19295
rect 35023 19261 35032 19295
rect 34980 19252 35032 19261
rect 38476 19320 38528 19372
rect 40040 19363 40092 19372
rect 40040 19329 40049 19363
rect 40049 19329 40083 19363
rect 40083 19329 40092 19363
rect 40040 19320 40092 19329
rect 41236 19295 41288 19304
rect 24308 19184 24360 19236
rect 24676 19184 24728 19236
rect 26332 19184 26384 19236
rect 29000 19184 29052 19236
rect 41236 19261 41245 19295
rect 41245 19261 41279 19295
rect 41279 19261 41288 19295
rect 41236 19252 41288 19261
rect 40316 19184 40368 19236
rect 18696 19116 18748 19168
rect 24860 19116 24912 19168
rect 28816 19159 28868 19168
rect 28816 19125 28825 19159
rect 28825 19125 28859 19159
rect 28859 19125 28868 19159
rect 28816 19116 28868 19125
rect 29828 19116 29880 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 18052 18912 18104 18964
rect 19432 18912 19484 18964
rect 20812 18912 20864 18964
rect 26240 18912 26292 18964
rect 33600 18955 33652 18964
rect 33600 18921 33609 18955
rect 33609 18921 33643 18955
rect 33643 18921 33652 18955
rect 33600 18912 33652 18921
rect 14648 18844 14700 18896
rect 15016 18844 15068 18896
rect 20076 18844 20128 18896
rect 22744 18887 22796 18896
rect 22744 18853 22753 18887
rect 22753 18853 22787 18887
rect 22787 18853 22796 18887
rect 22744 18844 22796 18853
rect 25504 18844 25556 18896
rect 14280 18776 14332 18828
rect 14924 18776 14976 18828
rect 16120 18776 16172 18828
rect 16304 18776 16356 18828
rect 11244 18708 11296 18760
rect 15016 18708 15068 18760
rect 16948 18751 17000 18760
rect 16948 18717 16957 18751
rect 16957 18717 16991 18751
rect 16991 18717 17000 18751
rect 16948 18708 17000 18717
rect 17408 18751 17460 18760
rect 17408 18717 17417 18751
rect 17417 18717 17451 18751
rect 17451 18717 17460 18751
rect 17408 18708 17460 18717
rect 28816 18776 28868 18828
rect 30012 18776 30064 18828
rect 40408 18819 40460 18828
rect 40408 18785 40417 18819
rect 40417 18785 40451 18819
rect 40451 18785 40460 18819
rect 40408 18776 40460 18785
rect 20904 18751 20956 18760
rect 20904 18717 20913 18751
rect 20913 18717 20947 18751
rect 20947 18717 20956 18751
rect 20904 18708 20956 18717
rect 22008 18708 22060 18760
rect 22284 18708 22336 18760
rect 29000 18708 29052 18760
rect 29828 18751 29880 18760
rect 29828 18717 29837 18751
rect 29837 18717 29871 18751
rect 29871 18717 29880 18751
rect 29828 18708 29880 18717
rect 30472 18708 30524 18760
rect 11704 18640 11756 18692
rect 13636 18640 13688 18692
rect 16672 18683 16724 18692
rect 16672 18649 16681 18683
rect 16681 18649 16715 18683
rect 16715 18649 16724 18683
rect 16672 18640 16724 18649
rect 17592 18683 17644 18692
rect 17592 18649 17601 18683
rect 17601 18649 17635 18683
rect 17635 18649 17644 18683
rect 17592 18640 17644 18649
rect 18880 18640 18932 18692
rect 20812 18640 20864 18692
rect 20996 18640 21048 18692
rect 23572 18640 23624 18692
rect 29920 18640 29972 18692
rect 30012 18640 30064 18692
rect 32312 18708 32364 18760
rect 32496 18751 32548 18760
rect 32496 18717 32530 18751
rect 32530 18717 32548 18751
rect 32496 18708 32548 18717
rect 38936 18751 38988 18760
rect 38936 18717 38945 18751
rect 38945 18717 38979 18751
rect 38979 18717 38988 18751
rect 38936 18708 38988 18717
rect 39028 18751 39080 18760
rect 39028 18717 39037 18751
rect 39037 18717 39071 18751
rect 39071 18717 39080 18751
rect 39028 18708 39080 18717
rect 39580 18708 39632 18760
rect 42064 18683 42116 18692
rect 42064 18649 42073 18683
rect 42073 18649 42107 18683
rect 42107 18649 42116 18683
rect 42064 18640 42116 18649
rect 15936 18572 15988 18624
rect 19984 18572 20036 18624
rect 24492 18572 24544 18624
rect 29092 18572 29144 18624
rect 29644 18572 29696 18624
rect 30748 18615 30800 18624
rect 30748 18581 30757 18615
rect 30757 18581 30791 18615
rect 30791 18581 30800 18615
rect 30748 18572 30800 18581
rect 39396 18572 39448 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 16212 18368 16264 18420
rect 22284 18411 22336 18420
rect 12900 18300 12952 18352
rect 13728 18232 13780 18284
rect 11520 18207 11572 18216
rect 11520 18173 11529 18207
rect 11529 18173 11563 18207
rect 11563 18173 11572 18207
rect 11520 18164 11572 18173
rect 15844 18275 15896 18284
rect 15844 18241 15856 18275
rect 15856 18241 15890 18275
rect 15890 18241 15896 18275
rect 15844 18232 15896 18241
rect 15936 18275 15988 18284
rect 15936 18241 15945 18275
rect 15945 18241 15979 18275
rect 15979 18241 15988 18275
rect 15936 18232 15988 18241
rect 16580 18232 16632 18284
rect 14924 18207 14976 18216
rect 14924 18173 14933 18207
rect 14933 18173 14967 18207
rect 14967 18173 14976 18207
rect 14924 18164 14976 18173
rect 15016 18207 15068 18216
rect 15016 18173 15025 18207
rect 15025 18173 15059 18207
rect 15059 18173 15068 18207
rect 16948 18232 17000 18284
rect 22284 18377 22293 18411
rect 22293 18377 22327 18411
rect 22327 18377 22336 18411
rect 22284 18368 22336 18377
rect 28724 18368 28776 18420
rect 18052 18232 18104 18284
rect 18696 18232 18748 18284
rect 18880 18275 18932 18284
rect 18880 18241 18889 18275
rect 18889 18241 18923 18275
rect 18923 18241 18932 18275
rect 18880 18232 18932 18241
rect 19984 18275 20036 18284
rect 19984 18241 19993 18275
rect 19993 18241 20027 18275
rect 20027 18241 20036 18275
rect 19984 18232 20036 18241
rect 28632 18232 28684 18284
rect 29092 18300 29144 18352
rect 29460 18343 29512 18352
rect 29460 18309 29461 18343
rect 29461 18309 29495 18343
rect 29495 18309 29512 18343
rect 29460 18300 29512 18309
rect 30012 18368 30064 18420
rect 38936 18411 38988 18420
rect 38936 18377 38945 18411
rect 38945 18377 38979 18411
rect 38979 18377 38988 18411
rect 38936 18368 38988 18377
rect 39580 18411 39632 18420
rect 39580 18377 39589 18411
rect 39589 18377 39623 18411
rect 39623 18377 39632 18411
rect 39580 18368 39632 18377
rect 30104 18300 30156 18352
rect 32312 18300 32364 18352
rect 15016 18164 15068 18173
rect 21640 18164 21692 18216
rect 30656 18275 30708 18284
rect 30656 18241 30665 18275
rect 30665 18241 30699 18275
rect 30699 18241 30708 18275
rect 38016 18300 38068 18352
rect 30656 18232 30708 18241
rect 30748 18164 30800 18216
rect 36360 18232 36412 18284
rect 37556 18275 37608 18284
rect 37556 18241 37565 18275
rect 37565 18241 37599 18275
rect 37599 18241 37608 18275
rect 37556 18232 37608 18241
rect 39396 18275 39448 18284
rect 39396 18241 39405 18275
rect 39405 18241 39439 18275
rect 39439 18241 39448 18275
rect 39396 18232 39448 18241
rect 41328 18207 41380 18216
rect 41328 18173 41337 18207
rect 41337 18173 41371 18207
rect 41371 18173 41380 18207
rect 41328 18164 41380 18173
rect 41696 18207 41748 18216
rect 41696 18173 41705 18207
rect 41705 18173 41739 18207
rect 41739 18173 41748 18207
rect 41696 18164 41748 18173
rect 41880 18207 41932 18216
rect 41880 18173 41889 18207
rect 41889 18173 41923 18207
rect 41923 18173 41932 18207
rect 41880 18164 41932 18173
rect 15200 18096 15252 18148
rect 15660 18096 15712 18148
rect 20076 18096 20128 18148
rect 32128 18096 32180 18148
rect 13544 18028 13596 18080
rect 14740 18028 14792 18080
rect 15108 18028 15160 18080
rect 16488 18028 16540 18080
rect 20168 18071 20220 18080
rect 20168 18037 20177 18071
rect 20177 18037 20211 18071
rect 20211 18037 20220 18071
rect 20168 18028 20220 18037
rect 29736 18071 29788 18080
rect 29736 18037 29745 18071
rect 29745 18037 29779 18071
rect 29779 18037 29788 18071
rect 29736 18028 29788 18037
rect 31024 18071 31076 18080
rect 31024 18037 31033 18071
rect 31033 18037 31067 18071
rect 31067 18037 31076 18071
rect 31024 18028 31076 18037
rect 34796 18071 34848 18080
rect 34796 18037 34805 18071
rect 34805 18037 34839 18071
rect 34839 18037 34848 18071
rect 34796 18028 34848 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 13728 17824 13780 17876
rect 14464 17824 14516 17876
rect 14372 17756 14424 17808
rect 14924 17824 14976 17876
rect 15384 17867 15436 17876
rect 15384 17833 15393 17867
rect 15393 17833 15427 17867
rect 15427 17833 15436 17867
rect 15384 17824 15436 17833
rect 16120 17824 16172 17876
rect 17592 17824 17644 17876
rect 26240 17824 26292 17876
rect 30012 17824 30064 17876
rect 40040 17824 40092 17876
rect 41696 17824 41748 17876
rect 41880 17824 41932 17876
rect 1952 17620 2004 17672
rect 11152 17620 11204 17672
rect 11244 17620 11296 17672
rect 13268 17663 13320 17672
rect 13268 17629 13277 17663
rect 13277 17629 13311 17663
rect 13311 17629 13320 17663
rect 13268 17620 13320 17629
rect 14096 17620 14148 17672
rect 14648 17688 14700 17740
rect 15936 17756 15988 17808
rect 29460 17756 29512 17808
rect 14740 17663 14792 17672
rect 14740 17629 14749 17663
rect 14749 17629 14783 17663
rect 14783 17629 14792 17663
rect 14740 17620 14792 17629
rect 13544 17595 13596 17604
rect 13544 17561 13553 17595
rect 13553 17561 13587 17595
rect 13587 17561 13596 17595
rect 13544 17552 13596 17561
rect 13728 17552 13780 17604
rect 14464 17595 14516 17604
rect 14464 17561 14473 17595
rect 14473 17561 14507 17595
rect 14507 17561 14516 17595
rect 14464 17552 14516 17561
rect 14556 17595 14608 17604
rect 14556 17561 14591 17595
rect 14591 17561 14608 17595
rect 14556 17552 14608 17561
rect 15292 17552 15344 17604
rect 15752 17552 15804 17604
rect 16488 17595 16540 17604
rect 16488 17561 16497 17595
rect 16497 17561 16531 17595
rect 16531 17561 16540 17595
rect 16488 17552 16540 17561
rect 16672 17595 16724 17604
rect 16672 17561 16697 17595
rect 16697 17561 16724 17595
rect 17960 17688 18012 17740
rect 17868 17663 17920 17672
rect 17868 17629 17877 17663
rect 17877 17629 17911 17663
rect 17911 17629 17920 17663
rect 18972 17688 19024 17740
rect 29368 17688 29420 17740
rect 36360 17731 36412 17740
rect 36360 17697 36369 17731
rect 36369 17697 36403 17731
rect 36403 17697 36412 17731
rect 36360 17688 36412 17697
rect 39028 17688 39080 17740
rect 17868 17620 17920 17629
rect 18328 17620 18380 17672
rect 20076 17620 20128 17672
rect 20904 17620 20956 17672
rect 27804 17620 27856 17672
rect 28724 17663 28776 17672
rect 28724 17629 28742 17663
rect 28742 17629 28776 17663
rect 28724 17620 28776 17629
rect 29920 17620 29972 17672
rect 31024 17620 31076 17672
rect 34796 17663 34848 17672
rect 34796 17629 34805 17663
rect 34805 17629 34839 17663
rect 34839 17629 34848 17663
rect 34796 17620 34848 17629
rect 34980 17663 35032 17672
rect 34980 17629 34989 17663
rect 34989 17629 35023 17663
rect 35023 17629 35032 17663
rect 34980 17620 35032 17629
rect 36636 17663 36688 17672
rect 36636 17629 36670 17663
rect 36670 17629 36688 17663
rect 36636 17620 36688 17629
rect 38476 17663 38528 17672
rect 38476 17629 38485 17663
rect 38485 17629 38519 17663
rect 38519 17629 38528 17663
rect 38476 17620 38528 17629
rect 38752 17663 38804 17672
rect 38752 17629 38761 17663
rect 38761 17629 38795 17663
rect 38795 17629 38804 17663
rect 38752 17620 38804 17629
rect 39764 17620 39816 17672
rect 41144 17620 41196 17672
rect 16672 17552 16724 17561
rect 19984 17552 20036 17604
rect 20168 17552 20220 17604
rect 2136 17484 2188 17536
rect 15384 17484 15436 17536
rect 17132 17484 17184 17536
rect 26884 17595 26936 17604
rect 26884 17561 26902 17595
rect 26902 17561 26936 17595
rect 30012 17595 30064 17604
rect 26884 17552 26936 17561
rect 23664 17484 23716 17536
rect 23848 17527 23900 17536
rect 23848 17493 23857 17527
rect 23857 17493 23891 17527
rect 23891 17493 23900 17527
rect 23848 17484 23900 17493
rect 28632 17484 28684 17536
rect 30012 17561 30021 17595
rect 30021 17561 30055 17595
rect 30055 17561 30064 17595
rect 30012 17552 30064 17561
rect 29000 17484 29052 17536
rect 30104 17527 30156 17536
rect 30104 17493 30113 17527
rect 30113 17493 30147 17527
rect 30147 17493 30156 17527
rect 30104 17484 30156 17493
rect 32588 17484 32640 17536
rect 34796 17484 34848 17536
rect 37924 17484 37976 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 13360 17280 13412 17332
rect 2136 17255 2188 17264
rect 2136 17221 2145 17255
rect 2145 17221 2179 17255
rect 2179 17221 2188 17255
rect 2136 17212 2188 17221
rect 13728 17255 13780 17264
rect 13728 17221 13737 17255
rect 13737 17221 13771 17255
rect 13771 17221 13780 17255
rect 13728 17212 13780 17221
rect 14096 17280 14148 17332
rect 17960 17280 18012 17332
rect 18972 17323 19024 17332
rect 18972 17289 18981 17323
rect 18981 17289 19015 17323
rect 19015 17289 19024 17323
rect 18972 17280 19024 17289
rect 15200 17255 15252 17264
rect 1952 17187 2004 17196
rect 1952 17153 1961 17187
rect 1961 17153 1995 17187
rect 1995 17153 2004 17187
rect 1952 17144 2004 17153
rect 11520 17187 11572 17196
rect 11520 17153 11529 17187
rect 11529 17153 11563 17187
rect 11563 17153 11572 17187
rect 11520 17144 11572 17153
rect 13452 17144 13504 17196
rect 13636 17187 13688 17196
rect 13636 17153 13645 17187
rect 13645 17153 13679 17187
rect 13679 17153 13688 17187
rect 15200 17221 15209 17255
rect 15209 17221 15243 17255
rect 15243 17221 15252 17255
rect 15200 17212 15252 17221
rect 17868 17212 17920 17264
rect 39764 17280 39816 17332
rect 13636 17144 13688 17153
rect 2780 17119 2832 17128
rect 2780 17085 2789 17119
rect 2789 17085 2823 17119
rect 2823 17085 2832 17119
rect 2780 17076 2832 17085
rect 14372 17144 14424 17196
rect 13820 16940 13872 16992
rect 14280 17076 14332 17128
rect 14924 17144 14976 17196
rect 15476 17187 15528 17196
rect 15476 17153 15485 17187
rect 15485 17153 15519 17187
rect 15519 17153 15528 17187
rect 15476 17144 15528 17153
rect 14740 17076 14792 17128
rect 15752 17144 15804 17196
rect 17224 17187 17276 17196
rect 16948 17119 17000 17128
rect 16948 17085 16957 17119
rect 16957 17085 16991 17119
rect 16991 17085 17000 17119
rect 16948 17076 17000 17085
rect 17224 17153 17233 17187
rect 17233 17153 17267 17187
rect 17267 17153 17276 17187
rect 17224 17144 17276 17153
rect 18236 17144 18288 17196
rect 18972 17144 19024 17196
rect 14372 17008 14424 17060
rect 29460 17212 29512 17264
rect 20076 17144 20128 17196
rect 21364 17144 21416 17196
rect 19984 17076 20036 17128
rect 20628 17119 20680 17128
rect 20628 17085 20637 17119
rect 20637 17085 20671 17119
rect 20671 17085 20680 17119
rect 20628 17076 20680 17085
rect 24768 17144 24820 17196
rect 25596 17187 25648 17196
rect 25596 17153 25605 17187
rect 25605 17153 25639 17187
rect 25639 17153 25648 17187
rect 25596 17144 25648 17153
rect 29368 17187 29420 17196
rect 29368 17153 29377 17187
rect 29377 17153 29411 17187
rect 29411 17153 29420 17187
rect 29368 17144 29420 17153
rect 34980 17212 35032 17264
rect 22100 17076 22152 17128
rect 26884 17076 26936 17128
rect 34888 17187 34940 17196
rect 34888 17153 34897 17187
rect 34897 17153 34931 17187
rect 34931 17153 34940 17187
rect 38752 17212 38804 17264
rect 34888 17144 34940 17153
rect 37924 17187 37976 17196
rect 37924 17153 37933 17187
rect 37933 17153 37967 17187
rect 37967 17153 37976 17187
rect 37924 17144 37976 17153
rect 14556 16940 14608 16992
rect 15108 16940 15160 16992
rect 16580 16940 16632 16992
rect 16672 16983 16724 16992
rect 16672 16949 16681 16983
rect 16681 16949 16715 16983
rect 16715 16949 16724 16983
rect 17132 16983 17184 16992
rect 16672 16940 16724 16949
rect 17132 16949 17141 16983
rect 17141 16949 17175 16983
rect 17175 16949 17184 16983
rect 17132 16940 17184 16949
rect 18052 16983 18104 16992
rect 18052 16949 18061 16983
rect 18061 16949 18095 16983
rect 18095 16949 18104 16983
rect 18052 16940 18104 16949
rect 18420 16983 18472 16992
rect 18420 16949 18429 16983
rect 18429 16949 18463 16983
rect 18463 16949 18472 16983
rect 18420 16940 18472 16949
rect 19248 16940 19300 16992
rect 22192 16940 22244 16992
rect 24492 16940 24544 16992
rect 30748 16983 30800 16992
rect 30748 16949 30757 16983
rect 30757 16949 30791 16983
rect 30791 16949 30800 16983
rect 30748 16940 30800 16949
rect 34612 16983 34664 16992
rect 34612 16949 34621 16983
rect 34621 16949 34655 16983
rect 34655 16949 34664 16983
rect 34612 16940 34664 16949
rect 37648 16983 37700 16992
rect 37648 16949 37657 16983
rect 37657 16949 37691 16983
rect 37691 16949 37700 16983
rect 37648 16940 37700 16949
rect 42156 16940 42208 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 7656 16736 7708 16788
rect 14372 16736 14424 16788
rect 14464 16736 14516 16788
rect 14924 16736 14976 16788
rect 15108 16779 15160 16788
rect 15108 16745 15117 16779
rect 15117 16745 15151 16779
rect 15151 16745 15160 16779
rect 15108 16736 15160 16745
rect 16488 16736 16540 16788
rect 13268 16668 13320 16720
rect 1860 16643 1912 16652
rect 1860 16609 1869 16643
rect 1869 16609 1903 16643
rect 1903 16609 1912 16643
rect 1860 16600 1912 16609
rect 13820 16600 13872 16652
rect 14464 16643 14516 16652
rect 14464 16609 14473 16643
rect 14473 16609 14507 16643
rect 14507 16609 14516 16643
rect 14464 16600 14516 16609
rect 15476 16668 15528 16720
rect 1400 16575 1452 16584
rect 1400 16541 1409 16575
rect 1409 16541 1443 16575
rect 1443 16541 1452 16575
rect 1400 16532 1452 16541
rect 13360 16532 13412 16584
rect 14280 16575 14332 16584
rect 14280 16541 14289 16575
rect 14289 16541 14323 16575
rect 14323 16541 14332 16575
rect 14280 16532 14332 16541
rect 15108 16575 15160 16584
rect 15108 16541 15117 16575
rect 15117 16541 15151 16575
rect 15151 16541 15160 16575
rect 17960 16668 18012 16720
rect 18420 16736 18472 16788
rect 21364 16779 21416 16788
rect 21364 16745 21373 16779
rect 21373 16745 21407 16779
rect 21407 16745 21416 16779
rect 21364 16736 21416 16745
rect 23848 16736 23900 16788
rect 24768 16736 24820 16788
rect 27712 16736 27764 16788
rect 27804 16736 27856 16788
rect 29368 16736 29420 16788
rect 16948 16600 17000 16652
rect 17684 16643 17736 16652
rect 17684 16609 17693 16643
rect 17693 16609 17727 16643
rect 17727 16609 17736 16643
rect 17684 16600 17736 16609
rect 15108 16532 15160 16541
rect 15936 16532 15988 16584
rect 16580 16532 16632 16584
rect 18052 16532 18104 16584
rect 19248 16575 19300 16584
rect 19248 16541 19257 16575
rect 19257 16541 19291 16575
rect 19291 16541 19300 16575
rect 19248 16532 19300 16541
rect 2136 16464 2188 16516
rect 17040 16507 17092 16516
rect 17040 16473 17049 16507
rect 17049 16473 17083 16507
rect 17083 16473 17092 16507
rect 17040 16464 17092 16473
rect 21180 16600 21232 16652
rect 20076 16532 20128 16584
rect 26240 16668 26292 16720
rect 22192 16643 22244 16652
rect 22192 16609 22201 16643
rect 22201 16609 22235 16643
rect 22235 16609 22244 16643
rect 22192 16600 22244 16609
rect 24492 16643 24544 16652
rect 24492 16609 24501 16643
rect 24501 16609 24535 16643
rect 24535 16609 24544 16643
rect 24492 16600 24544 16609
rect 23664 16532 23716 16584
rect 24860 16600 24912 16652
rect 25596 16575 25648 16584
rect 25596 16541 25605 16575
rect 25605 16541 25639 16575
rect 25639 16541 25648 16575
rect 25596 16532 25648 16541
rect 23756 16464 23808 16516
rect 24768 16464 24820 16516
rect 13544 16396 13596 16448
rect 15476 16439 15528 16448
rect 15476 16405 15485 16439
rect 15485 16405 15519 16439
rect 15519 16405 15528 16439
rect 15476 16396 15528 16405
rect 15752 16396 15804 16448
rect 21732 16396 21784 16448
rect 24676 16396 24728 16448
rect 25136 16396 25188 16448
rect 32772 16668 32824 16720
rect 33324 16668 33376 16720
rect 34796 16600 34848 16652
rect 41696 16643 41748 16652
rect 30104 16532 30156 16584
rect 30748 16532 30800 16584
rect 31024 16575 31076 16584
rect 31024 16541 31033 16575
rect 31033 16541 31067 16575
rect 31067 16541 31076 16575
rect 31024 16532 31076 16541
rect 31116 16464 31168 16516
rect 32588 16575 32640 16584
rect 32588 16541 32597 16575
rect 32597 16541 32631 16575
rect 32631 16541 32640 16575
rect 32864 16575 32916 16584
rect 32588 16532 32640 16541
rect 32864 16541 32872 16575
rect 32872 16541 32906 16575
rect 32906 16541 32916 16575
rect 32864 16532 32916 16541
rect 32956 16575 33008 16584
rect 32956 16541 32965 16575
rect 32965 16541 32999 16575
rect 32999 16541 33008 16575
rect 41696 16609 41705 16643
rect 41705 16609 41739 16643
rect 41739 16609 41748 16643
rect 41696 16600 41748 16609
rect 42156 16643 42208 16652
rect 42156 16609 42165 16643
rect 42165 16609 42199 16643
rect 42199 16609 42208 16643
rect 42156 16600 42208 16609
rect 32956 16532 33008 16541
rect 37648 16575 37700 16584
rect 32772 16464 32824 16516
rect 34612 16464 34664 16516
rect 37648 16541 37657 16575
rect 37657 16541 37691 16575
rect 37691 16541 37700 16575
rect 37648 16532 37700 16541
rect 35348 16464 35400 16516
rect 41420 16464 41472 16516
rect 26148 16396 26200 16448
rect 31024 16396 31076 16448
rect 32312 16439 32364 16448
rect 32312 16405 32321 16439
rect 32321 16405 32355 16439
rect 32355 16405 32364 16439
rect 32312 16396 32364 16405
rect 32588 16396 32640 16448
rect 34704 16396 34756 16448
rect 34796 16396 34848 16448
rect 37280 16396 37332 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 2136 16235 2188 16244
rect 2136 16201 2145 16235
rect 2145 16201 2179 16235
rect 2179 16201 2188 16235
rect 2136 16192 2188 16201
rect 1400 16099 1452 16108
rect 1400 16065 1409 16099
rect 1409 16065 1443 16099
rect 1443 16065 1452 16099
rect 1400 16056 1452 16065
rect 7104 16056 7156 16108
rect 13360 16124 13412 16176
rect 14372 16124 14424 16176
rect 14280 16056 14332 16108
rect 13268 15988 13320 16040
rect 14372 15988 14424 16040
rect 15476 16192 15528 16244
rect 18144 16192 18196 16244
rect 20720 16235 20772 16244
rect 20720 16201 20729 16235
rect 20729 16201 20763 16235
rect 20763 16201 20772 16235
rect 20720 16192 20772 16201
rect 41420 16235 41472 16244
rect 15752 16099 15804 16108
rect 15752 16065 15761 16099
rect 15761 16065 15795 16099
rect 15795 16065 15804 16099
rect 15752 16056 15804 16065
rect 17684 15988 17736 16040
rect 14464 15920 14516 15972
rect 21180 16124 21232 16176
rect 17960 16099 18012 16108
rect 17960 16065 17969 16099
rect 17969 16065 18003 16099
rect 18003 16065 18012 16099
rect 17960 16056 18012 16065
rect 22100 16056 22152 16108
rect 23664 16056 23716 16108
rect 19340 16031 19392 16040
rect 13360 15852 13412 15904
rect 14924 15895 14976 15904
rect 14924 15861 14933 15895
rect 14933 15861 14967 15895
rect 14967 15861 14976 15895
rect 14924 15852 14976 15861
rect 15108 15895 15160 15904
rect 15108 15861 15117 15895
rect 15117 15861 15151 15895
rect 15151 15861 15160 15895
rect 15108 15852 15160 15861
rect 15568 15852 15620 15904
rect 19340 15997 19349 16031
rect 19349 15997 19383 16031
rect 19383 15997 19392 16031
rect 19340 15988 19392 15997
rect 24492 16056 24544 16108
rect 24676 16056 24728 16108
rect 26148 16124 26200 16176
rect 31024 16167 31076 16176
rect 26240 16099 26292 16108
rect 26240 16065 26249 16099
rect 26249 16065 26283 16099
rect 26283 16065 26292 16099
rect 26240 16056 26292 16065
rect 31024 16133 31033 16167
rect 31033 16133 31067 16167
rect 31067 16133 31076 16167
rect 31024 16124 31076 16133
rect 32312 16124 32364 16176
rect 26700 16056 26752 16108
rect 25596 15988 25648 16040
rect 23756 15920 23808 15972
rect 24768 15920 24820 15972
rect 30748 16056 30800 16108
rect 31116 16099 31168 16108
rect 31116 16065 31125 16099
rect 31125 16065 31159 16099
rect 31159 16065 31168 16099
rect 32956 16124 33008 16176
rect 32588 16099 32640 16108
rect 31116 16056 31168 16065
rect 28816 16031 28868 16040
rect 28816 15997 28825 16031
rect 28825 15997 28859 16031
rect 28859 15997 28868 16031
rect 28816 15988 28868 15997
rect 29000 16031 29052 16040
rect 29000 15997 29009 16031
rect 29009 15997 29043 16031
rect 29043 15997 29052 16031
rect 29000 15988 29052 15997
rect 32588 16065 32597 16099
rect 32597 16065 32631 16099
rect 32631 16065 32640 16099
rect 32588 16056 32640 16065
rect 33692 16056 33744 16108
rect 34704 16056 34756 16108
rect 37280 16099 37332 16108
rect 37280 16065 37289 16099
rect 37289 16065 37323 16099
rect 37323 16065 37332 16099
rect 37280 16056 37332 16065
rect 41420 16201 41429 16235
rect 41429 16201 41463 16235
rect 41463 16201 41472 16235
rect 41420 16192 41472 16201
rect 32680 16031 32732 16040
rect 32680 15997 32689 16031
rect 32689 15997 32723 16031
rect 32723 15997 32732 16031
rect 32680 15988 32732 15997
rect 35348 16031 35400 16040
rect 21824 15852 21876 15904
rect 24584 15852 24636 15904
rect 24860 15852 24912 15904
rect 32588 15920 32640 15972
rect 35348 15997 35357 16031
rect 35357 15997 35391 16031
rect 35391 15997 35400 16031
rect 35348 15988 35400 15997
rect 37464 16031 37516 16040
rect 37464 15997 37473 16031
rect 37473 15997 37507 16031
rect 37507 15997 37516 16031
rect 37464 15988 37516 15997
rect 38936 16031 38988 16040
rect 38936 15997 38945 16031
rect 38945 15997 38979 16031
rect 38979 15997 38988 16031
rect 38936 15988 38988 15997
rect 40960 16056 41012 16108
rect 42340 16056 42392 16108
rect 41880 15988 41932 16040
rect 25596 15895 25648 15904
rect 25596 15861 25605 15895
rect 25605 15861 25639 15895
rect 25639 15861 25648 15895
rect 25596 15852 25648 15861
rect 26148 15852 26200 15904
rect 28908 15895 28960 15904
rect 28908 15861 28917 15895
rect 28917 15861 28951 15895
rect 28951 15861 28960 15895
rect 28908 15852 28960 15861
rect 32036 15852 32088 15904
rect 34612 15852 34664 15904
rect 36084 15852 36136 15904
rect 40316 15852 40368 15904
rect 40500 15852 40552 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 13268 15648 13320 15700
rect 13452 15648 13504 15700
rect 15108 15648 15160 15700
rect 18144 15691 18196 15700
rect 13636 15580 13688 15632
rect 14280 15580 14332 15632
rect 14004 15512 14056 15564
rect 15384 15555 15436 15564
rect 15384 15521 15392 15555
rect 15392 15521 15426 15555
rect 15426 15521 15436 15555
rect 15384 15512 15436 15521
rect 18144 15657 18153 15691
rect 18153 15657 18187 15691
rect 18187 15657 18196 15691
rect 18144 15648 18196 15657
rect 22468 15648 22520 15700
rect 16120 15555 16172 15564
rect 16120 15521 16129 15555
rect 16129 15521 16163 15555
rect 16163 15521 16172 15555
rect 16120 15512 16172 15521
rect 21732 15580 21784 15632
rect 28448 15648 28500 15700
rect 28816 15691 28868 15700
rect 28816 15657 28825 15691
rect 28825 15657 28859 15691
rect 28859 15657 28868 15691
rect 28816 15648 28868 15657
rect 1768 15487 1820 15496
rect 1768 15453 1777 15487
rect 1777 15453 1811 15487
rect 1811 15453 1820 15487
rect 1768 15444 1820 15453
rect 13360 15487 13412 15496
rect 13360 15453 13369 15487
rect 13369 15453 13403 15487
rect 13403 15453 13412 15487
rect 13360 15444 13412 15453
rect 13544 15487 13596 15496
rect 13544 15453 13553 15487
rect 13553 15453 13587 15487
rect 13587 15453 13596 15487
rect 13544 15444 13596 15453
rect 13820 15444 13872 15496
rect 14372 15487 14424 15496
rect 13176 15376 13228 15428
rect 13452 15376 13504 15428
rect 14372 15453 14381 15487
rect 14381 15453 14415 15487
rect 14415 15453 14424 15487
rect 14372 15444 14424 15453
rect 15200 15487 15252 15496
rect 14280 15419 14332 15428
rect 14280 15385 14289 15419
rect 14289 15385 14323 15419
rect 14323 15385 14332 15419
rect 14280 15376 14332 15385
rect 7104 15308 7156 15360
rect 7564 15308 7616 15360
rect 11152 15308 11204 15360
rect 12072 15308 12124 15360
rect 14464 15308 14516 15360
rect 14648 15351 14700 15360
rect 14648 15317 14657 15351
rect 14657 15317 14691 15351
rect 14691 15317 14700 15351
rect 14648 15308 14700 15317
rect 15200 15453 15209 15487
rect 15209 15453 15243 15487
rect 15243 15453 15252 15487
rect 15200 15444 15252 15453
rect 15660 15444 15712 15496
rect 15752 15444 15804 15496
rect 16396 15487 16448 15496
rect 16396 15453 16405 15487
rect 16405 15453 16439 15487
rect 16439 15453 16448 15487
rect 16396 15444 16448 15453
rect 17040 15444 17092 15496
rect 17408 15487 17460 15496
rect 17408 15453 17417 15487
rect 17417 15453 17451 15487
rect 17451 15453 17460 15487
rect 17408 15444 17460 15453
rect 19432 15512 19484 15564
rect 20720 15512 20772 15564
rect 18052 15487 18104 15496
rect 18052 15453 18061 15487
rect 18061 15453 18095 15487
rect 18095 15453 18104 15487
rect 18052 15444 18104 15453
rect 18328 15487 18380 15496
rect 18328 15453 18337 15487
rect 18337 15453 18371 15487
rect 18371 15453 18380 15487
rect 18328 15444 18380 15453
rect 20812 15487 20864 15496
rect 20812 15453 20821 15487
rect 20821 15453 20855 15487
rect 20855 15453 20864 15487
rect 20812 15444 20864 15453
rect 21364 15487 21416 15496
rect 21364 15453 21373 15487
rect 21373 15453 21407 15487
rect 21407 15453 21416 15487
rect 21364 15444 21416 15453
rect 21824 15487 21876 15496
rect 21824 15453 21833 15487
rect 21833 15453 21867 15487
rect 21867 15453 21876 15487
rect 21824 15444 21876 15453
rect 24860 15512 24912 15564
rect 24768 15444 24820 15496
rect 26700 15444 26752 15496
rect 27712 15487 27764 15496
rect 27712 15453 27746 15487
rect 27746 15453 27764 15487
rect 32588 15648 32640 15700
rect 33692 15691 33744 15700
rect 33692 15657 33701 15691
rect 33701 15657 33735 15691
rect 33735 15657 33744 15691
rect 33692 15648 33744 15657
rect 37464 15648 37516 15700
rect 34796 15580 34848 15632
rect 35532 15580 35584 15632
rect 29368 15512 29420 15564
rect 32956 15512 33008 15564
rect 34704 15555 34756 15564
rect 27712 15444 27764 15453
rect 29644 15444 29696 15496
rect 32864 15444 32916 15496
rect 33324 15487 33376 15496
rect 33324 15453 33333 15487
rect 33333 15453 33367 15487
rect 33367 15453 33376 15487
rect 34704 15521 34713 15555
rect 34713 15521 34747 15555
rect 34747 15521 34756 15555
rect 34704 15512 34756 15521
rect 33324 15444 33376 15453
rect 35900 15487 35952 15496
rect 35900 15453 35909 15487
rect 35909 15453 35943 15487
rect 35943 15453 35952 15487
rect 35900 15444 35952 15453
rect 36544 15444 36596 15496
rect 41512 15580 41564 15632
rect 40316 15555 40368 15564
rect 40316 15521 40325 15555
rect 40325 15521 40359 15555
rect 40359 15521 40368 15555
rect 40316 15512 40368 15521
rect 40500 15555 40552 15564
rect 40500 15521 40509 15555
rect 40509 15521 40543 15555
rect 40543 15521 40552 15555
rect 40500 15512 40552 15521
rect 42156 15555 42208 15564
rect 42156 15521 42165 15555
rect 42165 15521 42199 15555
rect 42199 15521 42208 15555
rect 42156 15512 42208 15521
rect 19340 15376 19392 15428
rect 20720 15376 20772 15428
rect 22652 15376 22704 15428
rect 15476 15308 15528 15360
rect 18420 15308 18472 15360
rect 20536 15308 20588 15360
rect 26884 15308 26936 15360
rect 30932 15351 30984 15360
rect 30932 15317 30941 15351
rect 30941 15317 30975 15351
rect 30975 15317 30984 15351
rect 30932 15308 30984 15317
rect 35348 15308 35400 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 13176 15147 13228 15156
rect 13176 15113 13185 15147
rect 13185 15113 13219 15147
rect 13219 15113 13228 15147
rect 13176 15104 13228 15113
rect 13544 15104 13596 15156
rect 15016 15104 15068 15156
rect 1768 15011 1820 15020
rect 1768 14977 1777 15011
rect 1777 14977 1811 15011
rect 1811 14977 1820 15011
rect 1768 14968 1820 14977
rect 13452 15011 13504 15020
rect 13452 14977 13461 15011
rect 13461 14977 13495 15011
rect 13495 14977 13504 15011
rect 13452 14968 13504 14977
rect 14648 15036 14700 15088
rect 15200 15036 15252 15088
rect 14188 14968 14240 15020
rect 14280 14968 14332 15020
rect 15108 14968 15160 15020
rect 17408 15104 17460 15156
rect 25596 15104 25648 15156
rect 19064 15036 19116 15088
rect 20444 15036 20496 15088
rect 22744 15079 22796 15088
rect 15476 15011 15528 15020
rect 15476 14977 15485 15011
rect 15485 14977 15519 15011
rect 15519 14977 15528 15011
rect 15476 14968 15528 14977
rect 2228 14900 2280 14952
rect 2780 14943 2832 14952
rect 2780 14909 2789 14943
rect 2789 14909 2823 14943
rect 2823 14909 2832 14943
rect 2780 14900 2832 14909
rect 16396 14968 16448 15020
rect 15936 14900 15988 14952
rect 18328 14968 18380 15020
rect 20076 14968 20128 15020
rect 20536 14968 20588 15020
rect 22744 15045 22753 15079
rect 22753 15045 22787 15079
rect 22787 15045 22796 15079
rect 22744 15036 22796 15045
rect 24400 15036 24452 15088
rect 24768 15079 24820 15088
rect 24768 15045 24777 15079
rect 24777 15045 24811 15079
rect 24811 15045 24820 15079
rect 24768 15036 24820 15045
rect 30932 15079 30984 15088
rect 26884 14968 26936 15020
rect 30932 15045 30941 15079
rect 30941 15045 30975 15079
rect 30975 15045 30984 15079
rect 30932 15036 30984 15045
rect 14096 14832 14148 14884
rect 18420 14832 18472 14884
rect 34704 14968 34756 15020
rect 35532 15011 35584 15020
rect 35532 14977 35541 15011
rect 35541 14977 35575 15011
rect 35575 14977 35584 15011
rect 35532 14968 35584 14977
rect 41328 14943 41380 14952
rect 41328 14909 41337 14943
rect 41337 14909 41371 14943
rect 41371 14909 41380 14943
rect 41328 14900 41380 14909
rect 41420 14900 41472 14952
rect 41972 14900 42024 14952
rect 22284 14832 22336 14884
rect 38476 14832 38528 14884
rect 17960 14764 18012 14816
rect 19616 14764 19668 14816
rect 22376 14764 22428 14816
rect 22652 14764 22704 14816
rect 23480 14764 23532 14816
rect 24676 14764 24728 14816
rect 25228 14764 25280 14816
rect 30196 14807 30248 14816
rect 30196 14773 30205 14807
rect 30205 14773 30239 14807
rect 30239 14773 30248 14807
rect 30196 14764 30248 14773
rect 31668 14764 31720 14816
rect 35808 14764 35860 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 2228 14603 2280 14612
rect 2228 14569 2237 14603
rect 2237 14569 2271 14603
rect 2271 14569 2280 14603
rect 2228 14560 2280 14569
rect 13820 14560 13872 14612
rect 15200 14560 15252 14612
rect 19616 14603 19668 14612
rect 2964 14356 3016 14408
rect 11612 14356 11664 14408
rect 13544 14424 13596 14476
rect 13452 14399 13504 14408
rect 13452 14365 13461 14399
rect 13461 14365 13495 14399
rect 13495 14365 13504 14399
rect 13452 14356 13504 14365
rect 11796 14220 11848 14272
rect 14372 14263 14424 14272
rect 14372 14229 14381 14263
rect 14381 14229 14415 14263
rect 14415 14229 14424 14263
rect 14372 14220 14424 14229
rect 15568 14492 15620 14544
rect 15660 14492 15712 14544
rect 19616 14569 19625 14603
rect 19625 14569 19659 14603
rect 19659 14569 19668 14603
rect 19616 14560 19668 14569
rect 20996 14560 21048 14612
rect 22192 14560 22244 14612
rect 22744 14560 22796 14612
rect 34520 14560 34572 14612
rect 35532 14603 35584 14612
rect 35532 14569 35541 14603
rect 35541 14569 35575 14603
rect 35575 14569 35584 14603
rect 35532 14560 35584 14569
rect 35900 14560 35952 14612
rect 36268 14560 36320 14612
rect 41420 14603 41472 14612
rect 41420 14569 41429 14603
rect 41429 14569 41463 14603
rect 41463 14569 41472 14603
rect 41420 14560 41472 14569
rect 41972 14603 42024 14612
rect 41972 14569 41981 14603
rect 41981 14569 42015 14603
rect 42015 14569 42024 14603
rect 41972 14560 42024 14569
rect 23572 14535 23624 14544
rect 17408 14424 17460 14476
rect 23572 14501 23581 14535
rect 23581 14501 23615 14535
rect 23615 14501 23624 14535
rect 23572 14492 23624 14501
rect 31852 14492 31904 14544
rect 18052 14424 18104 14476
rect 20168 14424 20220 14476
rect 15016 14399 15068 14408
rect 15016 14365 15025 14399
rect 15025 14365 15059 14399
rect 15059 14365 15068 14399
rect 15016 14356 15068 14365
rect 15108 14356 15160 14408
rect 15936 14399 15988 14408
rect 15936 14365 15945 14399
rect 15945 14365 15979 14399
rect 15979 14365 15988 14399
rect 15936 14356 15988 14365
rect 19432 14399 19484 14408
rect 19432 14365 19441 14399
rect 19441 14365 19475 14399
rect 19475 14365 19484 14399
rect 19432 14356 19484 14365
rect 20260 14399 20312 14408
rect 20260 14365 20269 14399
rect 20269 14365 20303 14399
rect 20303 14365 20312 14399
rect 20260 14356 20312 14365
rect 20444 14356 20496 14408
rect 16396 14288 16448 14340
rect 21732 14331 21784 14340
rect 21732 14297 21741 14331
rect 21741 14297 21775 14331
rect 21775 14297 21784 14331
rect 21732 14288 21784 14297
rect 16672 14220 16724 14272
rect 20444 14220 20496 14272
rect 26240 14399 26292 14408
rect 26240 14365 26249 14399
rect 26249 14365 26283 14399
rect 26283 14365 26292 14399
rect 26700 14399 26752 14408
rect 26240 14356 26292 14365
rect 26700 14365 26709 14399
rect 26709 14365 26743 14399
rect 26743 14365 26752 14399
rect 26700 14356 26752 14365
rect 26148 14288 26200 14340
rect 26884 14288 26936 14340
rect 29000 14220 29052 14272
rect 29736 14288 29788 14340
rect 31760 14356 31812 14408
rect 32036 14399 32088 14408
rect 32036 14365 32045 14399
rect 32045 14365 32079 14399
rect 32079 14365 32088 14399
rect 32036 14356 32088 14365
rect 32220 14356 32272 14408
rect 33600 14399 33652 14408
rect 33600 14365 33609 14399
rect 33609 14365 33643 14399
rect 33643 14365 33652 14399
rect 33600 14356 33652 14365
rect 33784 14399 33836 14408
rect 33784 14365 33793 14399
rect 33793 14365 33827 14399
rect 33827 14365 33836 14399
rect 33784 14356 33836 14365
rect 34612 14356 34664 14408
rect 35716 14399 35768 14408
rect 35716 14365 35725 14399
rect 35725 14365 35759 14399
rect 35759 14365 35768 14399
rect 35716 14356 35768 14365
rect 36084 14399 36136 14408
rect 36084 14365 36093 14399
rect 36093 14365 36127 14399
rect 36127 14365 36136 14399
rect 36084 14356 36136 14365
rect 30380 14288 30432 14340
rect 34520 14288 34572 14340
rect 35348 14288 35400 14340
rect 35532 14288 35584 14340
rect 37188 14356 37240 14408
rect 41236 14356 41288 14408
rect 30288 14220 30340 14272
rect 33416 14220 33468 14272
rect 34704 14263 34756 14272
rect 34704 14229 34713 14263
rect 34713 14229 34747 14263
rect 34747 14229 34756 14263
rect 34704 14220 34756 14229
rect 34980 14220 35032 14272
rect 36636 14263 36688 14272
rect 36636 14229 36645 14263
rect 36645 14229 36679 14263
rect 36679 14229 36688 14263
rect 36636 14220 36688 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 15936 14016 15988 14068
rect 14372 13991 14424 14000
rect 14372 13957 14406 13991
rect 14406 13957 14424 13991
rect 14372 13948 14424 13957
rect 15660 13948 15712 14000
rect 20260 14016 20312 14068
rect 24400 14016 24452 14068
rect 26148 14059 26200 14068
rect 26148 14025 26157 14059
rect 26157 14025 26191 14059
rect 26191 14025 26200 14059
rect 26148 14016 26200 14025
rect 16580 13948 16632 14000
rect 11796 13923 11848 13932
rect 11796 13889 11805 13923
rect 11805 13889 11839 13923
rect 11839 13889 11848 13923
rect 11796 13880 11848 13889
rect 14096 13923 14148 13932
rect 14096 13889 14105 13923
rect 14105 13889 14139 13923
rect 14139 13889 14148 13923
rect 14096 13880 14148 13889
rect 1952 13855 2004 13864
rect 1952 13821 1961 13855
rect 1961 13821 1995 13855
rect 1995 13821 2004 13855
rect 1952 13812 2004 13821
rect 2780 13812 2832 13864
rect 2872 13855 2924 13864
rect 2872 13821 2881 13855
rect 2881 13821 2915 13855
rect 2915 13821 2924 13855
rect 11980 13855 12032 13864
rect 2872 13812 2924 13821
rect 11980 13821 11989 13855
rect 11989 13821 12023 13855
rect 12023 13821 12032 13855
rect 11980 13812 12032 13821
rect 13636 13855 13688 13864
rect 13636 13821 13645 13855
rect 13645 13821 13679 13855
rect 13679 13821 13688 13855
rect 13636 13812 13688 13821
rect 16948 13812 17000 13864
rect 20168 13948 20220 14000
rect 20720 13948 20772 14000
rect 22100 13991 22152 14000
rect 22100 13957 22109 13991
rect 22109 13957 22143 13991
rect 22143 13957 22152 13991
rect 22100 13948 22152 13957
rect 22284 13948 22336 14000
rect 23112 13948 23164 14000
rect 31852 14016 31904 14068
rect 32220 14059 32272 14068
rect 32220 14025 32229 14059
rect 32229 14025 32263 14059
rect 32263 14025 32272 14059
rect 32220 14016 32272 14025
rect 35992 14016 36044 14068
rect 30012 13948 30064 14000
rect 18328 13812 18380 13864
rect 19984 13923 20036 13932
rect 19984 13889 19993 13923
rect 19993 13889 20027 13923
rect 20027 13889 20036 13923
rect 19984 13880 20036 13889
rect 20352 13880 20404 13932
rect 20352 13744 20404 13796
rect 21364 13880 21416 13932
rect 33600 13948 33652 14000
rect 22468 13880 22520 13932
rect 24584 13880 24636 13932
rect 25228 13923 25280 13932
rect 25228 13889 25237 13923
rect 25237 13889 25271 13923
rect 25271 13889 25280 13923
rect 25228 13880 25280 13889
rect 20720 13855 20772 13864
rect 20720 13821 20729 13855
rect 20729 13821 20763 13855
rect 20763 13821 20772 13855
rect 20720 13812 20772 13821
rect 24676 13812 24728 13864
rect 28172 13880 28224 13932
rect 30104 13923 30156 13932
rect 30104 13889 30113 13923
rect 30113 13889 30147 13923
rect 30147 13889 30156 13923
rect 30104 13880 30156 13889
rect 30288 13923 30340 13932
rect 30288 13889 30297 13923
rect 30297 13889 30331 13923
rect 30331 13889 30340 13923
rect 30288 13880 30340 13889
rect 30196 13812 30248 13864
rect 31668 13880 31720 13932
rect 33232 13923 33284 13932
rect 27528 13787 27580 13796
rect 27528 13753 27537 13787
rect 27537 13753 27571 13787
rect 27571 13753 27580 13787
rect 27528 13744 27580 13753
rect 31760 13812 31812 13864
rect 33232 13889 33241 13923
rect 33241 13889 33275 13923
rect 33275 13889 33284 13923
rect 33232 13880 33284 13889
rect 34428 13880 34480 13932
rect 33048 13744 33100 13796
rect 34796 13923 34848 13932
rect 34796 13889 34831 13923
rect 34831 13889 34848 13923
rect 34796 13880 34848 13889
rect 35716 13880 35768 13932
rect 35808 13880 35860 13932
rect 37372 13880 37424 13932
rect 34980 13855 35032 13864
rect 34980 13821 34989 13855
rect 34989 13821 35023 13855
rect 35023 13821 35032 13855
rect 34980 13812 35032 13821
rect 36176 13812 36228 13864
rect 34612 13744 34664 13796
rect 36820 13744 36872 13796
rect 16856 13719 16908 13728
rect 16856 13685 16865 13719
rect 16865 13685 16899 13719
rect 16899 13685 16908 13719
rect 16856 13676 16908 13685
rect 17868 13719 17920 13728
rect 17868 13685 17877 13719
rect 17877 13685 17911 13719
rect 17911 13685 17920 13719
rect 17868 13676 17920 13685
rect 19984 13676 20036 13728
rect 20444 13676 20496 13728
rect 25320 13719 25372 13728
rect 25320 13685 25329 13719
rect 25329 13685 25363 13719
rect 25363 13685 25372 13719
rect 25320 13676 25372 13685
rect 30748 13676 30800 13728
rect 31024 13676 31076 13728
rect 32864 13719 32916 13728
rect 32864 13685 32873 13719
rect 32873 13685 32907 13719
rect 32907 13685 32916 13719
rect 32864 13676 32916 13685
rect 34336 13719 34388 13728
rect 34336 13685 34345 13719
rect 34345 13685 34379 13719
rect 34379 13685 34388 13719
rect 34336 13676 34388 13685
rect 41788 13719 41840 13728
rect 41788 13685 41797 13719
rect 41797 13685 41831 13719
rect 41831 13685 41840 13719
rect 41788 13676 41840 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 1952 13472 2004 13524
rect 2780 13515 2832 13524
rect 2780 13481 2789 13515
rect 2789 13481 2823 13515
rect 2823 13481 2832 13515
rect 2780 13472 2832 13481
rect 11980 13472 12032 13524
rect 15200 13404 15252 13456
rect 16304 13404 16356 13456
rect 9404 13268 9456 13320
rect 10692 13268 10744 13320
rect 12808 13311 12860 13320
rect 12808 13277 12817 13311
rect 12817 13277 12851 13311
rect 12851 13277 12860 13311
rect 12808 13268 12860 13277
rect 16120 13311 16172 13320
rect 16120 13277 16129 13311
rect 16129 13277 16163 13311
rect 16163 13277 16172 13311
rect 16672 13336 16724 13388
rect 16120 13268 16172 13277
rect 16580 13311 16632 13320
rect 16580 13277 16589 13311
rect 16589 13277 16623 13311
rect 16623 13277 16632 13311
rect 16580 13268 16632 13277
rect 17868 13404 17920 13456
rect 16856 13336 16908 13388
rect 20260 13379 20312 13388
rect 20260 13345 20269 13379
rect 20269 13345 20303 13379
rect 20303 13345 20312 13379
rect 22652 13472 22704 13524
rect 25136 13472 25188 13524
rect 28172 13515 28224 13524
rect 28172 13481 28181 13515
rect 28181 13481 28215 13515
rect 28215 13481 28224 13515
rect 28172 13472 28224 13481
rect 28908 13472 28960 13524
rect 34796 13472 34848 13524
rect 22468 13379 22520 13388
rect 20260 13336 20312 13345
rect 22468 13345 22477 13379
rect 22477 13345 22511 13379
rect 22511 13345 22520 13379
rect 22468 13336 22520 13345
rect 20720 13268 20772 13320
rect 21548 13311 21600 13320
rect 21548 13277 21557 13311
rect 21557 13277 21591 13311
rect 21591 13277 21600 13311
rect 21548 13268 21600 13277
rect 12348 13132 12400 13184
rect 16488 13200 16540 13252
rect 16396 13132 16448 13184
rect 18052 13175 18104 13184
rect 18052 13141 18061 13175
rect 18061 13141 18095 13175
rect 18095 13141 18104 13175
rect 18052 13132 18104 13141
rect 20536 13132 20588 13184
rect 22376 13268 22428 13320
rect 24676 13311 24728 13320
rect 24676 13277 24685 13311
rect 24685 13277 24719 13311
rect 24719 13277 24728 13311
rect 24676 13268 24728 13277
rect 25228 13336 25280 13388
rect 25320 13311 25372 13320
rect 25320 13277 25329 13311
rect 25329 13277 25363 13311
rect 25363 13277 25372 13311
rect 25320 13268 25372 13277
rect 30288 13336 30340 13388
rect 33048 13404 33100 13456
rect 33416 13379 33468 13388
rect 33416 13345 33425 13379
rect 33425 13345 33459 13379
rect 33459 13345 33468 13379
rect 33416 13336 33468 13345
rect 29276 13268 29328 13320
rect 30104 13311 30156 13320
rect 30104 13277 30113 13311
rect 30113 13277 30147 13311
rect 30147 13277 30156 13311
rect 30104 13268 30156 13277
rect 31024 13311 31076 13320
rect 31024 13277 31033 13311
rect 31033 13277 31067 13311
rect 31067 13277 31076 13311
rect 31024 13268 31076 13277
rect 32220 13268 32272 13320
rect 34336 13268 34388 13320
rect 34520 13268 34572 13320
rect 24216 13132 24268 13184
rect 27252 13200 27304 13252
rect 30288 13243 30340 13252
rect 30288 13209 30297 13243
rect 30297 13209 30331 13243
rect 30331 13209 30340 13243
rect 30288 13200 30340 13209
rect 36544 13472 36596 13524
rect 36820 13515 36872 13524
rect 36820 13481 36829 13515
rect 36829 13481 36863 13515
rect 36863 13481 36872 13515
rect 36820 13472 36872 13481
rect 35716 13404 35768 13456
rect 41328 13379 41380 13388
rect 41328 13345 41337 13379
rect 41337 13345 41371 13379
rect 41371 13345 41380 13379
rect 41328 13336 41380 13345
rect 41788 13336 41840 13388
rect 35716 13311 35768 13320
rect 35716 13277 35725 13311
rect 35725 13277 35759 13311
rect 35759 13277 35768 13311
rect 35716 13268 35768 13277
rect 36176 13268 36228 13320
rect 37372 13311 37424 13320
rect 28356 13175 28408 13184
rect 28356 13141 28365 13175
rect 28365 13141 28399 13175
rect 28399 13141 28408 13175
rect 28356 13132 28408 13141
rect 28448 13132 28500 13184
rect 35348 13200 35400 13252
rect 35532 13200 35584 13252
rect 36268 13200 36320 13252
rect 37372 13277 37381 13311
rect 37381 13277 37415 13311
rect 37415 13277 37424 13311
rect 37372 13268 37424 13277
rect 41512 13200 41564 13252
rect 32312 13132 32364 13184
rect 35256 13132 35308 13184
rect 36176 13132 36228 13184
rect 37464 13175 37516 13184
rect 37464 13141 37473 13175
rect 37473 13141 37507 13175
rect 37507 13141 37516 13175
rect 37464 13132 37516 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 12808 12928 12860 12980
rect 12348 12903 12400 12912
rect 12348 12869 12357 12903
rect 12357 12869 12391 12903
rect 12391 12869 12400 12903
rect 12348 12860 12400 12869
rect 17224 12860 17276 12912
rect 18052 12860 18104 12912
rect 15200 12835 15252 12844
rect 15200 12801 15209 12835
rect 15209 12801 15243 12835
rect 15243 12801 15252 12835
rect 15200 12792 15252 12801
rect 12716 12724 12768 12776
rect 13728 12767 13780 12776
rect 13728 12733 13737 12767
rect 13737 12733 13771 12767
rect 13771 12733 13780 12767
rect 13728 12724 13780 12733
rect 15936 12767 15988 12776
rect 15936 12733 15945 12767
rect 15945 12733 15979 12767
rect 15979 12733 15988 12767
rect 15936 12724 15988 12733
rect 16304 12792 16356 12844
rect 16488 12792 16540 12844
rect 16948 12767 17000 12776
rect 16948 12733 16957 12767
rect 16957 12733 16991 12767
rect 16991 12733 17000 12767
rect 16948 12724 17000 12733
rect 17960 12792 18012 12844
rect 13820 12656 13872 12708
rect 16304 12656 16356 12708
rect 20260 12928 20312 12980
rect 21180 12971 21232 12980
rect 21180 12937 21189 12971
rect 21189 12937 21223 12971
rect 21223 12937 21232 12971
rect 21180 12928 21232 12937
rect 21548 12928 21600 12980
rect 20352 12792 20404 12844
rect 21088 12792 21140 12844
rect 28448 12928 28500 12980
rect 29276 12971 29328 12980
rect 29276 12937 29285 12971
rect 29285 12937 29319 12971
rect 29319 12937 29328 12971
rect 29276 12928 29328 12937
rect 30288 12928 30340 12980
rect 32220 12971 32272 12980
rect 27528 12860 27580 12912
rect 23940 12835 23992 12844
rect 23940 12801 23949 12835
rect 23949 12801 23983 12835
rect 23983 12801 23992 12835
rect 23940 12792 23992 12801
rect 24216 12835 24268 12844
rect 24216 12801 24225 12835
rect 24225 12801 24259 12835
rect 24259 12801 24268 12835
rect 24216 12792 24268 12801
rect 27252 12835 27304 12844
rect 27252 12801 27286 12835
rect 27286 12801 27304 12835
rect 27252 12792 27304 12801
rect 28816 12835 28868 12844
rect 28816 12801 28825 12835
rect 28825 12801 28859 12835
rect 28859 12801 28868 12835
rect 28816 12792 28868 12801
rect 29092 12835 29144 12844
rect 29092 12801 29101 12835
rect 29101 12801 29135 12835
rect 29135 12801 29144 12835
rect 29092 12792 29144 12801
rect 24124 12767 24176 12776
rect 24124 12733 24133 12767
rect 24133 12733 24167 12767
rect 24167 12733 24176 12767
rect 24124 12724 24176 12733
rect 25136 12767 25188 12776
rect 25136 12733 25145 12767
rect 25145 12733 25179 12767
rect 25179 12733 25188 12767
rect 25136 12724 25188 12733
rect 26976 12767 27028 12776
rect 26976 12733 26985 12767
rect 26985 12733 27019 12767
rect 27019 12733 27028 12767
rect 26976 12724 27028 12733
rect 29000 12767 29052 12776
rect 29000 12733 29009 12767
rect 29009 12733 29043 12767
rect 29043 12733 29052 12767
rect 29000 12724 29052 12733
rect 32220 12937 32229 12971
rect 32229 12937 32263 12971
rect 32263 12937 32272 12971
rect 32220 12928 32272 12937
rect 33232 12928 33284 12980
rect 33784 12928 33836 12980
rect 34704 12928 34756 12980
rect 35992 12971 36044 12980
rect 35992 12937 36001 12971
rect 36001 12937 36035 12971
rect 36035 12937 36044 12971
rect 35992 12928 36044 12937
rect 41512 12971 41564 12980
rect 41512 12937 41521 12971
rect 41521 12937 41555 12971
rect 41555 12937 41564 12971
rect 41512 12928 41564 12937
rect 30748 12835 30800 12844
rect 30748 12801 30757 12835
rect 30757 12801 30791 12835
rect 30791 12801 30800 12835
rect 30748 12792 30800 12801
rect 31208 12792 31260 12844
rect 31484 12792 31536 12844
rect 34796 12792 34848 12844
rect 37464 12860 37516 12912
rect 35716 12792 35768 12844
rect 36268 12835 36320 12844
rect 36268 12801 36277 12835
rect 36277 12801 36311 12835
rect 36311 12801 36320 12835
rect 36268 12792 36320 12801
rect 31024 12724 31076 12776
rect 35256 12767 35308 12776
rect 1676 12631 1728 12640
rect 1676 12597 1685 12631
rect 1685 12597 1719 12631
rect 1719 12597 1728 12631
rect 1676 12588 1728 12597
rect 16672 12588 16724 12640
rect 20536 12656 20588 12708
rect 22192 12631 22244 12640
rect 22192 12597 22201 12631
rect 22201 12597 22235 12631
rect 22235 12597 22244 12631
rect 22192 12588 22244 12597
rect 24676 12656 24728 12708
rect 26056 12656 26108 12708
rect 26240 12656 26292 12708
rect 24400 12631 24452 12640
rect 24400 12597 24409 12631
rect 24409 12597 24443 12631
rect 24443 12597 24452 12631
rect 24400 12588 24452 12597
rect 26332 12588 26384 12640
rect 26976 12588 27028 12640
rect 30380 12656 30432 12708
rect 30840 12656 30892 12708
rect 30472 12588 30524 12640
rect 35256 12733 35265 12767
rect 35265 12733 35299 12767
rect 35299 12733 35308 12767
rect 35256 12724 35308 12733
rect 35532 12724 35584 12776
rect 36360 12656 36412 12708
rect 36636 12835 36688 12844
rect 36636 12801 36645 12835
rect 36645 12801 36679 12835
rect 36679 12801 36688 12835
rect 36636 12792 36688 12801
rect 37188 12792 37240 12844
rect 41420 12835 41472 12844
rect 41420 12801 41429 12835
rect 41429 12801 41463 12835
rect 41463 12801 41472 12835
rect 41420 12792 41472 12801
rect 41696 12792 41748 12844
rect 40776 12631 40828 12640
rect 40776 12597 40785 12631
rect 40785 12597 40819 12631
rect 40819 12597 40828 12631
rect 40776 12588 40828 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 9404 12384 9456 12436
rect 11704 12384 11756 12436
rect 12716 12427 12768 12436
rect 12716 12393 12725 12427
rect 12725 12393 12759 12427
rect 12759 12393 12768 12427
rect 12716 12384 12768 12393
rect 16120 12384 16172 12436
rect 16580 12384 16632 12436
rect 17224 12427 17276 12436
rect 17224 12393 17233 12427
rect 17233 12393 17267 12427
rect 17267 12393 17276 12427
rect 17224 12384 17276 12393
rect 20168 12427 20220 12436
rect 20168 12393 20177 12427
rect 20177 12393 20211 12427
rect 20211 12393 20220 12427
rect 20168 12384 20220 12393
rect 20352 12427 20404 12436
rect 20352 12393 20361 12427
rect 20361 12393 20395 12427
rect 20395 12393 20404 12427
rect 20352 12384 20404 12393
rect 24400 12427 24452 12436
rect 24400 12393 24409 12427
rect 24409 12393 24443 12427
rect 24443 12393 24452 12427
rect 24400 12384 24452 12393
rect 24768 12427 24820 12436
rect 24768 12393 24777 12427
rect 24777 12393 24811 12427
rect 24811 12393 24820 12427
rect 24768 12384 24820 12393
rect 28816 12384 28868 12436
rect 34704 12384 34756 12436
rect 17868 12316 17920 12368
rect 19340 12359 19392 12368
rect 19340 12325 19349 12359
rect 19349 12325 19383 12359
rect 19383 12325 19392 12359
rect 19340 12316 19392 12325
rect 1676 12248 1728 12300
rect 2780 12291 2832 12300
rect 2780 12257 2789 12291
rect 2789 12257 2823 12291
rect 2823 12257 2832 12291
rect 2780 12248 2832 12257
rect 14096 12248 14148 12300
rect 13820 12180 13872 12232
rect 16304 12180 16356 12232
rect 16948 12180 17000 12232
rect 18328 12180 18380 12232
rect 20444 12248 20496 12300
rect 2136 12112 2188 12164
rect 14740 12112 14792 12164
rect 17500 12112 17552 12164
rect 16304 12044 16356 12096
rect 19156 12044 19208 12096
rect 21180 12223 21232 12232
rect 21180 12189 21189 12223
rect 21189 12189 21223 12223
rect 21223 12189 21232 12223
rect 21180 12180 21232 12189
rect 21272 12180 21324 12232
rect 25136 12180 25188 12232
rect 26056 12223 26108 12232
rect 26056 12189 26065 12223
rect 26065 12189 26099 12223
rect 26099 12189 26108 12223
rect 26056 12180 26108 12189
rect 26332 12223 26384 12232
rect 26332 12189 26366 12223
rect 26366 12189 26384 12223
rect 33416 12248 33468 12300
rect 33600 12248 33652 12300
rect 28632 12223 28684 12232
rect 26332 12180 26384 12189
rect 28632 12189 28641 12223
rect 28641 12189 28675 12223
rect 28675 12189 28684 12223
rect 28632 12180 28684 12189
rect 30472 12223 30524 12232
rect 30472 12189 30481 12223
rect 30481 12189 30515 12223
rect 30515 12189 30524 12223
rect 30472 12180 30524 12189
rect 32312 12223 32364 12232
rect 32312 12189 32321 12223
rect 32321 12189 32355 12223
rect 32355 12189 32364 12223
rect 32312 12180 32364 12189
rect 32864 12180 32916 12232
rect 34520 12248 34572 12300
rect 34796 12248 34848 12300
rect 20536 12155 20588 12164
rect 20536 12121 20545 12155
rect 20545 12121 20579 12155
rect 20579 12121 20588 12155
rect 20536 12112 20588 12121
rect 20996 12044 21048 12096
rect 21640 12044 21692 12096
rect 31944 12087 31996 12096
rect 31944 12053 31953 12087
rect 31953 12053 31987 12087
rect 31987 12053 31996 12087
rect 31944 12044 31996 12053
rect 33508 12044 33560 12096
rect 40776 12248 40828 12300
rect 42156 12291 42208 12300
rect 42156 12257 42165 12291
rect 42165 12257 42199 12291
rect 42199 12257 42208 12291
rect 42156 12248 42208 12257
rect 36084 12180 36136 12232
rect 35624 12112 35676 12164
rect 35808 12112 35860 12164
rect 36268 12112 36320 12164
rect 37004 12223 37056 12232
rect 37004 12189 37013 12223
rect 37013 12189 37047 12223
rect 37047 12189 37056 12223
rect 37004 12180 37056 12189
rect 41512 12112 41564 12164
rect 35164 12044 35216 12096
rect 35992 12044 36044 12096
rect 36360 12087 36412 12096
rect 36360 12053 36369 12087
rect 36369 12053 36403 12087
rect 36403 12053 36412 12087
rect 36360 12044 36412 12053
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 2136 11883 2188 11892
rect 2136 11849 2145 11883
rect 2145 11849 2179 11883
rect 2179 11849 2188 11883
rect 2136 11840 2188 11849
rect 14740 11883 14792 11892
rect 14740 11849 14749 11883
rect 14749 11849 14783 11883
rect 14783 11849 14792 11883
rect 14740 11840 14792 11849
rect 17224 11840 17276 11892
rect 2320 11704 2372 11756
rect 9404 11747 9456 11756
rect 9404 11713 9413 11747
rect 9413 11713 9447 11747
rect 9447 11713 9456 11747
rect 9404 11704 9456 11713
rect 16304 11704 16356 11756
rect 16488 11704 16540 11756
rect 18236 11636 18288 11688
rect 19524 11772 19576 11824
rect 19708 11772 19760 11824
rect 20352 11840 20404 11892
rect 23940 11840 23992 11892
rect 24124 11840 24176 11892
rect 29092 11840 29144 11892
rect 27160 11772 27212 11824
rect 33600 11772 33652 11824
rect 34428 11815 34480 11824
rect 34428 11781 34437 11815
rect 34437 11781 34471 11815
rect 34471 11781 34480 11815
rect 34428 11772 34480 11781
rect 21180 11704 21232 11756
rect 22468 11747 22520 11756
rect 22468 11713 22477 11747
rect 22477 11713 22511 11747
rect 22511 11713 22520 11747
rect 22468 11704 22520 11713
rect 22560 11704 22612 11756
rect 23480 11704 23532 11756
rect 26976 11747 27028 11756
rect 26976 11713 26985 11747
rect 26985 11713 27019 11747
rect 27019 11713 27028 11747
rect 26976 11704 27028 11713
rect 31944 11704 31996 11756
rect 33048 11704 33100 11756
rect 33692 11747 33744 11756
rect 33692 11713 33701 11747
rect 33701 11713 33735 11747
rect 33735 11713 33744 11747
rect 33692 11704 33744 11713
rect 34980 11772 35032 11824
rect 36176 11840 36228 11892
rect 37004 11840 37056 11892
rect 41512 11883 41564 11892
rect 41512 11849 41521 11883
rect 41521 11849 41555 11883
rect 41555 11849 41564 11883
rect 41512 11840 41564 11849
rect 34612 11747 34664 11756
rect 34612 11713 34621 11747
rect 34621 11713 34655 11747
rect 34655 11713 34664 11747
rect 36084 11772 36136 11824
rect 34612 11704 34664 11713
rect 36268 11704 36320 11756
rect 37004 11704 37056 11756
rect 41420 11704 41472 11756
rect 9220 11500 9272 11552
rect 19340 11500 19392 11552
rect 19432 11543 19484 11552
rect 19432 11509 19441 11543
rect 19441 11509 19475 11543
rect 19475 11509 19484 11543
rect 19432 11500 19484 11509
rect 24584 11500 24636 11552
rect 25320 11500 25372 11552
rect 26056 11636 26108 11688
rect 35992 11636 36044 11688
rect 36820 11636 36872 11688
rect 35624 11568 35676 11620
rect 36268 11568 36320 11620
rect 30472 11543 30524 11552
rect 30472 11509 30481 11543
rect 30481 11509 30515 11543
rect 30515 11509 30524 11543
rect 30472 11500 30524 11509
rect 33232 11543 33284 11552
rect 33232 11509 33241 11543
rect 33241 11509 33275 11543
rect 33275 11509 33284 11543
rect 33232 11500 33284 11509
rect 34336 11543 34388 11552
rect 34336 11509 34345 11543
rect 34345 11509 34379 11543
rect 34379 11509 34388 11543
rect 34336 11500 34388 11509
rect 35992 11500 36044 11552
rect 40316 11500 40368 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 19524 11339 19576 11348
rect 19524 11305 19533 11339
rect 19533 11305 19567 11339
rect 19567 11305 19576 11339
rect 19524 11296 19576 11305
rect 20996 11339 21048 11348
rect 20996 11305 21005 11339
rect 21005 11305 21039 11339
rect 21039 11305 21048 11339
rect 20996 11296 21048 11305
rect 21180 11296 21232 11348
rect 22836 11339 22888 11348
rect 22836 11305 22845 11339
rect 22845 11305 22879 11339
rect 22879 11305 22888 11339
rect 22836 11296 22888 11305
rect 24032 11296 24084 11348
rect 35900 11228 35952 11280
rect 19432 11160 19484 11212
rect 1676 11135 1728 11144
rect 1676 11101 1685 11135
rect 1685 11101 1719 11135
rect 1719 11101 1728 11135
rect 1676 11092 1728 11101
rect 17224 11135 17276 11144
rect 17224 11101 17233 11135
rect 17233 11101 17267 11135
rect 17267 11101 17276 11135
rect 17224 11092 17276 11101
rect 17500 11092 17552 11144
rect 18512 11092 18564 11144
rect 19708 11135 19760 11144
rect 19708 11101 19717 11135
rect 19717 11101 19751 11135
rect 19751 11101 19760 11135
rect 19708 11092 19760 11101
rect 21088 11135 21140 11144
rect 19156 11024 19208 11076
rect 21088 11101 21097 11135
rect 21097 11101 21131 11135
rect 21131 11101 21140 11135
rect 21088 11092 21140 11101
rect 33692 11160 33744 11212
rect 36360 11228 36412 11280
rect 36452 11228 36504 11280
rect 36176 11203 36228 11212
rect 36176 11169 36185 11203
rect 36185 11169 36219 11203
rect 36219 11169 36228 11203
rect 36176 11160 36228 11169
rect 22192 11092 22244 11144
rect 23388 11092 23440 11144
rect 25780 11092 25832 11144
rect 33508 11135 33560 11144
rect 33508 11101 33514 11135
rect 33514 11101 33548 11135
rect 33548 11101 33560 11135
rect 33508 11092 33560 11101
rect 34428 11092 34480 11144
rect 35440 11092 35492 11144
rect 35716 11092 35768 11144
rect 35992 11135 36044 11144
rect 35992 11101 36001 11135
rect 36001 11101 36035 11135
rect 36035 11101 36044 11135
rect 35992 11092 36044 11101
rect 36452 11092 36504 11144
rect 36820 11135 36872 11144
rect 36820 11101 36829 11135
rect 36829 11101 36863 11135
rect 36863 11101 36872 11135
rect 36820 11092 36872 11101
rect 37004 11135 37056 11144
rect 37004 11101 37013 11135
rect 37013 11101 37047 11135
rect 37047 11101 37056 11135
rect 37004 11092 37056 11101
rect 40316 11203 40368 11212
rect 40316 11169 40325 11203
rect 40325 11169 40359 11203
rect 40359 11169 40368 11203
rect 40316 11160 40368 11169
rect 14556 10956 14608 11008
rect 17132 10999 17184 11008
rect 17132 10965 17141 10999
rect 17141 10965 17175 10999
rect 17175 10965 17184 10999
rect 17132 10956 17184 10965
rect 17316 10956 17368 11008
rect 19248 10956 19300 11008
rect 19432 10956 19484 11008
rect 20996 11024 21048 11076
rect 41420 11024 41472 11076
rect 42156 11067 42208 11076
rect 42156 11033 42165 11067
rect 42165 11033 42199 11067
rect 42199 11033 42208 11067
rect 42156 11024 42208 11033
rect 25688 10999 25740 11008
rect 25688 10965 25697 10999
rect 25697 10965 25731 10999
rect 25731 10965 25740 10999
rect 25688 10956 25740 10965
rect 33324 10999 33376 11008
rect 33324 10965 33333 10999
rect 33333 10965 33367 10999
rect 33367 10965 33376 10999
rect 33324 10956 33376 10965
rect 33416 10956 33468 11008
rect 35624 10999 35676 11008
rect 35624 10965 35633 10999
rect 35633 10965 35667 10999
rect 35667 10965 35676 10999
rect 35624 10956 35676 10965
rect 37556 10999 37608 11008
rect 37556 10965 37565 10999
rect 37565 10965 37599 10999
rect 37599 10965 37608 10999
rect 37556 10956 37608 10965
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 18696 10752 18748 10804
rect 18144 10727 18196 10736
rect 18144 10693 18153 10727
rect 18153 10693 18187 10727
rect 18187 10693 18196 10727
rect 18144 10684 18196 10693
rect 19248 10684 19300 10736
rect 21088 10752 21140 10804
rect 25780 10752 25832 10804
rect 28356 10795 28408 10804
rect 28356 10761 28365 10795
rect 28365 10761 28399 10795
rect 28399 10761 28408 10795
rect 28356 10752 28408 10761
rect 33324 10752 33376 10804
rect 35624 10752 35676 10804
rect 41420 10795 41472 10804
rect 41420 10761 41429 10795
rect 41429 10761 41463 10795
rect 41463 10761 41472 10795
rect 41420 10752 41472 10761
rect 1676 10659 1728 10668
rect 1676 10625 1685 10659
rect 1685 10625 1719 10659
rect 1719 10625 1728 10659
rect 1676 10616 1728 10625
rect 14096 10616 14148 10668
rect 14740 10659 14792 10668
rect 14740 10625 14749 10659
rect 14749 10625 14783 10659
rect 14783 10625 14792 10659
rect 14740 10616 14792 10625
rect 14832 10616 14884 10668
rect 18512 10659 18564 10668
rect 18512 10625 18521 10659
rect 18521 10625 18555 10659
rect 18555 10625 18564 10659
rect 18512 10616 18564 10625
rect 19064 10616 19116 10668
rect 19432 10659 19484 10668
rect 19432 10625 19441 10659
rect 19441 10625 19475 10659
rect 19475 10625 19484 10659
rect 19432 10616 19484 10625
rect 19984 10616 20036 10668
rect 30288 10684 30340 10736
rect 30472 10684 30524 10736
rect 35440 10684 35492 10736
rect 29920 10616 29972 10668
rect 30840 10616 30892 10668
rect 32588 10616 32640 10668
rect 33324 10616 33376 10668
rect 35348 10616 35400 10668
rect 35900 10616 35952 10668
rect 2044 10548 2096 10600
rect 2780 10591 2832 10600
rect 2780 10557 2789 10591
rect 2789 10557 2823 10591
rect 2823 10557 2832 10591
rect 2780 10548 2832 10557
rect 16948 10591 17000 10600
rect 16488 10480 16540 10532
rect 16948 10557 16957 10591
rect 16957 10557 16991 10591
rect 16991 10557 17000 10591
rect 16948 10548 17000 10557
rect 19156 10591 19208 10600
rect 19156 10557 19165 10591
rect 19165 10557 19199 10591
rect 19199 10557 19208 10591
rect 19156 10548 19208 10557
rect 22836 10591 22888 10600
rect 22836 10557 22845 10591
rect 22845 10557 22879 10591
rect 22879 10557 22888 10591
rect 22836 10548 22888 10557
rect 18052 10412 18104 10464
rect 18236 10480 18288 10532
rect 19248 10455 19300 10464
rect 19248 10421 19257 10455
rect 19257 10421 19291 10455
rect 19291 10421 19300 10455
rect 19248 10412 19300 10421
rect 28908 10591 28960 10600
rect 28908 10557 28917 10591
rect 28917 10557 28951 10591
rect 28951 10557 28960 10591
rect 33048 10591 33100 10600
rect 28908 10548 28960 10557
rect 33048 10557 33057 10591
rect 33057 10557 33091 10591
rect 33091 10557 33100 10591
rect 33048 10548 33100 10557
rect 37188 10616 37240 10668
rect 42248 10616 42300 10668
rect 36268 10548 36320 10600
rect 25320 10412 25372 10464
rect 30564 10412 30616 10464
rect 31116 10412 31168 10464
rect 32312 10412 32364 10464
rect 33048 10412 33100 10464
rect 35716 10455 35768 10464
rect 35716 10421 35725 10455
rect 35725 10421 35759 10455
rect 35759 10421 35768 10455
rect 35716 10412 35768 10421
rect 40316 10412 40368 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 2044 10251 2096 10260
rect 2044 10217 2053 10251
rect 2053 10217 2087 10251
rect 2087 10217 2096 10251
rect 2044 10208 2096 10217
rect 14832 10251 14884 10260
rect 14832 10217 14841 10251
rect 14841 10217 14875 10251
rect 14875 10217 14884 10251
rect 14832 10208 14884 10217
rect 15936 10208 15988 10260
rect 16488 10251 16540 10260
rect 16488 10217 16497 10251
rect 16497 10217 16531 10251
rect 16531 10217 16540 10251
rect 16488 10208 16540 10217
rect 17500 10208 17552 10260
rect 18236 10208 18288 10260
rect 18696 10251 18748 10260
rect 18696 10217 18705 10251
rect 18705 10217 18739 10251
rect 18739 10217 18748 10251
rect 18696 10208 18748 10217
rect 19984 10208 20036 10260
rect 22560 10251 22612 10260
rect 22560 10217 22569 10251
rect 22569 10217 22603 10251
rect 22603 10217 22612 10251
rect 22560 10208 22612 10217
rect 23480 10208 23532 10260
rect 32588 10251 32640 10260
rect 32588 10217 32597 10251
rect 32597 10217 32631 10251
rect 32631 10217 32640 10251
rect 32588 10208 32640 10217
rect 35348 10208 35400 10260
rect 36176 10140 36228 10192
rect 14740 10072 14792 10124
rect 16856 10072 16908 10124
rect 17316 10115 17368 10124
rect 17316 10081 17325 10115
rect 17325 10081 17359 10115
rect 17359 10081 17368 10115
rect 17316 10072 17368 10081
rect 19064 10072 19116 10124
rect 33048 10115 33100 10124
rect 2136 10047 2188 10056
rect 2136 10013 2145 10047
rect 2145 10013 2179 10047
rect 2179 10013 2188 10047
rect 2136 10004 2188 10013
rect 3240 10004 3292 10056
rect 15384 10004 15436 10056
rect 15476 9936 15528 9988
rect 15660 10004 15712 10056
rect 19248 10004 19300 10056
rect 33048 10081 33057 10115
rect 33057 10081 33091 10115
rect 33091 10081 33100 10115
rect 33048 10072 33100 10081
rect 33416 10072 33468 10124
rect 22192 10004 22244 10056
rect 22376 10047 22428 10056
rect 22376 10013 22385 10047
rect 22385 10013 22419 10047
rect 22419 10013 22428 10047
rect 22376 10004 22428 10013
rect 22560 10004 22612 10056
rect 25320 10004 25372 10056
rect 27344 10047 27396 10056
rect 27344 10013 27353 10047
rect 27353 10013 27387 10047
rect 27387 10013 27396 10047
rect 27344 10004 27396 10013
rect 30840 10004 30892 10056
rect 31484 10004 31536 10056
rect 33232 10004 33284 10056
rect 35440 10004 35492 10056
rect 35716 10047 35768 10056
rect 35716 10013 35725 10047
rect 35725 10013 35759 10047
rect 35759 10013 35768 10047
rect 35716 10004 35768 10013
rect 36820 10072 36872 10124
rect 40316 10115 40368 10124
rect 40316 10081 40325 10115
rect 40325 10081 40359 10115
rect 40359 10081 40368 10115
rect 40316 10072 40368 10081
rect 42156 10115 42208 10124
rect 42156 10081 42165 10115
rect 42165 10081 42199 10115
rect 42199 10081 42208 10115
rect 42156 10072 42208 10081
rect 37556 10004 37608 10056
rect 16120 9868 16172 9920
rect 16488 9911 16540 9920
rect 16488 9877 16513 9911
rect 16513 9877 16540 9911
rect 17960 9936 18012 9988
rect 19432 9936 19484 9988
rect 25688 9979 25740 9988
rect 25688 9945 25722 9979
rect 25722 9945 25740 9979
rect 25688 9936 25740 9945
rect 27620 9979 27672 9988
rect 27620 9945 27654 9979
rect 27654 9945 27672 9979
rect 27620 9936 27672 9945
rect 31116 9979 31168 9988
rect 31116 9945 31134 9979
rect 31134 9945 31168 9979
rect 31116 9936 31168 9945
rect 41420 9936 41472 9988
rect 16488 9868 16540 9877
rect 18236 9868 18288 9920
rect 21732 9911 21784 9920
rect 21732 9877 21741 9911
rect 21741 9877 21775 9911
rect 21775 9877 21784 9911
rect 21732 9868 21784 9877
rect 29552 9868 29604 9920
rect 30380 9868 30432 9920
rect 34704 9911 34756 9920
rect 34704 9877 34713 9911
rect 34713 9877 34747 9911
rect 34747 9877 34756 9911
rect 34704 9868 34756 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 18144 9664 18196 9716
rect 28908 9664 28960 9716
rect 29920 9664 29972 9716
rect 30564 9664 30616 9716
rect 15476 9596 15528 9648
rect 15660 9596 15712 9648
rect 4712 9528 4764 9580
rect 15384 9528 15436 9580
rect 16948 9596 17000 9648
rect 16304 9528 16356 9580
rect 18788 9596 18840 9648
rect 21732 9528 21784 9580
rect 22192 9528 22244 9580
rect 23572 9571 23624 9580
rect 23572 9537 23606 9571
rect 23606 9537 23624 9571
rect 25780 9596 25832 9648
rect 23572 9528 23624 9537
rect 15936 9460 15988 9512
rect 17132 9460 17184 9512
rect 18144 9503 18196 9512
rect 18144 9469 18153 9503
rect 18153 9469 18187 9503
rect 18187 9469 18196 9503
rect 18144 9460 18196 9469
rect 16120 9392 16172 9444
rect 18512 9460 18564 9512
rect 18696 9460 18748 9512
rect 18788 9392 18840 9444
rect 1768 9324 1820 9376
rect 2228 9367 2280 9376
rect 2228 9333 2237 9367
rect 2237 9333 2271 9367
rect 2271 9333 2280 9367
rect 2228 9324 2280 9333
rect 2872 9367 2924 9376
rect 2872 9333 2881 9367
rect 2881 9333 2915 9367
rect 2915 9333 2924 9367
rect 2872 9324 2924 9333
rect 22468 9460 22520 9512
rect 23020 9460 23072 9512
rect 22928 9392 22980 9444
rect 25504 9528 25556 9580
rect 27160 9596 27212 9648
rect 29184 9528 29236 9580
rect 30840 9596 30892 9648
rect 33324 9639 33376 9648
rect 33324 9605 33333 9639
rect 33333 9605 33367 9639
rect 33367 9605 33376 9639
rect 33324 9596 33376 9605
rect 34704 9596 34756 9648
rect 41420 9639 41472 9648
rect 41420 9605 41429 9639
rect 41429 9605 41463 9639
rect 41463 9605 41472 9639
rect 41420 9596 41472 9605
rect 30380 9571 30432 9580
rect 30380 9537 30389 9571
rect 30389 9537 30423 9571
rect 30423 9537 30432 9571
rect 30380 9528 30432 9537
rect 32312 9571 32364 9580
rect 32312 9537 32321 9571
rect 32321 9537 32355 9571
rect 32355 9537 32364 9571
rect 32312 9528 32364 9537
rect 34336 9528 34388 9580
rect 41144 9528 41196 9580
rect 26240 9460 26292 9512
rect 30564 9503 30616 9512
rect 30564 9469 30573 9503
rect 30573 9469 30607 9503
rect 30607 9469 30616 9503
rect 30564 9460 30616 9469
rect 33416 9460 33468 9512
rect 25136 9435 25188 9444
rect 25136 9401 25145 9435
rect 25145 9401 25179 9435
rect 25179 9401 25188 9435
rect 25136 9392 25188 9401
rect 27620 9392 27672 9444
rect 22652 9324 22704 9376
rect 22836 9367 22888 9376
rect 22836 9333 22845 9367
rect 22845 9333 22879 9367
rect 22879 9333 22888 9367
rect 22836 9324 22888 9333
rect 25228 9324 25280 9376
rect 32128 9367 32180 9376
rect 32128 9333 32137 9367
rect 32137 9333 32171 9367
rect 32171 9333 32180 9367
rect 32128 9324 32180 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 17960 9163 18012 9172
rect 17960 9129 17969 9163
rect 17969 9129 18003 9163
rect 18003 9129 18012 9163
rect 17960 9120 18012 9129
rect 17868 9052 17920 9104
rect 21548 9120 21600 9172
rect 22376 9120 22428 9172
rect 22560 9120 22612 9172
rect 29184 9120 29236 9172
rect 2228 8984 2280 9036
rect 3240 9027 3292 9036
rect 3240 8993 3249 9027
rect 3249 8993 3283 9027
rect 3283 8993 3292 9027
rect 3240 8984 3292 8993
rect 16488 9027 16540 9036
rect 1400 8959 1452 8968
rect 1400 8925 1409 8959
rect 1409 8925 1443 8959
rect 1443 8925 1452 8959
rect 1400 8916 1452 8925
rect 15384 8916 15436 8968
rect 16488 8993 16497 9027
rect 16497 8993 16531 9027
rect 16531 8993 16540 9027
rect 16488 8984 16540 8993
rect 21732 8984 21784 9036
rect 31484 9027 31536 9036
rect 31484 8993 31493 9027
rect 31493 8993 31527 9027
rect 31527 8993 31536 9027
rect 31484 8984 31536 8993
rect 15660 8959 15712 8968
rect 15660 8925 15669 8959
rect 15669 8925 15703 8959
rect 15703 8925 15712 8959
rect 15660 8916 15712 8925
rect 16120 8959 16172 8968
rect 16120 8925 16129 8959
rect 16129 8925 16163 8959
rect 16163 8925 16172 8959
rect 16120 8916 16172 8925
rect 16304 8959 16356 8968
rect 16304 8925 16313 8959
rect 16313 8925 16347 8959
rect 16347 8925 16356 8959
rect 16304 8916 16356 8925
rect 18052 8916 18104 8968
rect 20996 8916 21048 8968
rect 21548 8916 21600 8968
rect 20720 8848 20772 8900
rect 22652 8916 22704 8968
rect 25504 8916 25556 8968
rect 28632 8916 28684 8968
rect 29552 8959 29604 8968
rect 29552 8925 29561 8959
rect 29561 8925 29595 8959
rect 29595 8925 29604 8959
rect 29552 8916 29604 8925
rect 32128 8916 32180 8968
rect 26240 8848 26292 8900
rect 15568 8823 15620 8832
rect 15568 8789 15577 8823
rect 15577 8789 15611 8823
rect 15611 8789 15620 8823
rect 15568 8780 15620 8789
rect 19432 8780 19484 8832
rect 20628 8780 20680 8832
rect 23756 8780 23808 8832
rect 27160 8823 27212 8832
rect 27160 8789 27169 8823
rect 27169 8789 27203 8823
rect 27203 8789 27212 8823
rect 27160 8780 27212 8789
rect 29184 8780 29236 8832
rect 31300 8780 31352 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 16120 8619 16172 8628
rect 16120 8585 16129 8619
rect 16129 8585 16163 8619
rect 16163 8585 16172 8619
rect 16120 8576 16172 8585
rect 21548 8576 21600 8628
rect 22192 8619 22244 8628
rect 22192 8585 22201 8619
rect 22201 8585 22235 8619
rect 22235 8585 22244 8619
rect 22192 8576 22244 8585
rect 25228 8576 25280 8628
rect 28632 8619 28684 8628
rect 28632 8585 28641 8619
rect 28641 8585 28675 8619
rect 28675 8585 28684 8619
rect 28632 8576 28684 8585
rect 30564 8576 30616 8628
rect 2872 8508 2924 8560
rect 15568 8508 15620 8560
rect 16304 8508 16356 8560
rect 19432 8508 19484 8560
rect 1768 8483 1820 8492
rect 1768 8449 1777 8483
rect 1777 8449 1811 8483
rect 1811 8449 1820 8483
rect 1768 8440 1820 8449
rect 14740 8483 14792 8492
rect 14740 8449 14749 8483
rect 14749 8449 14783 8483
rect 14783 8449 14792 8483
rect 14740 8440 14792 8449
rect 17868 8440 17920 8492
rect 22836 8508 22888 8560
rect 27160 8508 27212 8560
rect 20720 8483 20772 8492
rect 20720 8449 20729 8483
rect 20729 8449 20763 8483
rect 20763 8449 20772 8483
rect 20720 8440 20772 8449
rect 20996 8483 21048 8492
rect 20996 8449 21005 8483
rect 21005 8449 21039 8483
rect 21039 8449 21048 8483
rect 20996 8440 21048 8449
rect 21732 8440 21784 8492
rect 22008 8483 22060 8492
rect 22008 8449 22017 8483
rect 22017 8449 22051 8483
rect 22051 8449 22060 8483
rect 22008 8440 22060 8449
rect 23020 8483 23072 8492
rect 23020 8449 23029 8483
rect 23029 8449 23063 8483
rect 23063 8449 23072 8483
rect 23020 8440 23072 8449
rect 27344 8440 27396 8492
rect 30840 8508 30892 8560
rect 29184 8440 29236 8492
rect 2780 8415 2832 8424
rect 2780 8381 2789 8415
rect 2789 8381 2823 8415
rect 2823 8381 2832 8415
rect 2780 8372 2832 8381
rect 17132 8372 17184 8424
rect 17408 8415 17460 8424
rect 17408 8381 17417 8415
rect 17417 8381 17451 8415
rect 17451 8381 17460 8415
rect 17408 8372 17460 8381
rect 30288 8372 30340 8424
rect 17224 8236 17276 8288
rect 18604 8236 18656 8288
rect 20260 8304 20312 8356
rect 31300 8347 31352 8356
rect 31300 8313 31309 8347
rect 31309 8313 31343 8347
rect 31343 8313 31352 8347
rect 31300 8304 31352 8313
rect 19156 8236 19208 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 15660 8032 15712 8084
rect 16304 8032 16356 8084
rect 17868 8032 17920 8084
rect 20628 8075 20680 8084
rect 20628 8041 20637 8075
rect 20637 8041 20671 8075
rect 20671 8041 20680 8075
rect 20628 8032 20680 8041
rect 22008 8032 22060 8084
rect 23572 8032 23624 8084
rect 15936 7939 15988 7948
rect 15936 7905 15945 7939
rect 15945 7905 15979 7939
rect 15979 7905 15988 7939
rect 15936 7896 15988 7905
rect 16856 7939 16908 7948
rect 16856 7905 16865 7939
rect 16865 7905 16899 7939
rect 16899 7905 16908 7939
rect 16856 7896 16908 7905
rect 16120 7828 16172 7880
rect 23020 7896 23072 7948
rect 25320 7939 25372 7948
rect 25320 7905 25329 7939
rect 25329 7905 25363 7939
rect 25363 7905 25372 7939
rect 25320 7896 25372 7905
rect 22928 7871 22980 7880
rect 22928 7837 22937 7871
rect 22937 7837 22971 7871
rect 22971 7837 22980 7871
rect 22928 7828 22980 7837
rect 23756 7871 23808 7880
rect 23756 7837 23765 7871
rect 23765 7837 23799 7871
rect 23799 7837 23808 7871
rect 23756 7828 23808 7837
rect 41604 7828 41656 7880
rect 17132 7803 17184 7812
rect 17132 7769 17166 7803
rect 17166 7769 17184 7803
rect 17132 7760 17184 7769
rect 18788 7760 18840 7812
rect 20720 7760 20772 7812
rect 25596 7803 25648 7812
rect 25596 7769 25630 7803
rect 25630 7769 25648 7803
rect 25596 7760 25648 7769
rect 23572 7735 23624 7744
rect 23572 7701 23581 7735
rect 23581 7701 23615 7735
rect 23615 7701 23624 7735
rect 23572 7692 23624 7701
rect 40500 7692 40552 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 17868 7488 17920 7540
rect 18788 7531 18840 7540
rect 18788 7497 18797 7531
rect 18797 7497 18831 7531
rect 18831 7497 18840 7531
rect 18788 7488 18840 7497
rect 17224 7420 17276 7472
rect 23572 7420 23624 7472
rect 17408 7395 17460 7404
rect 17408 7361 17417 7395
rect 17417 7361 17451 7395
rect 17451 7361 17460 7395
rect 18604 7395 18656 7404
rect 17408 7352 17460 7361
rect 18604 7361 18613 7395
rect 18613 7361 18647 7395
rect 18647 7361 18656 7395
rect 18604 7352 18656 7361
rect 20628 7352 20680 7404
rect 23020 7395 23072 7404
rect 23020 7361 23029 7395
rect 23029 7361 23063 7395
rect 23063 7361 23072 7395
rect 23020 7352 23072 7361
rect 25596 7488 25648 7540
rect 25504 7352 25556 7404
rect 41880 7395 41932 7404
rect 41880 7361 41889 7395
rect 41889 7361 41923 7395
rect 41923 7361 41932 7395
rect 41880 7352 41932 7361
rect 20996 7284 21048 7336
rect 17132 7259 17184 7268
rect 17132 7225 17141 7259
rect 17141 7225 17175 7259
rect 17175 7225 17184 7259
rect 17132 7216 17184 7225
rect 24584 7216 24636 7268
rect 40960 7191 41012 7200
rect 40960 7157 40969 7191
rect 40969 7157 41003 7191
rect 41003 7157 41012 7191
rect 40960 7148 41012 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 4068 6808 4120 6860
rect 13636 6808 13688 6860
rect 40960 6808 41012 6860
rect 4620 6740 4672 6792
rect 20260 6783 20312 6792
rect 20260 6749 20269 6783
rect 20269 6749 20303 6783
rect 20303 6749 20312 6783
rect 20260 6740 20312 6749
rect 40500 6715 40552 6724
rect 40500 6681 40509 6715
rect 40509 6681 40543 6715
rect 40543 6681 40552 6715
rect 40500 6672 40552 6681
rect 42156 6715 42208 6724
rect 42156 6681 42165 6715
rect 42165 6681 42199 6715
rect 42199 6681 42208 6715
rect 42156 6672 42208 6681
rect 4160 6647 4212 6656
rect 4160 6613 4169 6647
rect 4169 6613 4203 6647
rect 4203 6613 4212 6647
rect 4160 6604 4212 6613
rect 20720 6604 20772 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 7656 6400 7708 6452
rect 4160 6375 4212 6384
rect 4160 6341 4169 6375
rect 4169 6341 4203 6375
rect 4203 6341 4212 6375
rect 4160 6332 4212 6341
rect 3976 6239 4028 6248
rect 3976 6205 3985 6239
rect 3985 6205 4019 6239
rect 4019 6205 4028 6239
rect 3976 6196 4028 6205
rect 5080 6239 5132 6248
rect 5080 6205 5089 6239
rect 5089 6205 5123 6239
rect 5123 6205 5132 6239
rect 5080 6196 5132 6205
rect 1400 6103 1452 6112
rect 1400 6069 1409 6103
rect 1409 6069 1443 6103
rect 1443 6069 1452 6103
rect 1400 6060 1452 6069
rect 1952 6060 2004 6112
rect 2780 6103 2832 6112
rect 2780 6069 2789 6103
rect 2789 6069 2823 6103
rect 2823 6069 2832 6103
rect 2780 6060 2832 6069
rect 40316 6060 40368 6112
rect 41788 6103 41840 6112
rect 41788 6069 41797 6103
rect 41797 6069 41831 6103
rect 41831 6069 41840 6103
rect 41788 6060 41840 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 3976 5856 4028 5908
rect 1400 5763 1452 5772
rect 1400 5729 1409 5763
rect 1409 5729 1443 5763
rect 1443 5729 1452 5763
rect 1400 5720 1452 5729
rect 1860 5763 1912 5772
rect 1860 5729 1869 5763
rect 1869 5729 1903 5763
rect 1903 5729 1912 5763
rect 1860 5720 1912 5729
rect 2136 5720 2188 5772
rect 4988 5652 5040 5704
rect 41696 5720 41748 5772
rect 38476 5652 38528 5704
rect 39856 5695 39908 5704
rect 39856 5661 39865 5695
rect 39865 5661 39899 5695
rect 39899 5661 39908 5695
rect 39856 5652 39908 5661
rect 41236 5652 41288 5704
rect 41972 5695 42024 5704
rect 41972 5661 41981 5695
rect 41981 5661 42015 5695
rect 42015 5661 42024 5695
rect 41972 5652 42024 5661
rect 1584 5627 1636 5636
rect 1584 5593 1593 5627
rect 1593 5593 1627 5627
rect 1627 5593 1636 5627
rect 1584 5584 1636 5593
rect 38660 5516 38712 5568
rect 41972 5516 42024 5568
rect 42064 5559 42116 5568
rect 42064 5525 42073 5559
rect 42073 5525 42107 5559
rect 42107 5525 42116 5559
rect 42064 5516 42116 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 2780 5244 2832 5296
rect 38660 5287 38712 5296
rect 38660 5253 38669 5287
rect 38669 5253 38703 5287
rect 38703 5253 38712 5287
rect 38660 5244 38712 5253
rect 1952 5219 2004 5228
rect 1952 5185 1961 5219
rect 1961 5185 1995 5219
rect 1995 5185 2004 5219
rect 1952 5176 2004 5185
rect 38476 5219 38528 5228
rect 38476 5185 38485 5219
rect 38485 5185 38519 5219
rect 38519 5185 38528 5219
rect 38476 5176 38528 5185
rect 41052 5176 41104 5228
rect 41420 5219 41472 5228
rect 41420 5185 41429 5219
rect 41429 5185 41463 5219
rect 41463 5185 41472 5219
rect 41420 5176 41472 5185
rect 2780 5151 2832 5160
rect 2780 5117 2789 5151
rect 2789 5117 2823 5151
rect 2823 5117 2832 5151
rect 2780 5108 2832 5117
rect 43168 5108 43220 5160
rect 4620 4972 4672 5024
rect 40040 4972 40092 5024
rect 41512 5015 41564 5024
rect 41512 4981 41521 5015
rect 41521 4981 41555 5015
rect 41555 4981 41564 5015
rect 41512 4972 41564 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 1584 4768 1636 4820
rect 4804 4700 4856 4752
rect 1492 4564 1544 4616
rect 2136 4564 2188 4616
rect 5540 4632 5592 4684
rect 40316 4675 40368 4684
rect 40316 4641 40325 4675
rect 40325 4641 40359 4675
rect 40359 4641 40368 4675
rect 40316 4632 40368 4641
rect 41512 4632 41564 4684
rect 41880 4675 41932 4684
rect 41880 4641 41889 4675
rect 41889 4641 41923 4675
rect 41923 4641 41932 4675
rect 41880 4632 41932 4641
rect 3240 4564 3292 4616
rect 4712 4564 4764 4616
rect 36728 4607 36780 4616
rect 36728 4573 36737 4607
rect 36737 4573 36771 4607
rect 36771 4573 36780 4607
rect 36728 4564 36780 4573
rect 37556 4564 37608 4616
rect 39028 4564 39080 4616
rect 39120 4607 39172 4616
rect 39120 4573 39129 4607
rect 39129 4573 39163 4607
rect 39163 4573 39172 4607
rect 39120 4564 39172 4573
rect 5172 4496 5224 4548
rect 11244 4496 11296 4548
rect 4804 4428 4856 4480
rect 39764 4428 39816 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 10140 4156 10192 4208
rect 18604 4156 18656 4208
rect 39764 4199 39816 4208
rect 39764 4165 39773 4199
rect 39773 4165 39807 4199
rect 39807 4165 39816 4199
rect 39764 4156 39816 4165
rect 2412 4088 2464 4140
rect 3148 4131 3200 4140
rect 3148 4097 3157 4131
rect 3157 4097 3191 4131
rect 3191 4097 3200 4131
rect 3148 4088 3200 4097
rect 4988 4131 5040 4140
rect 4988 4097 4997 4131
rect 4997 4097 5031 4131
rect 5031 4097 5040 4131
rect 4988 4088 5040 4097
rect 37832 4131 37884 4140
rect 4804 4063 4856 4072
rect 4804 4029 4813 4063
rect 4813 4029 4847 4063
rect 4847 4029 4856 4063
rect 4804 4020 4856 4029
rect 7564 4020 7616 4072
rect 10140 4020 10192 4072
rect 10232 4020 10284 4072
rect 11428 4020 11480 4072
rect 10692 3952 10744 4004
rect 37832 4097 37841 4131
rect 37841 4097 37875 4131
rect 37875 4097 37884 4131
rect 37832 4088 37884 4097
rect 22468 4020 22520 4072
rect 22836 4063 22888 4072
rect 22836 4029 22845 4063
rect 22845 4029 22879 4063
rect 22879 4029 22888 4063
rect 22836 4020 22888 4029
rect 23204 4063 23256 4072
rect 23204 4029 23213 4063
rect 23213 4029 23247 4063
rect 23247 4029 23256 4063
rect 23204 4020 23256 4029
rect 39028 4088 39080 4140
rect 39120 4020 39172 4072
rect 41328 4063 41380 4072
rect 41328 4029 41337 4063
rect 41337 4029 41371 4063
rect 41371 4029 41380 4063
rect 41328 4020 41380 4029
rect 3056 3884 3108 3936
rect 4896 3884 4948 3936
rect 6368 3927 6420 3936
rect 6368 3893 6377 3927
rect 6377 3893 6411 3927
rect 6411 3893 6420 3927
rect 6368 3884 6420 3893
rect 9864 3927 9916 3936
rect 9864 3893 9873 3927
rect 9873 3893 9907 3927
rect 9907 3893 9916 3927
rect 9864 3884 9916 3893
rect 11336 3884 11388 3936
rect 11520 3927 11572 3936
rect 11520 3893 11529 3927
rect 11529 3893 11563 3927
rect 11563 3893 11572 3927
rect 11520 3884 11572 3893
rect 18144 3927 18196 3936
rect 18144 3893 18153 3927
rect 18153 3893 18187 3927
rect 18187 3893 18196 3927
rect 18144 3884 18196 3893
rect 19524 3884 19576 3936
rect 21824 3884 21876 3936
rect 34704 3927 34756 3936
rect 34704 3893 34713 3927
rect 34713 3893 34747 3927
rect 34747 3893 34756 3927
rect 34704 3884 34756 3893
rect 35624 3927 35676 3936
rect 35624 3893 35633 3927
rect 35633 3893 35667 3927
rect 35667 3893 35676 3927
rect 35624 3884 35676 3893
rect 37464 3884 37516 3936
rect 37648 3884 37700 3936
rect 38660 3927 38712 3936
rect 38660 3893 38669 3927
rect 38669 3893 38703 3927
rect 38703 3893 38712 3927
rect 38660 3884 38712 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 8116 3680 8168 3732
rect 3056 3587 3108 3596
rect 3056 3553 3065 3587
rect 3065 3553 3099 3587
rect 3099 3553 3108 3587
rect 3056 3544 3108 3553
rect 3240 3587 3292 3596
rect 3240 3553 3249 3587
rect 3249 3553 3283 3587
rect 3283 3553 3292 3587
rect 3240 3544 3292 3553
rect 4712 3587 4764 3596
rect 4712 3553 4721 3587
rect 4721 3553 4755 3587
rect 4755 3553 4764 3587
rect 4712 3544 4764 3553
rect 4896 3587 4948 3596
rect 4896 3553 4905 3587
rect 4905 3553 4939 3587
rect 4939 3553 4948 3587
rect 4896 3544 4948 3553
rect 5172 3587 5224 3596
rect 5172 3553 5181 3587
rect 5181 3553 5215 3587
rect 5215 3553 5224 3587
rect 5172 3544 5224 3553
rect 9864 3612 9916 3664
rect 9220 3587 9272 3596
rect 9220 3553 9229 3587
rect 9229 3553 9263 3587
rect 9263 3553 9272 3587
rect 9220 3544 9272 3553
rect 9680 3587 9732 3596
rect 9680 3553 9689 3587
rect 9689 3553 9723 3587
rect 9723 3553 9732 3587
rect 9680 3544 9732 3553
rect 11336 3587 11388 3596
rect 11336 3553 11345 3587
rect 11345 3553 11379 3587
rect 11379 3553 11388 3587
rect 11336 3544 11388 3553
rect 11704 3544 11756 3596
rect 16856 3680 16908 3732
rect 22468 3723 22520 3732
rect 22468 3689 22477 3723
rect 22477 3689 22511 3723
rect 22511 3689 22520 3723
rect 22468 3680 22520 3689
rect 16672 3544 16724 3596
rect 16856 3587 16908 3596
rect 16856 3553 16865 3587
rect 16865 3553 16899 3587
rect 16899 3553 16908 3587
rect 16856 3544 16908 3553
rect 19524 3587 19576 3596
rect 19524 3553 19533 3587
rect 19533 3553 19567 3587
rect 19567 3553 19576 3587
rect 19524 3544 19576 3553
rect 19984 3587 20036 3596
rect 19984 3553 19993 3587
rect 19993 3553 20027 3587
rect 20027 3553 20036 3587
rect 19984 3544 20036 3553
rect 1400 3519 1452 3528
rect 1400 3485 1409 3519
rect 1409 3485 1443 3519
rect 1443 3485 1452 3519
rect 1400 3476 1452 3485
rect 4252 3519 4304 3528
rect 4252 3485 4261 3519
rect 4261 3485 4295 3519
rect 4295 3485 4304 3519
rect 4252 3476 4304 3485
rect 7196 3476 7248 3528
rect 5356 3340 5408 3392
rect 7380 3340 7432 3392
rect 14280 3476 14332 3528
rect 18604 3519 18656 3528
rect 18604 3485 18613 3519
rect 18613 3485 18647 3519
rect 18647 3485 18656 3519
rect 18604 3476 18656 3485
rect 11612 3408 11664 3460
rect 16764 3408 16816 3460
rect 12164 3340 12216 3392
rect 16948 3340 17000 3392
rect 18328 3340 18380 3392
rect 23480 3476 23532 3528
rect 34704 3587 34756 3596
rect 34704 3553 34713 3587
rect 34713 3553 34747 3587
rect 34747 3553 34756 3587
rect 34704 3544 34756 3553
rect 34888 3544 34940 3596
rect 36728 3544 36780 3596
rect 37372 3544 37424 3596
rect 41788 3544 41840 3596
rect 27620 3476 27672 3528
rect 27804 3519 27856 3528
rect 27804 3485 27813 3519
rect 27813 3485 27847 3519
rect 27847 3485 27856 3519
rect 27804 3476 27856 3485
rect 20536 3408 20588 3460
rect 23664 3383 23716 3392
rect 23664 3349 23673 3383
rect 23673 3349 23707 3383
rect 23707 3349 23716 3383
rect 23664 3340 23716 3349
rect 35532 3408 35584 3460
rect 37188 3451 37240 3460
rect 37188 3417 37197 3451
rect 37197 3417 37231 3451
rect 37231 3417 37240 3451
rect 37188 3408 37240 3417
rect 39764 3408 39816 3460
rect 41972 3451 42024 3460
rect 41972 3417 41981 3451
rect 41981 3417 42015 3451
rect 42015 3417 42024 3451
rect 41972 3408 42024 3417
rect 36360 3340 36412 3392
rect 41236 3340 41288 3392
rect 42156 3340 42208 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 4252 3136 4304 3188
rect 664 3068 716 3120
rect 5356 3111 5408 3120
rect 5356 3077 5365 3111
rect 5365 3077 5399 3111
rect 5399 3077 5408 3111
rect 5356 3068 5408 3077
rect 1400 3043 1452 3052
rect 1400 3009 1409 3043
rect 1409 3009 1443 3043
rect 1443 3009 1452 3043
rect 1400 3000 1452 3009
rect 5540 3043 5592 3052
rect 5540 3009 5549 3043
rect 5549 3009 5583 3043
rect 5583 3009 5592 3043
rect 9588 3136 9640 3188
rect 12072 3136 12124 3188
rect 16764 3179 16816 3188
rect 7380 3111 7432 3120
rect 7380 3077 7389 3111
rect 7389 3077 7423 3111
rect 7423 3077 7432 3111
rect 7380 3068 7432 3077
rect 5540 3000 5592 3009
rect 7196 3043 7248 3052
rect 7196 3009 7205 3043
rect 7205 3009 7239 3043
rect 7239 3009 7248 3043
rect 7196 3000 7248 3009
rect 10232 3043 10284 3052
rect 10232 3009 10241 3043
rect 10241 3009 10275 3043
rect 10275 3009 10284 3043
rect 10232 3000 10284 3009
rect 12256 3068 12308 3120
rect 16764 3145 16773 3179
rect 16773 3145 16807 3179
rect 16807 3145 16816 3179
rect 16764 3136 16816 3145
rect 16948 3136 17000 3188
rect 20536 3179 20588 3188
rect 18328 3111 18380 3120
rect 11520 3043 11572 3052
rect 11520 3009 11529 3043
rect 11529 3009 11563 3043
rect 11563 3009 11572 3043
rect 11520 3000 11572 3009
rect 14280 3043 14332 3052
rect 14280 3009 14289 3043
rect 14289 3009 14323 3043
rect 14323 3009 14332 3043
rect 14280 3000 14332 3009
rect 18328 3077 18337 3111
rect 18337 3077 18371 3111
rect 18371 3077 18380 3111
rect 18328 3068 18380 3077
rect 20536 3145 20545 3179
rect 20545 3145 20579 3179
rect 20579 3145 20588 3179
rect 20536 3136 20588 3145
rect 22836 3136 22888 3188
rect 23664 3111 23716 3120
rect 18144 3043 18196 3052
rect 1584 2975 1636 2984
rect 1584 2941 1593 2975
rect 1593 2941 1627 2975
rect 1627 2941 1636 2975
rect 1584 2932 1636 2941
rect 2780 2975 2832 2984
rect 2780 2941 2789 2975
rect 2789 2941 2823 2975
rect 2823 2941 2832 2975
rect 2780 2932 2832 2941
rect 7104 2932 7156 2984
rect 3240 2864 3292 2916
rect 9128 2864 9180 2916
rect 10968 2864 11020 2916
rect 15200 2932 15252 2984
rect 15476 2975 15528 2984
rect 15476 2941 15485 2975
rect 15485 2941 15519 2975
rect 15519 2941 15528 2975
rect 15476 2932 15528 2941
rect 18144 3009 18153 3043
rect 18153 3009 18187 3043
rect 18187 3009 18196 3043
rect 18144 3000 18196 3009
rect 20628 3043 20680 3052
rect 20628 3009 20637 3043
rect 20637 3009 20671 3043
rect 20671 3009 20680 3043
rect 20628 3000 20680 3009
rect 23664 3077 23673 3111
rect 23673 3077 23707 3111
rect 23707 3077 23716 3111
rect 23664 3068 23716 3077
rect 23480 3043 23532 3052
rect 18696 2975 18748 2984
rect 18696 2941 18705 2975
rect 18705 2941 18739 2975
rect 18739 2941 18748 2975
rect 18696 2932 18748 2941
rect 23480 3009 23489 3043
rect 23489 3009 23523 3043
rect 23523 3009 23532 3043
rect 23480 3000 23532 3009
rect 27804 3043 27856 3052
rect 27804 3009 27813 3043
rect 27813 3009 27847 3043
rect 27847 3009 27856 3043
rect 27804 3000 27856 3009
rect 35624 3068 35676 3120
rect 38660 3068 38712 3120
rect 40040 3111 40092 3120
rect 40040 3077 40049 3111
rect 40049 3077 40083 3111
rect 40083 3077 40092 3111
rect 40040 3068 40092 3077
rect 37556 3043 37608 3052
rect 37556 3009 37565 3043
rect 37565 3009 37599 3043
rect 37599 3009 37608 3043
rect 37556 3000 37608 3009
rect 39856 3043 39908 3052
rect 39856 3009 39865 3043
rect 39865 3009 39899 3043
rect 39899 3009 39908 3043
rect 39856 3000 39908 3009
rect 23848 2932 23900 2984
rect 27988 2975 28040 2984
rect 27988 2941 27997 2975
rect 27997 2941 28031 2975
rect 28031 2941 28040 2975
rect 27988 2932 28040 2941
rect 28356 2975 28408 2984
rect 28356 2941 28365 2975
rect 28365 2941 28399 2975
rect 28399 2941 28408 2975
rect 28356 2932 28408 2941
rect 35808 2932 35860 2984
rect 36084 2975 36136 2984
rect 36084 2941 36093 2975
rect 36093 2941 36127 2975
rect 36127 2941 36136 2975
rect 36084 2932 36136 2941
rect 39304 2975 39356 2984
rect 39304 2941 39313 2975
rect 39313 2941 39347 2975
rect 39347 2941 39356 2975
rect 39304 2932 39356 2941
rect 40592 2975 40644 2984
rect 40592 2941 40601 2975
rect 40601 2941 40635 2975
rect 40635 2941 40644 2975
rect 40592 2932 40644 2941
rect 35440 2864 35492 2916
rect 38936 2864 38988 2916
rect 6552 2796 6604 2848
rect 10784 2796 10836 2848
rect 22008 2839 22060 2848
rect 22008 2805 22017 2839
rect 22017 2805 22051 2839
rect 22051 2805 22060 2839
rect 22008 2796 22060 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 1584 2592 1636 2644
rect 3424 2592 3476 2644
rect 11612 2635 11664 2644
rect 4620 2524 4672 2576
rect 6828 2524 6880 2576
rect 3976 2456 4028 2508
rect 6368 2499 6420 2508
rect 6368 2465 6377 2499
rect 6377 2465 6411 2499
rect 6411 2465 6420 2499
rect 6368 2456 6420 2465
rect 6552 2499 6604 2508
rect 6552 2465 6561 2499
rect 6561 2465 6595 2499
rect 6595 2465 6604 2499
rect 6552 2456 6604 2465
rect 6736 2456 6788 2508
rect 9128 2499 9180 2508
rect 9128 2465 9137 2499
rect 9137 2465 9171 2499
rect 9171 2465 9180 2499
rect 9128 2456 9180 2465
rect 2136 2431 2188 2440
rect 2136 2397 2145 2431
rect 2145 2397 2179 2431
rect 2179 2397 2188 2431
rect 2136 2388 2188 2397
rect 2964 2388 3016 2440
rect 10784 2499 10836 2508
rect 10784 2465 10793 2499
rect 10793 2465 10827 2499
rect 10827 2465 10836 2499
rect 10784 2456 10836 2465
rect 11612 2601 11621 2635
rect 11621 2601 11655 2635
rect 11655 2601 11664 2635
rect 11612 2592 11664 2601
rect 15200 2635 15252 2644
rect 15200 2601 15209 2635
rect 15209 2601 15243 2635
rect 15243 2601 15252 2635
rect 15200 2592 15252 2601
rect 27988 2592 28040 2644
rect 35808 2635 35860 2644
rect 35808 2601 35817 2635
rect 35817 2601 35851 2635
rect 35851 2601 35860 2635
rect 35808 2592 35860 2601
rect 37188 2592 37240 2644
rect 13728 2456 13780 2508
rect 21824 2499 21876 2508
rect 10692 2320 10744 2372
rect 11428 2388 11480 2440
rect 20628 2388 20680 2440
rect 21824 2465 21833 2499
rect 21833 2465 21867 2499
rect 21867 2465 21876 2499
rect 21824 2456 21876 2465
rect 22008 2499 22060 2508
rect 22008 2465 22017 2499
rect 22017 2465 22051 2499
rect 22051 2465 22060 2499
rect 22008 2456 22060 2465
rect 22560 2499 22612 2508
rect 22560 2465 22569 2499
rect 22569 2465 22603 2499
rect 22603 2465 22612 2499
rect 22560 2456 22612 2465
rect 41420 2524 41472 2576
rect 37464 2499 37516 2508
rect 37464 2465 37473 2499
rect 37473 2465 37507 2499
rect 37507 2465 37516 2499
rect 37464 2456 37516 2465
rect 37648 2499 37700 2508
rect 37648 2465 37657 2499
rect 37657 2465 37691 2499
rect 37691 2465 37700 2499
rect 37648 2456 37700 2465
rect 41328 2499 41380 2508
rect 41328 2465 41337 2499
rect 41337 2465 41371 2499
rect 41371 2465 41380 2499
rect 41328 2456 41380 2465
rect 42064 2456 42116 2508
rect 27620 2388 27672 2440
rect 35900 2431 35952 2440
rect 35900 2397 35909 2431
rect 35909 2397 35943 2431
rect 35943 2397 35952 2431
rect 36360 2431 36412 2440
rect 35900 2388 35952 2397
rect 36360 2397 36369 2431
rect 36369 2397 36403 2431
rect 36403 2397 36412 2431
rect 36360 2388 36412 2397
rect 37832 2320 37884 2372
rect 39948 2320 40000 2372
rect 41696 2320 41748 2372
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 10232 2048 10284 2100
rect 35900 2048 35952 2100
<< metal2 >>
rect 18 43200 74 44000
rect 662 43200 718 44000
rect 1950 43330 2006 44000
rect 2594 43330 2650 44000
rect 1950 43302 2084 43330
rect 1950 43200 2006 43302
rect 1860 41132 1912 41138
rect 1860 41074 1912 41080
rect 1872 40905 1900 41074
rect 1858 40896 1914 40905
rect 1858 40831 1914 40840
rect 2056 40594 2084 43302
rect 2594 43302 2728 43330
rect 2594 43200 2650 43302
rect 2700 41002 2728 43302
rect 3238 43200 3294 44000
rect 4526 43330 4582 44000
rect 5170 43330 5226 44000
rect 4526 43302 4936 43330
rect 4526 43200 4582 43302
rect 2870 42936 2926 42945
rect 2870 42871 2926 42880
rect 2688 40996 2740 41002
rect 2688 40938 2740 40944
rect 2780 40928 2832 40934
rect 2780 40870 2832 40876
rect 2044 40588 2096 40594
rect 2044 40530 2096 40536
rect 2792 40118 2820 40870
rect 2780 40112 2832 40118
rect 2780 40054 2832 40060
rect 1584 39976 1636 39982
rect 1584 39918 1636 39924
rect 1400 39432 1452 39438
rect 1400 39374 1452 39380
rect 1412 38554 1440 39374
rect 1596 38962 1624 39918
rect 2884 39506 2912 42871
rect 2962 41576 3018 41585
rect 2962 41511 3018 41520
rect 2872 39500 2924 39506
rect 2872 39442 2924 39448
rect 2136 39364 2188 39370
rect 2136 39306 2188 39312
rect 2148 39098 2176 39306
rect 2136 39092 2188 39098
rect 2136 39034 2188 39040
rect 1584 38956 1636 38962
rect 1584 38898 1636 38904
rect 2412 38888 2464 38894
rect 2412 38830 2464 38836
rect 1400 38548 1452 38554
rect 1400 38490 1452 38496
rect 1676 37664 1728 37670
rect 1676 37606 1728 37612
rect 1688 37330 1716 37606
rect 1676 37324 1728 37330
rect 1676 37266 1728 37272
rect 2044 37188 2096 37194
rect 2044 37130 2096 37136
rect 2056 36922 2084 37130
rect 2044 36916 2096 36922
rect 2044 36858 2096 36864
rect 2228 36848 2280 36854
rect 2228 36790 2280 36796
rect 1952 36168 2004 36174
rect 1952 36110 2004 36116
rect 1964 35698 1992 36110
rect 2240 35894 2268 36790
rect 2240 35866 2360 35894
rect 1952 35692 2004 35698
rect 1952 35634 2004 35640
rect 1676 28960 1728 28966
rect 1676 28902 1728 28908
rect 1688 28626 1716 28902
rect 1676 28620 1728 28626
rect 1676 28562 1728 28568
rect 2136 28484 2188 28490
rect 2136 28426 2188 28432
rect 2148 28218 2176 28426
rect 2136 28212 2188 28218
rect 2136 28154 2188 28160
rect 1400 23112 1452 23118
rect 1400 23054 1452 23060
rect 1412 22098 1440 23054
rect 2136 22636 2188 22642
rect 2136 22578 2188 22584
rect 1584 22432 1636 22438
rect 1584 22374 1636 22380
rect 1596 22098 1624 22374
rect 1400 22092 1452 22098
rect 1400 22034 1452 22040
rect 1584 22092 1636 22098
rect 1584 22034 1636 22040
rect 1860 22092 1912 22098
rect 1860 22034 1912 22040
rect 1872 21865 1900 22034
rect 1858 21856 1914 21865
rect 1858 21791 1914 21800
rect 1860 21480 1912 21486
rect 1860 21422 1912 21428
rect 1872 21146 1900 21422
rect 1860 21140 1912 21146
rect 1860 21082 1912 21088
rect 1400 20256 1452 20262
rect 1400 20198 1452 20204
rect 1412 19922 1440 20198
rect 1400 19916 1452 19922
rect 1400 19858 1452 19864
rect 1860 19916 1912 19922
rect 1860 19858 1912 19864
rect 1872 19825 1900 19858
rect 1858 19816 1914 19825
rect 1858 19751 1914 19760
rect 2044 19780 2096 19786
rect 2044 19722 2096 19728
rect 2056 19514 2084 19722
rect 2044 19508 2096 19514
rect 2044 19450 2096 19456
rect 2148 19378 2176 22578
rect 2136 19372 2188 19378
rect 2136 19314 2188 19320
rect 2148 19258 2176 19314
rect 2056 19230 2176 19258
rect 1952 17672 2004 17678
rect 1952 17614 2004 17620
rect 1964 17202 1992 17614
rect 1952 17196 2004 17202
rect 1952 17138 2004 17144
rect 1860 16652 1912 16658
rect 1860 16594 1912 16600
rect 1400 16584 1452 16590
rect 1400 16526 1452 16532
rect 1412 16114 1440 16526
rect 1872 16425 1900 16594
rect 1858 16416 1914 16425
rect 1858 16351 1914 16360
rect 1400 16108 1452 16114
rect 1400 16050 1452 16056
rect 1768 15496 1820 15502
rect 1768 15438 1820 15444
rect 1780 15026 1808 15438
rect 1768 15020 1820 15026
rect 1768 14962 1820 14968
rect 1952 13864 2004 13870
rect 1952 13806 2004 13812
rect 1964 13530 1992 13806
rect 1952 13524 2004 13530
rect 1952 13466 2004 13472
rect 1676 12640 1728 12646
rect 1676 12582 1728 12588
rect 1688 12306 1716 12582
rect 1676 12300 1728 12306
rect 1676 12242 1728 12248
rect 2056 11234 2084 19230
rect 2136 17536 2188 17542
rect 2136 17478 2188 17484
rect 2148 17270 2176 17478
rect 2136 17264 2188 17270
rect 2136 17206 2188 17212
rect 2136 16516 2188 16522
rect 2136 16458 2188 16464
rect 2148 16250 2176 16458
rect 2136 16244 2188 16250
rect 2136 16186 2188 16192
rect 2228 14952 2280 14958
rect 2228 14894 2280 14900
rect 2240 14618 2268 14894
rect 2228 14612 2280 14618
rect 2228 14554 2280 14560
rect 2136 12164 2188 12170
rect 2136 12106 2188 12112
rect 2148 11898 2176 12106
rect 2136 11892 2188 11898
rect 2136 11834 2188 11840
rect 2332 11762 2360 35866
rect 2320 11756 2372 11762
rect 2320 11698 2372 11704
rect 2056 11206 2176 11234
rect 1676 11144 1728 11150
rect 1676 11086 1728 11092
rect 1688 10674 1716 11086
rect 1676 10668 1728 10674
rect 1676 10610 1728 10616
rect 2044 10600 2096 10606
rect 2044 10542 2096 10548
rect 2056 10266 2084 10542
rect 2044 10260 2096 10266
rect 2044 10202 2096 10208
rect 2148 10062 2176 11206
rect 2136 10056 2188 10062
rect 2136 9998 2188 10004
rect 1768 9376 1820 9382
rect 1768 9318 1820 9324
rect 1400 8968 1452 8974
rect 1398 8936 1400 8945
rect 1452 8936 1454 8945
rect 1398 8871 1454 8880
rect 1780 8498 1808 9318
rect 1768 8492 1820 8498
rect 1768 8434 1820 8440
rect 1400 6112 1452 6118
rect 1400 6054 1452 6060
rect 1952 6112 2004 6118
rect 1952 6054 2004 6060
rect 1412 5778 1440 6054
rect 1400 5772 1452 5778
rect 1400 5714 1452 5720
rect 1860 5772 1912 5778
rect 1860 5714 1912 5720
rect 1584 5636 1636 5642
rect 1584 5578 1636 5584
rect 1596 4826 1624 5578
rect 1872 5545 1900 5714
rect 1858 5536 1914 5545
rect 1858 5471 1914 5480
rect 1964 5234 1992 6054
rect 2148 5778 2176 9998
rect 2228 9376 2280 9382
rect 2228 9318 2280 9324
rect 2240 9042 2268 9318
rect 2228 9036 2280 9042
rect 2228 8978 2280 8984
rect 2136 5772 2188 5778
rect 2136 5714 2188 5720
rect 1952 5228 2004 5234
rect 1952 5170 2004 5176
rect 1584 4820 1636 4826
rect 1584 4762 1636 4768
rect 1492 4616 1544 4622
rect 1492 4558 1544 4564
rect 2136 4616 2188 4622
rect 2136 4558 2188 4564
rect 1400 3528 1452 3534
rect 1398 3496 1400 3505
rect 1452 3496 1454 3505
rect 1398 3431 1454 3440
rect 664 3120 716 3126
rect 664 3062 716 3068
rect 676 800 704 3062
rect 1400 3052 1452 3058
rect 1504 3040 1532 4558
rect 1452 3012 1532 3040
rect 1400 2994 1452 3000
rect 1584 2984 1636 2990
rect 1584 2926 1636 2932
rect 1596 2650 1624 2926
rect 1584 2644 1636 2650
rect 1584 2586 1636 2592
rect 2148 2446 2176 4558
rect 2424 4146 2452 38830
rect 2778 38176 2834 38185
rect 2778 38111 2834 38120
rect 2792 37806 2820 38111
rect 2780 37800 2832 37806
rect 2780 37742 2832 37748
rect 2976 37262 3004 41511
rect 3700 41132 3752 41138
rect 3700 41074 3752 41080
rect 3240 40520 3292 40526
rect 3240 40462 3292 40468
rect 3056 40452 3108 40458
rect 3056 40394 3108 40400
rect 3068 40186 3096 40394
rect 3056 40180 3108 40186
rect 3056 40122 3108 40128
rect 3252 39642 3280 40462
rect 3514 40216 3570 40225
rect 3514 40151 3570 40160
rect 3528 40118 3556 40151
rect 3712 40118 3740 41074
rect 3792 41064 3844 41070
rect 3792 41006 3844 41012
rect 4712 41064 4764 41070
rect 4712 41006 4764 41012
rect 3516 40112 3568 40118
rect 3516 40054 3568 40060
rect 3700 40112 3752 40118
rect 3700 40054 3752 40060
rect 3240 39636 3292 39642
rect 3240 39578 3292 39584
rect 3804 38962 3832 41006
rect 4214 40828 4522 40848
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40752 4522 40772
rect 4724 40050 4752 41006
rect 4908 40594 4936 43302
rect 5170 43302 5304 43330
rect 5170 43200 5226 43302
rect 4896 40588 4948 40594
rect 4896 40530 4948 40536
rect 4712 40044 4764 40050
rect 4712 39986 4764 39992
rect 4620 39976 4672 39982
rect 4620 39918 4672 39924
rect 4214 39740 4522 39760
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39664 4522 39684
rect 4632 39574 4660 39918
rect 4988 39908 5040 39914
rect 4988 39850 5040 39856
rect 4620 39568 4672 39574
rect 4620 39510 4672 39516
rect 3792 38956 3844 38962
rect 3792 38898 3844 38904
rect 4214 38652 4522 38672
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38576 4522 38596
rect 4436 38276 4488 38282
rect 4436 38218 4488 38224
rect 4252 38208 4304 38214
rect 4252 38150 4304 38156
rect 4264 37942 4292 38150
rect 4252 37936 4304 37942
rect 4252 37878 4304 37884
rect 4448 37874 4476 38218
rect 4436 37868 4488 37874
rect 4436 37810 4488 37816
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 4632 37346 4660 39510
rect 4804 39364 4856 39370
rect 4804 39306 4856 39312
rect 4816 39098 4844 39306
rect 4804 39092 4856 39098
rect 4804 39034 4856 39040
rect 4712 38956 4764 38962
rect 4712 38898 4764 38904
rect 4540 37318 4660 37346
rect 2964 37256 3016 37262
rect 2964 37198 3016 37204
rect 3606 36816 3662 36825
rect 3606 36751 3662 36760
rect 2870 36136 2926 36145
rect 2870 36071 2926 36080
rect 2780 36032 2832 36038
rect 2780 35974 2832 35980
rect 2792 35766 2820 35974
rect 2780 35760 2832 35766
rect 2780 35702 2832 35708
rect 2884 35630 2912 36071
rect 2872 35624 2924 35630
rect 2872 35566 2924 35572
rect 2778 28656 2834 28665
rect 2778 28591 2780 28600
rect 2832 28591 2834 28600
rect 2780 28562 2832 28568
rect 2596 28076 2648 28082
rect 2596 28018 2648 28024
rect 2608 19718 2636 28018
rect 3620 24274 3648 36751
rect 4540 36718 4568 37318
rect 4620 37256 4672 37262
rect 4620 37198 4672 37204
rect 4632 36786 4660 37198
rect 4620 36780 4672 36786
rect 4620 36722 4672 36728
rect 4528 36712 4580 36718
rect 4528 36654 4580 36660
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 4528 36304 4580 36310
rect 4528 36246 4580 36252
rect 4540 35894 4568 36246
rect 4632 36174 4660 36722
rect 4620 36168 4672 36174
rect 4620 36110 4672 36116
rect 4540 35866 4660 35894
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 3608 24268 3660 24274
rect 3608 24210 3660 24216
rect 3424 24132 3476 24138
rect 3424 24074 3476 24080
rect 3436 23866 3464 24074
rect 3424 23860 3476 23866
rect 3424 23802 3476 23808
rect 3332 23724 3384 23730
rect 3332 23666 3384 23672
rect 2688 21480 2740 21486
rect 2688 21422 2740 21428
rect 2780 21480 2832 21486
rect 2780 21422 2832 21428
rect 2700 21146 2728 21422
rect 2792 21185 2820 21422
rect 2778 21176 2834 21185
rect 2688 21140 2740 21146
rect 2778 21111 2834 21120
rect 2688 21082 2740 21088
rect 3344 20942 3372 23666
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 3332 20936 3384 20942
rect 3332 20878 3384 20884
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 2596 19712 2648 19718
rect 2596 19654 2648 19660
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 2778 17776 2834 17785
rect 2778 17711 2834 17720
rect 2792 17134 2820 17711
rect 2780 17128 2832 17134
rect 2780 17070 2832 17076
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 2778 15056 2834 15065
rect 2778 14991 2834 15000
rect 2792 14958 2820 14991
rect 2780 14952 2832 14958
rect 2780 14894 2832 14900
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 2964 14408 3016 14414
rect 2964 14350 3016 14356
rect 2780 13864 2832 13870
rect 2780 13806 2832 13812
rect 2872 13864 2924 13870
rect 2872 13806 2924 13812
rect 2792 13530 2820 13806
rect 2884 13705 2912 13806
rect 2870 13696 2926 13705
rect 2870 13631 2926 13640
rect 2780 13524 2832 13530
rect 2780 13466 2832 13472
rect 2778 12336 2834 12345
rect 2778 12271 2780 12280
rect 2832 12271 2834 12280
rect 2780 12242 2832 12248
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 2792 10305 2820 10542
rect 2778 10296 2834 10305
rect 2778 10231 2834 10240
rect 2872 9376 2924 9382
rect 2872 9318 2924 9324
rect 2884 8566 2912 9318
rect 2872 8560 2924 8566
rect 2872 8502 2924 8508
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2792 8265 2820 8366
rect 2778 8256 2834 8265
rect 2778 8191 2834 8200
rect 2780 6112 2832 6118
rect 2780 6054 2832 6060
rect 2792 5302 2820 6054
rect 2780 5296 2832 5302
rect 2780 5238 2832 5244
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 2792 4865 2820 5102
rect 2778 4856 2834 4865
rect 2778 4791 2834 4800
rect 2412 4140 2464 4146
rect 2412 4082 2464 4088
rect 2780 2984 2832 2990
rect 2780 2926 2832 2932
rect 2136 2440 2188 2446
rect 2136 2382 2188 2388
rect 2792 1465 2820 2926
rect 2976 2446 3004 14350
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 3240 10056 3292 10062
rect 3240 9998 3292 10004
rect 3252 9042 3280 9998
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 3240 9036 3292 9042
rect 3240 8978 3292 8984
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 4066 6896 4122 6905
rect 4066 6831 4068 6840
rect 4120 6831 4122 6840
rect 4068 6802 4120 6808
rect 4632 6798 4660 35866
rect 4724 9586 4752 38898
rect 4896 37188 4948 37194
rect 4896 37130 4948 37136
rect 4908 36854 4936 37130
rect 4896 36848 4948 36854
rect 4896 36790 4948 36796
rect 4908 36378 4936 36790
rect 5000 36718 5028 39850
rect 5276 39506 5304 43302
rect 5814 43200 5870 44000
rect 6458 43200 6514 44000
rect 7746 43330 7802 44000
rect 7746 43302 7972 43330
rect 7746 43200 7802 43302
rect 7944 41206 7972 43302
rect 8390 43200 8446 44000
rect 9034 43200 9090 44000
rect 9678 43200 9734 44000
rect 10966 43200 11022 44000
rect 11610 43200 11666 44000
rect 12254 43200 12310 44000
rect 12898 43200 12954 44000
rect 14186 43200 14242 44000
rect 14830 43200 14886 44000
rect 15474 43200 15530 44000
rect 16762 43200 16818 44000
rect 17406 43200 17462 44000
rect 18050 43200 18106 44000
rect 18694 43200 18750 44000
rect 19982 43200 20038 44000
rect 20626 43200 20682 44000
rect 21270 43200 21326 44000
rect 21914 43200 21970 44000
rect 23202 43330 23258 44000
rect 23202 43302 23428 43330
rect 23202 43200 23258 43302
rect 5816 41200 5868 41206
rect 5816 41142 5868 41148
rect 7932 41200 7984 41206
rect 7932 41142 7984 41148
rect 5632 40452 5684 40458
rect 5632 40394 5684 40400
rect 5644 40050 5672 40394
rect 5632 40044 5684 40050
rect 5632 39986 5684 39992
rect 5264 39500 5316 39506
rect 5264 39442 5316 39448
rect 5828 36786 5856 41142
rect 8024 40928 8076 40934
rect 8024 40870 8076 40876
rect 7196 40112 7248 40118
rect 7196 40054 7248 40060
rect 6736 40044 6788 40050
rect 6736 39986 6788 39992
rect 6460 39840 6512 39846
rect 6460 39782 6512 39788
rect 6472 39506 6500 39782
rect 6748 39506 6776 39986
rect 6460 39500 6512 39506
rect 6460 39442 6512 39448
rect 6736 39500 6788 39506
rect 6736 39442 6788 39448
rect 5540 36780 5592 36786
rect 5540 36722 5592 36728
rect 5816 36780 5868 36786
rect 5816 36722 5868 36728
rect 4988 36712 5040 36718
rect 4988 36654 5040 36660
rect 4896 36372 4948 36378
rect 4896 36314 4948 36320
rect 5000 36310 5028 36654
rect 5080 36576 5132 36582
rect 5080 36518 5132 36524
rect 4988 36304 5040 36310
rect 4988 36246 5040 36252
rect 5092 36174 5120 36518
rect 5080 36168 5132 36174
rect 5080 36110 5132 36116
rect 5092 35698 5120 36110
rect 5172 36100 5224 36106
rect 5172 36042 5224 36048
rect 5080 35692 5132 35698
rect 5080 35634 5132 35640
rect 4804 35624 4856 35630
rect 4804 35566 4856 35572
rect 4816 34746 4844 35566
rect 4804 34740 4856 34746
rect 4804 34682 4856 34688
rect 4712 9580 4764 9586
rect 4712 9522 4764 9528
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 4172 6390 4200 6598
rect 4160 6384 4212 6390
rect 4160 6326 4212 6332
rect 3976 6248 4028 6254
rect 3976 6190 4028 6196
rect 3988 5914 4016 6190
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 3240 4616 3292 4622
rect 3240 4558 3292 4564
rect 3146 4176 3202 4185
rect 3146 4111 3148 4120
rect 3200 4111 3202 4120
rect 3148 4082 3200 4088
rect 3056 3936 3108 3942
rect 3056 3878 3108 3884
rect 3068 3602 3096 3878
rect 3252 3602 3280 4558
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 3056 3596 3108 3602
rect 3056 3538 3108 3544
rect 3240 3596 3292 3602
rect 3240 3538 3292 3544
rect 4252 3528 4304 3534
rect 4252 3470 4304 3476
rect 4264 3194 4292 3470
rect 4252 3188 4304 3194
rect 4252 3130 4304 3136
rect 3240 2916 3292 2922
rect 3240 2858 3292 2864
rect 2964 2440 3016 2446
rect 2964 2382 3016 2388
rect 2778 1456 2834 1465
rect 2778 1391 2834 1400
rect 3252 800 3280 2858
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 3436 2145 3464 2586
rect 4632 2582 4660 4966
rect 4816 4758 4844 34682
rect 5080 6248 5132 6254
rect 5080 6190 5132 6196
rect 4988 5704 5040 5710
rect 4988 5646 5040 5652
rect 4804 4752 4856 4758
rect 4804 4694 4856 4700
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 4724 3602 4752 4558
rect 4804 4480 4856 4486
rect 4804 4422 4856 4428
rect 4816 4078 4844 4422
rect 5000 4146 5028 5646
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 4804 4072 4856 4078
rect 4804 4014 4856 4020
rect 4896 3936 4948 3942
rect 4896 3878 4948 3884
rect 4908 3602 4936 3878
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 4896 3596 4948 3602
rect 4896 3538 4948 3544
rect 4620 2576 4672 2582
rect 4620 2518 4672 2524
rect 3976 2508 4028 2514
rect 3976 2450 4028 2456
rect 3422 2136 3478 2145
rect 3422 2071 3478 2080
rect 3988 1170 4016 2450
rect 3896 1142 4016 1170
rect 3896 800 3924 1142
rect 4540 870 4660 898
rect 4540 800 4568 870
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 1950 0 2006 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 4632 762 4660 870
rect 5092 762 5120 6190
rect 5184 4554 5212 36042
rect 5448 20868 5500 20874
rect 5448 20810 5500 20816
rect 5460 20058 5488 20810
rect 5552 20466 5580 36722
rect 5630 24304 5686 24313
rect 5630 24239 5632 24248
rect 5684 24239 5686 24248
rect 5632 24210 5684 24216
rect 6368 21548 6420 21554
rect 6368 21490 6420 21496
rect 6380 20942 6408 21490
rect 5724 20936 5776 20942
rect 5724 20878 5776 20884
rect 6368 20936 6420 20942
rect 6368 20878 6420 20884
rect 5736 20602 5764 20878
rect 5724 20596 5776 20602
rect 5724 20538 5776 20544
rect 6380 20466 6408 20878
rect 5540 20460 5592 20466
rect 5540 20402 5592 20408
rect 6368 20460 6420 20466
rect 6368 20402 6420 20408
rect 5448 20052 5500 20058
rect 5448 19994 5500 20000
rect 6380 19854 6408 20402
rect 6748 19922 6776 39442
rect 7208 26234 7236 40054
rect 7472 36032 7524 36038
rect 7472 35974 7524 35980
rect 7116 26206 7236 26234
rect 7116 21486 7144 26206
rect 7104 21480 7156 21486
rect 7104 21422 7156 21428
rect 6736 19916 6788 19922
rect 6736 19858 6788 19864
rect 6368 19848 6420 19854
rect 6368 19790 6420 19796
rect 6748 16574 6776 19858
rect 6748 16546 6868 16574
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 5172 4548 5224 4554
rect 5172 4490 5224 4496
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 5184 800 5212 3538
rect 5356 3392 5408 3398
rect 5356 3334 5408 3340
rect 5368 3126 5396 3334
rect 5356 3120 5408 3126
rect 5356 3062 5408 3068
rect 5552 3058 5580 4626
rect 6368 3936 6420 3942
rect 6368 3878 6420 3884
rect 5540 3052 5592 3058
rect 5540 2994 5592 3000
rect 6380 2514 6408 3878
rect 6552 2848 6604 2854
rect 6552 2790 6604 2796
rect 6564 2514 6592 2790
rect 6840 2582 6868 16546
rect 7116 16114 7144 21422
rect 7484 21146 7512 35974
rect 8036 29850 8064 40870
rect 9128 40520 9180 40526
rect 9128 40462 9180 40468
rect 8208 40112 8260 40118
rect 8208 40054 8260 40060
rect 8220 39545 8248 40054
rect 9140 40050 9168 40462
rect 9128 40044 9180 40050
rect 9128 39986 9180 39992
rect 9692 39982 9720 43200
rect 10968 40928 11020 40934
rect 10968 40870 11020 40876
rect 10980 40594 11008 40870
rect 11624 40594 11652 43200
rect 10968 40588 11020 40594
rect 10968 40530 11020 40536
rect 11612 40588 11664 40594
rect 11612 40530 11664 40536
rect 12268 39982 12296 43200
rect 12912 41070 12940 43200
rect 14200 41414 14228 43200
rect 20640 41414 20668 43200
rect 14200 41386 14320 41414
rect 12900 41064 12952 41070
rect 12900 41006 12952 41012
rect 12992 41064 13044 41070
rect 12992 41006 13044 41012
rect 13544 41064 13596 41070
rect 13544 41006 13596 41012
rect 9312 39976 9364 39982
rect 9312 39918 9364 39924
rect 9680 39976 9732 39982
rect 9680 39918 9732 39924
rect 12256 39976 12308 39982
rect 12256 39918 12308 39924
rect 9324 39642 9352 39918
rect 12440 39908 12492 39914
rect 12440 39850 12492 39856
rect 9312 39636 9364 39642
rect 9312 39578 9364 39584
rect 8206 39536 8262 39545
rect 8206 39471 8262 39480
rect 12452 39438 12480 39850
rect 13004 39642 13032 41006
rect 13360 40656 13412 40662
rect 13360 40598 13412 40604
rect 13176 40520 13228 40526
rect 13176 40462 13228 40468
rect 13188 40390 13216 40462
rect 13176 40384 13228 40390
rect 13176 40326 13228 40332
rect 12992 39636 13044 39642
rect 12992 39578 13044 39584
rect 9220 39432 9272 39438
rect 9220 39374 9272 39380
rect 10232 39432 10284 39438
rect 10232 39374 10284 39380
rect 10876 39432 10928 39438
rect 10876 39374 10928 39380
rect 12440 39432 12492 39438
rect 12440 39374 12492 39380
rect 13084 39432 13136 39438
rect 13084 39374 13136 39380
rect 8944 39364 8996 39370
rect 8944 39306 8996 39312
rect 8852 38956 8904 38962
rect 8852 38898 8904 38904
rect 8864 38350 8892 38898
rect 8956 38894 8984 39306
rect 8944 38888 8996 38894
rect 8944 38830 8996 38836
rect 9232 38758 9260 39374
rect 9586 38992 9642 39001
rect 9586 38927 9588 38936
rect 9640 38927 9642 38936
rect 9588 38898 9640 38904
rect 9220 38752 9272 38758
rect 9220 38694 9272 38700
rect 8852 38344 8904 38350
rect 8852 38286 8904 38292
rect 8864 35894 8892 38286
rect 8864 35866 8984 35894
rect 8024 29844 8076 29850
rect 8024 29786 8076 29792
rect 7472 21140 7524 21146
rect 7472 21082 7524 21088
rect 8116 21140 8168 21146
rect 8116 21082 8168 21088
rect 8128 20466 8156 21082
rect 8116 20460 8168 20466
rect 8116 20402 8168 20408
rect 7656 20392 7708 20398
rect 7656 20334 7708 20340
rect 7668 16794 7696 20334
rect 7656 16788 7708 16794
rect 7656 16730 7708 16736
rect 7104 16108 7156 16114
rect 7104 16050 7156 16056
rect 7116 15366 7144 16050
rect 7104 15360 7156 15366
rect 7104 15302 7156 15308
rect 7564 15360 7616 15366
rect 7564 15302 7616 15308
rect 7576 4078 7604 15302
rect 7668 6458 7696 16730
rect 7656 6452 7708 6458
rect 7656 6394 7708 6400
rect 7564 4072 7616 4078
rect 7564 4014 7616 4020
rect 8128 3738 8156 20402
rect 8956 19514 8984 35866
rect 9232 22642 9260 38694
rect 9220 22636 9272 22642
rect 9220 22578 9272 22584
rect 8944 19508 8996 19514
rect 8944 19450 8996 19456
rect 9404 13320 9456 13326
rect 9404 13262 9456 13268
rect 9416 12442 9444 13262
rect 9404 12436 9456 12442
rect 9404 12378 9456 12384
rect 9416 11762 9444 12378
rect 9404 11756 9456 11762
rect 9404 11698 9456 11704
rect 9220 11552 9272 11558
rect 9220 11494 9272 11500
rect 8116 3732 8168 3738
rect 8116 3674 8168 3680
rect 9232 3602 9260 11494
rect 9220 3596 9272 3602
rect 9220 3538 9272 3544
rect 7196 3528 7248 3534
rect 7196 3470 7248 3476
rect 7208 3058 7236 3470
rect 7380 3392 7432 3398
rect 7380 3334 7432 3340
rect 7392 3126 7420 3334
rect 9600 3194 9628 38898
rect 10244 36786 10272 39374
rect 10416 39296 10468 39302
rect 10416 39238 10468 39244
rect 10428 38962 10456 39238
rect 10888 38962 10916 39374
rect 10416 38956 10468 38962
rect 10416 38898 10468 38904
rect 10876 38956 10928 38962
rect 10876 38898 10928 38904
rect 10324 38888 10376 38894
rect 10324 38830 10376 38836
rect 10232 36780 10284 36786
rect 10232 36722 10284 36728
rect 10336 31210 10364 38830
rect 10888 38350 10916 38898
rect 12348 38888 12400 38894
rect 12346 38856 12348 38865
rect 12400 38856 12402 38865
rect 12346 38791 12402 38800
rect 11980 38752 12032 38758
rect 11980 38694 12032 38700
rect 10876 38344 10928 38350
rect 10876 38286 10928 38292
rect 10888 37874 10916 38286
rect 11428 38208 11480 38214
rect 11428 38150 11480 38156
rect 10876 37868 10928 37874
rect 10876 37810 10928 37816
rect 10324 31204 10376 31210
rect 10324 31146 10376 31152
rect 10324 20528 10376 20534
rect 10324 20470 10376 20476
rect 10336 19854 10364 20470
rect 10324 19848 10376 19854
rect 10324 19790 10376 19796
rect 11244 19848 11296 19854
rect 11244 19790 11296 19796
rect 11256 19378 11284 19790
rect 10692 19372 10744 19378
rect 10692 19314 10744 19320
rect 11244 19372 11296 19378
rect 11244 19314 11296 19320
rect 10704 13326 10732 19314
rect 11256 18766 11284 19314
rect 11244 18760 11296 18766
rect 11244 18702 11296 18708
rect 11256 17678 11284 18702
rect 11152 17672 11204 17678
rect 11152 17614 11204 17620
rect 11244 17672 11296 17678
rect 11244 17614 11296 17620
rect 11164 15366 11192 17614
rect 11152 15360 11204 15366
rect 11152 15302 11204 15308
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 11244 4548 11296 4554
rect 11244 4490 11296 4496
rect 10140 4208 10192 4214
rect 10140 4150 10192 4156
rect 10152 4078 10180 4150
rect 10140 4072 10192 4078
rect 10140 4014 10192 4020
rect 10232 4072 10284 4078
rect 10232 4014 10284 4020
rect 9864 3936 9916 3942
rect 9864 3878 9916 3884
rect 9876 3670 9904 3878
rect 9864 3664 9916 3670
rect 9864 3606 9916 3612
rect 9680 3596 9732 3602
rect 9680 3538 9732 3544
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 7380 3120 7432 3126
rect 7380 3062 7432 3068
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 7104 2984 7156 2990
rect 7104 2926 7156 2932
rect 6828 2576 6880 2582
rect 6828 2518 6880 2524
rect 6368 2508 6420 2514
rect 6368 2450 6420 2456
rect 6552 2508 6604 2514
rect 6552 2450 6604 2456
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 6472 870 6592 898
rect 6472 800 6500 870
rect 4632 734 5120 762
rect 5170 0 5226 800
rect 6458 0 6514 800
rect 6564 762 6592 870
rect 6748 762 6776 2450
rect 7116 800 7144 2926
rect 9128 2916 9180 2922
rect 9128 2858 9180 2864
rect 9140 2514 9168 2858
rect 9128 2508 9180 2514
rect 9128 2450 9180 2456
rect 9692 800 9720 3538
rect 10244 3058 10272 4014
rect 10692 4004 10744 4010
rect 10692 3946 10744 3952
rect 10232 3052 10284 3058
rect 10232 2994 10284 3000
rect 10244 2106 10272 2994
rect 10704 2378 10732 3946
rect 10968 2916 11020 2922
rect 10968 2858 11020 2864
rect 10784 2848 10836 2854
rect 10784 2790 10836 2796
rect 10796 2514 10824 2790
rect 10784 2508 10836 2514
rect 10784 2450 10836 2456
rect 10692 2372 10744 2378
rect 10692 2314 10744 2320
rect 10232 2100 10284 2106
rect 10232 2042 10284 2048
rect 10980 800 11008 2858
rect 11256 2774 11284 4490
rect 11440 4078 11468 38150
rect 11992 37942 12020 38694
rect 11980 37936 12032 37942
rect 11980 37878 12032 37884
rect 11980 30116 12032 30122
rect 11980 30058 12032 30064
rect 11992 29578 12020 30058
rect 11980 29572 12032 29578
rect 11980 29514 12032 29520
rect 12072 29572 12124 29578
rect 12072 29514 12124 29520
rect 12084 29170 12112 29514
rect 12072 29164 12124 29170
rect 12072 29106 12124 29112
rect 11888 27532 11940 27538
rect 12084 27520 12112 29106
rect 11940 27492 12112 27520
rect 11888 27474 11940 27480
rect 12084 26450 12112 27492
rect 12072 26444 12124 26450
rect 12072 26386 12124 26392
rect 11612 19916 11664 19922
rect 11612 19858 11664 19864
rect 11624 19718 11652 19858
rect 11612 19712 11664 19718
rect 11612 19654 11664 19660
rect 11520 18216 11572 18222
rect 11520 18158 11572 18164
rect 11532 17202 11560 18158
rect 11520 17196 11572 17202
rect 11520 17138 11572 17144
rect 11624 14414 11652 19654
rect 12164 19440 12216 19446
rect 12164 19382 12216 19388
rect 11704 18692 11756 18698
rect 11704 18634 11756 18640
rect 11612 14408 11664 14414
rect 11612 14350 11664 14356
rect 11716 12889 11744 18634
rect 12072 15360 12124 15366
rect 12072 15302 12124 15308
rect 11796 14272 11848 14278
rect 11796 14214 11848 14220
rect 11808 13938 11836 14214
rect 11796 13932 11848 13938
rect 11796 13874 11848 13880
rect 11980 13864 12032 13870
rect 11980 13806 12032 13812
rect 11992 13530 12020 13806
rect 11980 13524 12032 13530
rect 11980 13466 12032 13472
rect 11702 12880 11758 12889
rect 11702 12815 11758 12824
rect 11716 12442 11744 12815
rect 11704 12436 11756 12442
rect 11704 12378 11756 12384
rect 11428 4072 11480 4078
rect 11428 4014 11480 4020
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 11520 3936 11572 3942
rect 11520 3878 11572 3884
rect 11348 3602 11376 3878
rect 11336 3596 11388 3602
rect 11336 3538 11388 3544
rect 11532 3058 11560 3878
rect 11704 3596 11756 3602
rect 11704 3538 11756 3544
rect 11612 3460 11664 3466
rect 11612 3402 11664 3408
rect 11520 3052 11572 3058
rect 11520 2994 11572 3000
rect 11256 2746 11468 2774
rect 11440 2446 11468 2746
rect 11624 2650 11652 3402
rect 11612 2644 11664 2650
rect 11612 2586 11664 2592
rect 11428 2440 11480 2446
rect 11428 2382 11480 2388
rect 11716 1714 11744 3538
rect 12084 3194 12112 15302
rect 12176 3398 12204 19382
rect 12360 16574 12388 38791
rect 13096 36106 13124 39374
rect 13084 36100 13136 36106
rect 13084 36042 13136 36048
rect 13188 31754 13216 40326
rect 13268 39976 13320 39982
rect 13372 39964 13400 40598
rect 13452 40384 13504 40390
rect 13452 40326 13504 40332
rect 13464 40118 13492 40326
rect 13452 40112 13504 40118
rect 13452 40054 13504 40060
rect 13452 39976 13504 39982
rect 13372 39936 13452 39964
rect 13268 39918 13320 39924
rect 13452 39918 13504 39924
rect 13280 39642 13308 39918
rect 13268 39636 13320 39642
rect 13268 39578 13320 39584
rect 13556 38962 13584 41006
rect 14096 40928 14148 40934
rect 14096 40870 14148 40876
rect 14108 40594 14136 40870
rect 14292 40594 14320 41386
rect 19574 41372 19882 41392
rect 20640 41386 20760 41414
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41296 19882 41316
rect 14740 40928 14792 40934
rect 14740 40870 14792 40876
rect 20168 40928 20220 40934
rect 20168 40870 20220 40876
rect 14096 40588 14148 40594
rect 14096 40530 14148 40536
rect 14280 40588 14332 40594
rect 14280 40530 14332 40536
rect 14280 40452 14332 40458
rect 14280 40394 14332 40400
rect 14292 39642 14320 40394
rect 14752 39982 14780 40870
rect 20180 40594 20208 40870
rect 20732 40594 20760 41386
rect 21824 41064 21876 41070
rect 21824 41006 21876 41012
rect 21836 40730 21864 41006
rect 21928 41002 21956 43200
rect 23400 41414 23428 43302
rect 23846 43200 23902 44000
rect 24490 43200 24546 44000
rect 25134 43200 25190 44000
rect 26422 43200 26478 44000
rect 27066 43330 27122 44000
rect 27066 43302 27384 43330
rect 27066 43200 27122 43302
rect 23400 41386 23520 41414
rect 22008 41064 22060 41070
rect 22008 41006 22060 41012
rect 21916 40996 21968 41002
rect 21916 40938 21968 40944
rect 21824 40724 21876 40730
rect 21824 40666 21876 40672
rect 20168 40588 20220 40594
rect 20168 40530 20220 40536
rect 20720 40588 20772 40594
rect 20720 40530 20772 40536
rect 20352 40452 20404 40458
rect 20352 40394 20404 40400
rect 19574 40284 19882 40304
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40208 19882 40228
rect 20364 40186 20392 40394
rect 22020 40186 22048 41006
rect 23492 40594 23520 41386
rect 23480 40588 23532 40594
rect 23480 40530 23532 40536
rect 20352 40180 20404 40186
rect 20352 40122 20404 40128
rect 22008 40180 22060 40186
rect 22008 40122 22060 40128
rect 20260 40044 20312 40050
rect 20260 39986 20312 39992
rect 21640 40044 21692 40050
rect 21640 39986 21692 39992
rect 14740 39976 14792 39982
rect 14740 39918 14792 39924
rect 15936 39976 15988 39982
rect 15936 39918 15988 39924
rect 14280 39636 14332 39642
rect 14280 39578 14332 39584
rect 15948 39574 15976 39918
rect 20272 39914 20300 39986
rect 20260 39908 20312 39914
rect 20260 39850 20312 39856
rect 14096 39568 14148 39574
rect 14096 39510 14148 39516
rect 15936 39568 15988 39574
rect 15936 39510 15988 39516
rect 14108 39438 14136 39510
rect 14096 39432 14148 39438
rect 14096 39374 14148 39380
rect 14108 39030 14136 39374
rect 19574 39196 19882 39216
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39120 19882 39140
rect 14096 39024 14148 39030
rect 14096 38966 14148 38972
rect 13544 38956 13596 38962
rect 13544 38898 13596 38904
rect 20272 38418 20300 39850
rect 21652 39302 21680 39986
rect 23860 39982 23888 43200
rect 24504 41206 24532 43200
rect 24492 41200 24544 41206
rect 24492 41142 24544 41148
rect 24952 40928 25004 40934
rect 24952 40870 25004 40876
rect 24584 40452 24636 40458
rect 24584 40394 24636 40400
rect 23296 39976 23348 39982
rect 23296 39918 23348 39924
rect 23480 39976 23532 39982
rect 23480 39918 23532 39924
rect 23848 39976 23900 39982
rect 23848 39918 23900 39924
rect 23308 39642 23336 39918
rect 23296 39636 23348 39642
rect 23296 39578 23348 39584
rect 22744 39432 22796 39438
rect 22744 39374 22796 39380
rect 21640 39296 21692 39302
rect 21640 39238 21692 39244
rect 20260 38412 20312 38418
rect 20260 38354 20312 38360
rect 19574 38108 19882 38128
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38032 19882 38052
rect 17500 37868 17552 37874
rect 17500 37810 17552 37816
rect 16580 37800 16632 37806
rect 16580 37742 16632 37748
rect 16592 37262 16620 37742
rect 17512 37466 17540 37810
rect 17868 37664 17920 37670
rect 17868 37606 17920 37612
rect 18328 37664 18380 37670
rect 18328 37606 18380 37612
rect 17500 37460 17552 37466
rect 17500 37402 17552 37408
rect 17880 37330 17908 37606
rect 17868 37324 17920 37330
rect 17868 37266 17920 37272
rect 14096 37256 14148 37262
rect 14096 37198 14148 37204
rect 16580 37256 16632 37262
rect 16580 37198 16632 37204
rect 17224 37256 17276 37262
rect 17224 37198 17276 37204
rect 14108 36174 14136 37198
rect 15568 37188 15620 37194
rect 15568 37130 15620 37136
rect 15580 36922 15608 37130
rect 16856 37120 16908 37126
rect 16856 37062 16908 37068
rect 15568 36916 15620 36922
rect 15568 36858 15620 36864
rect 14556 36848 14608 36854
rect 14556 36790 14608 36796
rect 14280 36780 14332 36786
rect 14280 36722 14332 36728
rect 14096 36168 14148 36174
rect 14096 36110 14148 36116
rect 14108 33998 14136 36110
rect 14292 35834 14320 36722
rect 14568 36718 14596 36790
rect 15660 36780 15712 36786
rect 15660 36722 15712 36728
rect 15936 36780 15988 36786
rect 15936 36722 15988 36728
rect 14556 36712 14608 36718
rect 14556 36654 14608 36660
rect 14372 36576 14424 36582
rect 14372 36518 14424 36524
rect 14384 36174 14412 36518
rect 14462 36408 14518 36417
rect 14462 36343 14464 36352
rect 14516 36343 14518 36352
rect 14464 36314 14516 36320
rect 14372 36168 14424 36174
rect 14372 36110 14424 36116
rect 14280 35828 14332 35834
rect 14280 35770 14332 35776
rect 14372 34400 14424 34406
rect 14372 34342 14424 34348
rect 14384 33998 14412 34342
rect 14096 33992 14148 33998
rect 14096 33934 14148 33940
rect 14372 33992 14424 33998
rect 14372 33934 14424 33940
rect 14108 32434 14136 33934
rect 14096 32428 14148 32434
rect 14096 32370 14148 32376
rect 14108 31890 14136 32370
rect 14096 31884 14148 31890
rect 14096 31826 14148 31832
rect 13188 31726 13400 31754
rect 13084 29504 13136 29510
rect 13084 29446 13136 29452
rect 13096 29170 13124 29446
rect 13084 29164 13136 29170
rect 13084 29106 13136 29112
rect 12716 28076 12768 28082
rect 12716 28018 12768 28024
rect 12532 27872 12584 27878
rect 12532 27814 12584 27820
rect 12544 27470 12572 27814
rect 12532 27464 12584 27470
rect 12532 27406 12584 27412
rect 12728 27130 12756 28018
rect 13268 27328 13320 27334
rect 13268 27270 13320 27276
rect 12716 27124 12768 27130
rect 12716 27066 12768 27072
rect 13280 26926 13308 27270
rect 13268 26920 13320 26926
rect 13268 26862 13320 26868
rect 12900 26376 12952 26382
rect 12900 26318 12952 26324
rect 12912 24818 12940 26318
rect 12900 24812 12952 24818
rect 12900 24754 12952 24760
rect 12900 22024 12952 22030
rect 12900 21966 12952 21972
rect 12912 20398 12940 21966
rect 12900 20392 12952 20398
rect 12900 20334 12952 20340
rect 12912 19378 12940 20334
rect 13372 19922 13400 31726
rect 14372 31748 14424 31754
rect 14372 31690 14424 31696
rect 14384 31482 14412 31690
rect 14372 31476 14424 31482
rect 14372 31418 14424 31424
rect 14372 31272 14424 31278
rect 14372 31214 14424 31220
rect 14384 30734 14412 31214
rect 14372 30728 14424 30734
rect 14372 30670 14424 30676
rect 13728 30660 13780 30666
rect 13728 30602 13780 30608
rect 13740 30190 13768 30602
rect 14188 30592 14240 30598
rect 14188 30534 14240 30540
rect 14004 30388 14056 30394
rect 14004 30330 14056 30336
rect 14016 30258 14044 30330
rect 14200 30258 14228 30534
rect 14384 30394 14412 30670
rect 14372 30388 14424 30394
rect 14372 30330 14424 30336
rect 14004 30252 14056 30258
rect 14004 30194 14056 30200
rect 14188 30252 14240 30258
rect 14188 30194 14240 30200
rect 13728 30184 13780 30190
rect 13728 30126 13780 30132
rect 14016 29102 14044 30194
rect 14280 29640 14332 29646
rect 14280 29582 14332 29588
rect 14096 29504 14148 29510
rect 14096 29446 14148 29452
rect 14108 29238 14136 29446
rect 14096 29232 14148 29238
rect 14096 29174 14148 29180
rect 14004 29096 14056 29102
rect 14004 29038 14056 29044
rect 13452 28960 13504 28966
rect 13452 28902 13504 28908
rect 13464 28626 13492 28902
rect 13452 28620 13504 28626
rect 13452 28562 13504 28568
rect 14016 28558 14044 29038
rect 14004 28552 14056 28558
rect 14004 28494 14056 28500
rect 14016 28150 14044 28494
rect 14292 28422 14320 29582
rect 14384 28626 14412 30330
rect 14568 30258 14596 36654
rect 15672 36174 15700 36722
rect 15752 36576 15804 36582
rect 15752 36518 15804 36524
rect 15660 36168 15712 36174
rect 15660 36110 15712 36116
rect 15476 36032 15528 36038
rect 15476 35974 15528 35980
rect 15488 35766 15516 35974
rect 15476 35760 15528 35766
rect 15476 35702 15528 35708
rect 15292 35692 15344 35698
rect 15292 35634 15344 35640
rect 15304 35562 15332 35634
rect 15292 35556 15344 35562
rect 15292 35498 15344 35504
rect 14740 35488 14792 35494
rect 14740 35430 14792 35436
rect 14648 34604 14700 34610
rect 14648 34546 14700 34552
rect 14464 30252 14516 30258
rect 14464 30194 14516 30200
rect 14556 30252 14608 30258
rect 14556 30194 14608 30200
rect 14476 30054 14504 30194
rect 14464 30048 14516 30054
rect 14464 29990 14516 29996
rect 14476 29714 14504 29990
rect 14660 29730 14688 34546
rect 14752 34406 14780 35430
rect 15304 34542 15332 35498
rect 15764 35290 15792 36518
rect 15948 36378 15976 36722
rect 15936 36372 15988 36378
rect 15936 36314 15988 36320
rect 16868 36310 16896 37062
rect 17132 36712 17184 36718
rect 17132 36654 17184 36660
rect 16948 36372 17000 36378
rect 16948 36314 17000 36320
rect 16856 36304 16908 36310
rect 16856 36246 16908 36252
rect 16212 36168 16264 36174
rect 16212 36110 16264 36116
rect 16672 36168 16724 36174
rect 16672 36110 16724 36116
rect 16224 36038 16252 36110
rect 16212 36032 16264 36038
rect 16212 35974 16264 35980
rect 15752 35284 15804 35290
rect 15752 35226 15804 35232
rect 16224 35018 16252 35974
rect 16684 35698 16712 36110
rect 16672 35692 16724 35698
rect 16672 35634 16724 35640
rect 16856 35692 16908 35698
rect 16856 35634 16908 35640
rect 16684 35222 16712 35634
rect 16672 35216 16724 35222
rect 16672 35158 16724 35164
rect 16672 35080 16724 35086
rect 16672 35022 16724 35028
rect 15476 35012 15528 35018
rect 15476 34954 15528 34960
rect 16212 35012 16264 35018
rect 16212 34954 16264 34960
rect 15488 34610 15516 34954
rect 16684 34610 16712 35022
rect 15476 34604 15528 34610
rect 15476 34546 15528 34552
rect 16672 34604 16724 34610
rect 16672 34546 16724 34552
rect 15292 34536 15344 34542
rect 15292 34478 15344 34484
rect 16580 34536 16632 34542
rect 16580 34478 16632 34484
rect 14740 34400 14792 34406
rect 14740 34342 14792 34348
rect 15304 34134 15332 34478
rect 15292 34128 15344 34134
rect 15292 34070 15344 34076
rect 15108 32768 15160 32774
rect 15108 32710 15160 32716
rect 15120 32434 15148 32710
rect 15108 32428 15160 32434
rect 15108 32370 15160 32376
rect 15844 32224 15896 32230
rect 15844 32166 15896 32172
rect 15568 31952 15620 31958
rect 15568 31894 15620 31900
rect 15580 31414 15608 31894
rect 15200 31408 15252 31414
rect 15200 31350 15252 31356
rect 15568 31408 15620 31414
rect 15568 31350 15620 31356
rect 14740 31340 14792 31346
rect 14740 31282 14792 31288
rect 14752 30938 14780 31282
rect 15212 30938 15240 31350
rect 15856 31346 15884 32166
rect 16212 31816 16264 31822
rect 16212 31758 16264 31764
rect 15936 31476 15988 31482
rect 15936 31418 15988 31424
rect 15844 31340 15896 31346
rect 15844 31282 15896 31288
rect 14740 30932 14792 30938
rect 14740 30874 14792 30880
rect 15200 30932 15252 30938
rect 15200 30874 15252 30880
rect 15660 30660 15712 30666
rect 15660 30602 15712 30608
rect 15672 30546 15700 30602
rect 15844 30592 15896 30598
rect 15672 30518 15792 30546
rect 15844 30534 15896 30540
rect 14924 30320 14976 30326
rect 14924 30262 14976 30268
rect 14832 30252 14884 30258
rect 14832 30194 14884 30200
rect 14464 29708 14516 29714
rect 14660 29702 14780 29730
rect 14464 29650 14516 29656
rect 14752 29646 14780 29702
rect 14556 29640 14608 29646
rect 14556 29582 14608 29588
rect 14740 29640 14792 29646
rect 14740 29582 14792 29588
rect 14568 28762 14596 29582
rect 14752 29034 14780 29582
rect 14740 29028 14792 29034
rect 14740 28970 14792 28976
rect 14556 28756 14608 28762
rect 14556 28698 14608 28704
rect 14372 28620 14424 28626
rect 14372 28562 14424 28568
rect 14280 28416 14332 28422
rect 14280 28358 14332 28364
rect 14556 28416 14608 28422
rect 14556 28358 14608 28364
rect 14004 28144 14056 28150
rect 14004 28086 14056 28092
rect 14568 28082 14596 28358
rect 14648 28144 14700 28150
rect 14648 28086 14700 28092
rect 14464 28076 14516 28082
rect 14464 28018 14516 28024
rect 14556 28076 14608 28082
rect 14556 28018 14608 28024
rect 14476 27470 14504 28018
rect 14660 27470 14688 28086
rect 14464 27464 14516 27470
rect 14464 27406 14516 27412
rect 14648 27464 14700 27470
rect 14648 27406 14700 27412
rect 14476 26926 14504 27406
rect 14740 26988 14792 26994
rect 14740 26930 14792 26936
rect 14464 26920 14516 26926
rect 14464 26862 14516 26868
rect 14476 26518 14504 26862
rect 14464 26512 14516 26518
rect 14464 26454 14516 26460
rect 14752 26450 14780 26930
rect 14740 26444 14792 26450
rect 14740 26386 14792 26392
rect 14752 26042 14780 26386
rect 14740 26036 14792 26042
rect 14740 25978 14792 25984
rect 14556 25288 14608 25294
rect 14556 25230 14608 25236
rect 14568 24954 14596 25230
rect 14556 24948 14608 24954
rect 14556 24890 14608 24896
rect 13452 24812 13504 24818
rect 13452 24754 13504 24760
rect 13464 24410 13492 24754
rect 13912 24676 13964 24682
rect 13912 24618 13964 24624
rect 13820 24608 13872 24614
rect 13820 24550 13872 24556
rect 13452 24404 13504 24410
rect 13452 24346 13504 24352
rect 13832 24274 13860 24550
rect 13820 24268 13872 24274
rect 13820 24210 13872 24216
rect 13924 24206 13952 24618
rect 14188 24608 14240 24614
rect 14188 24550 14240 24556
rect 13912 24200 13964 24206
rect 13912 24142 13964 24148
rect 14096 20800 14148 20806
rect 14096 20742 14148 20748
rect 14200 20754 14228 24550
rect 14844 24410 14872 30194
rect 14936 29782 14964 30262
rect 15764 30190 15792 30518
rect 15752 30184 15804 30190
rect 15752 30126 15804 30132
rect 14924 29776 14976 29782
rect 14924 29718 14976 29724
rect 14924 29640 14976 29646
rect 14924 29582 14976 29588
rect 15476 29640 15528 29646
rect 15476 29582 15528 29588
rect 14936 28694 14964 29582
rect 15292 29504 15344 29510
rect 15292 29446 15344 29452
rect 14924 28688 14976 28694
rect 14924 28630 14976 28636
rect 15108 27872 15160 27878
rect 15108 27814 15160 27820
rect 15120 27470 15148 27814
rect 15108 27464 15160 27470
rect 15108 27406 15160 27412
rect 15304 26994 15332 29446
rect 15488 29170 15516 29582
rect 15764 29306 15792 30126
rect 15752 29300 15804 29306
rect 15752 29242 15804 29248
rect 15476 29164 15528 29170
rect 15476 29106 15528 29112
rect 15764 28626 15792 29242
rect 15856 28966 15884 30534
rect 15948 29646 15976 31418
rect 16224 30938 16252 31758
rect 16488 31272 16540 31278
rect 16488 31214 16540 31220
rect 16212 30932 16264 30938
rect 16212 30874 16264 30880
rect 16224 30734 16252 30874
rect 16500 30734 16528 31214
rect 16592 30870 16620 34478
rect 16684 33658 16712 34546
rect 16672 33652 16724 33658
rect 16672 33594 16724 33600
rect 16868 33522 16896 35634
rect 16960 35154 16988 36314
rect 17144 35834 17172 36654
rect 17236 36378 17264 37198
rect 18052 37120 18104 37126
rect 18052 37062 18104 37068
rect 18064 36786 18092 37062
rect 17500 36780 17552 36786
rect 17500 36722 17552 36728
rect 18052 36780 18104 36786
rect 18052 36722 18104 36728
rect 17512 36582 17540 36722
rect 18144 36712 18196 36718
rect 18144 36654 18196 36660
rect 17316 36576 17368 36582
rect 17316 36518 17368 36524
rect 17500 36576 17552 36582
rect 17500 36518 17552 36524
rect 17328 36378 17356 36518
rect 17224 36372 17276 36378
rect 17224 36314 17276 36320
rect 17316 36372 17368 36378
rect 17316 36314 17368 36320
rect 17960 36168 18012 36174
rect 17960 36110 18012 36116
rect 17132 35828 17184 35834
rect 17132 35770 17184 35776
rect 17224 35692 17276 35698
rect 17224 35634 17276 35640
rect 16948 35148 17000 35154
rect 16948 35090 17000 35096
rect 17236 35086 17264 35634
rect 17972 35630 18000 36110
rect 17960 35624 18012 35630
rect 17960 35566 18012 35572
rect 17224 35080 17276 35086
rect 17224 35022 17276 35028
rect 17236 34746 17264 35022
rect 17224 34740 17276 34746
rect 17224 34682 17276 34688
rect 18156 34610 18184 36654
rect 18234 36408 18290 36417
rect 18234 36343 18290 36352
rect 18248 36310 18276 36343
rect 18236 36304 18288 36310
rect 18236 36246 18288 36252
rect 18340 36242 18368 37606
rect 20812 37460 20864 37466
rect 20812 37402 20864 37408
rect 18604 37256 18656 37262
rect 18604 37198 18656 37204
rect 20720 37256 20772 37262
rect 20720 37198 20772 37204
rect 18616 36922 18644 37198
rect 20536 37188 20588 37194
rect 20536 37130 20588 37136
rect 19248 37120 19300 37126
rect 19248 37062 19300 37068
rect 18604 36916 18656 36922
rect 18604 36858 18656 36864
rect 19260 36718 19288 37062
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 20548 36922 20576 37130
rect 20536 36916 20588 36922
rect 20536 36858 20588 36864
rect 20352 36780 20404 36786
rect 20404 36740 20484 36768
rect 20352 36722 20404 36728
rect 19248 36712 19300 36718
rect 19248 36654 19300 36660
rect 18512 36576 18564 36582
rect 18512 36518 18564 36524
rect 18328 36236 18380 36242
rect 18380 36196 18460 36224
rect 18328 36178 18380 36184
rect 18328 35488 18380 35494
rect 18328 35430 18380 35436
rect 18236 35148 18288 35154
rect 18236 35090 18288 35096
rect 18248 34610 18276 35090
rect 18340 35000 18368 35430
rect 18432 35154 18460 36196
rect 18524 36106 18552 36518
rect 19248 36168 19300 36174
rect 19248 36110 19300 36116
rect 18512 36100 18564 36106
rect 18512 36042 18564 36048
rect 19064 35488 19116 35494
rect 19064 35430 19116 35436
rect 18420 35148 18472 35154
rect 18420 35090 18472 35096
rect 18420 35012 18472 35018
rect 18340 34972 18420 35000
rect 18144 34604 18196 34610
rect 18144 34546 18196 34552
rect 18236 34604 18288 34610
rect 18236 34546 18288 34552
rect 18156 34474 18184 34546
rect 18144 34468 18196 34474
rect 18144 34410 18196 34416
rect 18156 34134 18184 34410
rect 18144 34128 18196 34134
rect 18144 34070 18196 34076
rect 18340 33998 18368 34972
rect 18420 34954 18472 34960
rect 18972 34672 19024 34678
rect 18972 34614 19024 34620
rect 18420 34604 18472 34610
rect 18420 34546 18472 34552
rect 18512 34604 18564 34610
rect 18512 34546 18564 34552
rect 18328 33992 18380 33998
rect 18328 33934 18380 33940
rect 18236 33924 18288 33930
rect 18236 33866 18288 33872
rect 16856 33516 16908 33522
rect 16856 33458 16908 33464
rect 17408 33380 17460 33386
rect 17408 33322 17460 33328
rect 16856 32904 16908 32910
rect 16856 32846 16908 32852
rect 16868 32026 16896 32846
rect 16856 32020 16908 32026
rect 16856 31962 16908 31968
rect 17420 31822 17448 33322
rect 17960 33312 18012 33318
rect 17960 33254 18012 33260
rect 17972 32910 18000 33254
rect 18248 32910 18276 33866
rect 18432 32978 18460 34546
rect 18524 34202 18552 34546
rect 18984 34202 19012 34614
rect 18512 34196 18564 34202
rect 18512 34138 18564 34144
rect 18972 34196 19024 34202
rect 18972 34138 19024 34144
rect 18696 33992 18748 33998
rect 18696 33934 18748 33940
rect 18420 32972 18472 32978
rect 18420 32914 18472 32920
rect 17960 32904 18012 32910
rect 17960 32846 18012 32852
rect 18236 32904 18288 32910
rect 18236 32846 18288 32852
rect 18512 32904 18564 32910
rect 18512 32846 18564 32852
rect 18328 32836 18380 32842
rect 18328 32778 18380 32784
rect 18236 32428 18288 32434
rect 18236 32370 18288 32376
rect 18248 32026 18276 32370
rect 18340 32366 18368 32778
rect 18420 32768 18472 32774
rect 18420 32710 18472 32716
rect 18328 32360 18380 32366
rect 18328 32302 18380 32308
rect 18236 32020 18288 32026
rect 18236 31962 18288 31968
rect 18432 31822 18460 32710
rect 18524 32230 18552 32846
rect 18708 32774 18736 33934
rect 18788 33924 18840 33930
rect 18788 33866 18840 33872
rect 18800 32910 18828 33866
rect 19076 33658 19104 35430
rect 19260 34592 19288 36110
rect 19432 36032 19484 36038
rect 19432 35974 19484 35980
rect 19444 35714 19472 35974
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 19444 35686 19564 35714
rect 19536 35170 19564 35686
rect 19616 35692 19668 35698
rect 19616 35634 19668 35640
rect 19628 35290 19656 35634
rect 20168 35556 20220 35562
rect 20168 35498 20220 35504
rect 19616 35284 19668 35290
rect 19616 35226 19668 35232
rect 19536 35142 19748 35170
rect 19720 35086 19748 35142
rect 19984 35148 20036 35154
rect 19984 35090 20036 35096
rect 19708 35080 19760 35086
rect 19708 35022 19760 35028
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 19432 34672 19484 34678
rect 19432 34614 19484 34620
rect 19340 34604 19392 34610
rect 19260 34564 19340 34592
rect 19340 34546 19392 34552
rect 19444 33998 19472 34614
rect 19432 33992 19484 33998
rect 19432 33934 19484 33940
rect 19996 33930 20024 35090
rect 20076 35012 20128 35018
rect 20076 34954 20128 34960
rect 20088 34134 20116 34954
rect 20180 34474 20208 35498
rect 20260 34944 20312 34950
rect 20260 34886 20312 34892
rect 20168 34468 20220 34474
rect 20168 34410 20220 34416
rect 20168 34196 20220 34202
rect 20168 34138 20220 34144
rect 20076 34128 20128 34134
rect 20076 34070 20128 34076
rect 20088 33998 20116 34070
rect 20076 33992 20128 33998
rect 20076 33934 20128 33940
rect 19984 33924 20036 33930
rect 19984 33866 20036 33872
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 19064 33652 19116 33658
rect 19064 33594 19116 33600
rect 19156 33584 19208 33590
rect 19156 33526 19208 33532
rect 18880 33516 18932 33522
rect 18880 33458 18932 33464
rect 19064 33516 19116 33522
rect 19064 33458 19116 33464
rect 18892 33114 18920 33458
rect 18880 33108 18932 33114
rect 18880 33050 18932 33056
rect 18788 32904 18840 32910
rect 18788 32846 18840 32852
rect 18696 32768 18748 32774
rect 18696 32710 18748 32716
rect 18800 32570 18828 32846
rect 18788 32564 18840 32570
rect 18788 32506 18840 32512
rect 18892 32502 18920 33050
rect 19076 32842 19104 33458
rect 19168 33386 19196 33526
rect 19996 33454 20024 33866
rect 19984 33448 20036 33454
rect 19984 33390 20036 33396
rect 19156 33380 19208 33386
rect 19156 33322 19208 33328
rect 20180 32978 20208 34138
rect 20272 33046 20300 34886
rect 20260 33040 20312 33046
rect 20260 32982 20312 32988
rect 20168 32972 20220 32978
rect 20168 32914 20220 32920
rect 20076 32904 20128 32910
rect 20076 32846 20128 32852
rect 19064 32836 19116 32842
rect 19064 32778 19116 32784
rect 19076 32570 19104 32778
rect 19984 32768 20036 32774
rect 19984 32710 20036 32716
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 19064 32564 19116 32570
rect 19064 32506 19116 32512
rect 18880 32496 18932 32502
rect 18880 32438 18932 32444
rect 19340 32428 19392 32434
rect 19340 32370 19392 32376
rect 19352 32314 19380 32370
rect 19260 32286 19380 32314
rect 19260 32230 19288 32286
rect 18512 32224 18564 32230
rect 18512 32166 18564 32172
rect 19248 32224 19300 32230
rect 19248 32166 19300 32172
rect 17408 31816 17460 31822
rect 17408 31758 17460 31764
rect 17776 31816 17828 31822
rect 17776 31758 17828 31764
rect 18420 31816 18472 31822
rect 18420 31758 18472 31764
rect 16948 31748 17000 31754
rect 16948 31690 17000 31696
rect 17592 31748 17644 31754
rect 17592 31690 17644 31696
rect 16960 31346 16988 31690
rect 16948 31340 17000 31346
rect 16948 31282 17000 31288
rect 16580 30864 16632 30870
rect 16580 30806 16632 30812
rect 16212 30728 16264 30734
rect 16212 30670 16264 30676
rect 16488 30728 16540 30734
rect 16488 30670 16540 30676
rect 16224 29646 16252 30670
rect 16592 30054 16620 30806
rect 16672 30728 16724 30734
rect 16672 30670 16724 30676
rect 16684 30394 16712 30670
rect 16960 30598 16988 31282
rect 17604 30938 17632 31690
rect 17788 31482 17816 31758
rect 17776 31476 17828 31482
rect 17776 31418 17828 31424
rect 17592 30932 17644 30938
rect 17592 30874 17644 30880
rect 17224 30728 17276 30734
rect 17224 30670 17276 30676
rect 17776 30728 17828 30734
rect 17776 30670 17828 30676
rect 16948 30592 17000 30598
rect 16948 30534 17000 30540
rect 16672 30388 16724 30394
rect 16672 30330 16724 30336
rect 17236 30190 17264 30670
rect 17224 30184 17276 30190
rect 17224 30126 17276 30132
rect 16580 30048 16632 30054
rect 16580 29990 16632 29996
rect 16764 29776 16816 29782
rect 16764 29718 16816 29724
rect 15936 29640 15988 29646
rect 15936 29582 15988 29588
rect 16212 29640 16264 29646
rect 16212 29582 16264 29588
rect 16224 29306 16252 29582
rect 16212 29300 16264 29306
rect 16212 29242 16264 29248
rect 16488 29232 16540 29238
rect 16488 29174 16540 29180
rect 15844 28960 15896 28966
rect 15844 28902 15896 28908
rect 15752 28620 15804 28626
rect 15752 28562 15804 28568
rect 15856 28558 15884 28902
rect 16396 28620 16448 28626
rect 16396 28562 16448 28568
rect 15844 28552 15896 28558
rect 15844 28494 15896 28500
rect 15856 28082 15884 28494
rect 15936 28484 15988 28490
rect 15936 28426 15988 28432
rect 15948 28082 15976 28426
rect 15844 28076 15896 28082
rect 15844 28018 15896 28024
rect 15936 28076 15988 28082
rect 15936 28018 15988 28024
rect 15660 28008 15712 28014
rect 15660 27950 15712 27956
rect 15672 26994 15700 27950
rect 15292 26988 15344 26994
rect 15292 26930 15344 26936
rect 15660 26988 15712 26994
rect 15660 26930 15712 26936
rect 15384 26852 15436 26858
rect 15384 26794 15436 26800
rect 15396 26518 15424 26794
rect 15476 26580 15528 26586
rect 15476 26522 15528 26528
rect 15384 26512 15436 26518
rect 15384 26454 15436 26460
rect 15292 26308 15344 26314
rect 15292 26250 15344 26256
rect 15200 26240 15252 26246
rect 15200 26182 15252 26188
rect 15212 25906 15240 26182
rect 15200 25900 15252 25906
rect 15200 25842 15252 25848
rect 15200 25764 15252 25770
rect 15200 25706 15252 25712
rect 14924 24812 14976 24818
rect 14924 24754 14976 24760
rect 14832 24404 14884 24410
rect 14832 24346 14884 24352
rect 14936 24274 14964 24754
rect 14924 24268 14976 24274
rect 14924 24210 14976 24216
rect 15212 24070 15240 25706
rect 15304 25498 15332 26250
rect 15292 25492 15344 25498
rect 15292 25434 15344 25440
rect 15292 25356 15344 25362
rect 15292 25298 15344 25304
rect 15304 24410 15332 25298
rect 15396 25294 15424 26454
rect 15384 25288 15436 25294
rect 15384 25230 15436 25236
rect 15488 24818 15516 26522
rect 15568 26376 15620 26382
rect 15568 26318 15620 26324
rect 15580 26042 15608 26318
rect 15568 26036 15620 26042
rect 15568 25978 15620 25984
rect 15568 25832 15620 25838
rect 15568 25774 15620 25780
rect 15580 25294 15608 25774
rect 15844 25764 15896 25770
rect 15844 25706 15896 25712
rect 15568 25288 15620 25294
rect 15568 25230 15620 25236
rect 15476 24812 15528 24818
rect 15476 24754 15528 24760
rect 15580 24410 15608 25230
rect 15856 24886 15884 25706
rect 15844 24880 15896 24886
rect 15844 24822 15896 24828
rect 15948 24750 15976 28018
rect 16408 27538 16436 28562
rect 16500 28490 16528 29174
rect 16776 29170 16804 29718
rect 17132 29504 17184 29510
rect 17132 29446 17184 29452
rect 16764 29164 16816 29170
rect 16764 29106 16816 29112
rect 16948 28552 17000 28558
rect 16948 28494 17000 28500
rect 16488 28484 16540 28490
rect 16488 28426 16540 28432
rect 16396 27532 16448 27538
rect 16396 27474 16448 27480
rect 16408 26450 16436 27474
rect 16500 27470 16528 28426
rect 16764 27872 16816 27878
rect 16764 27814 16816 27820
rect 16488 27464 16540 27470
rect 16488 27406 16540 27412
rect 16776 27402 16804 27814
rect 16764 27396 16816 27402
rect 16764 27338 16816 27344
rect 16672 26988 16724 26994
rect 16672 26930 16724 26936
rect 16396 26444 16448 26450
rect 16396 26386 16448 26392
rect 16408 25226 16436 26386
rect 16684 26314 16712 26930
rect 16960 26926 16988 28494
rect 17040 28144 17092 28150
rect 17040 28086 17092 28092
rect 17052 27470 17080 28086
rect 17144 28082 17172 29446
rect 17236 29238 17264 30126
rect 17788 30122 17816 30670
rect 18236 30592 18288 30598
rect 18236 30534 18288 30540
rect 17776 30116 17828 30122
rect 17776 30058 17828 30064
rect 17224 29232 17276 29238
rect 17224 29174 17276 29180
rect 17224 29028 17276 29034
rect 17224 28970 17276 28976
rect 17132 28076 17184 28082
rect 17132 28018 17184 28024
rect 17144 27538 17172 28018
rect 17132 27532 17184 27538
rect 17132 27474 17184 27480
rect 17040 27464 17092 27470
rect 17040 27406 17092 27412
rect 16948 26920 17000 26926
rect 16948 26862 17000 26868
rect 16856 26784 16908 26790
rect 16856 26726 16908 26732
rect 16764 26376 16816 26382
rect 16764 26318 16816 26324
rect 16672 26308 16724 26314
rect 16672 26250 16724 26256
rect 16776 25294 16804 26318
rect 16868 25906 16896 26726
rect 16948 26308 17000 26314
rect 16948 26250 17000 26256
rect 16856 25900 16908 25906
rect 16856 25842 16908 25848
rect 16868 25362 16896 25842
rect 16856 25356 16908 25362
rect 16856 25298 16908 25304
rect 16764 25288 16816 25294
rect 16764 25230 16816 25236
rect 16396 25220 16448 25226
rect 16396 25162 16448 25168
rect 16028 24948 16080 24954
rect 16028 24890 16080 24896
rect 15936 24744 15988 24750
rect 15936 24686 15988 24692
rect 15292 24404 15344 24410
rect 15292 24346 15344 24352
rect 15568 24404 15620 24410
rect 15568 24346 15620 24352
rect 15752 24132 15804 24138
rect 15752 24074 15804 24080
rect 14464 24064 14516 24070
rect 14464 24006 14516 24012
rect 15200 24064 15252 24070
rect 15200 24006 15252 24012
rect 14476 23730 14504 24006
rect 14464 23724 14516 23730
rect 14464 23666 14516 23672
rect 14372 23656 14424 23662
rect 14372 23598 14424 23604
rect 14384 22030 14412 23598
rect 15764 23594 15792 24074
rect 16040 23866 16068 24890
rect 16408 24818 16436 25162
rect 16396 24812 16448 24818
rect 16396 24754 16448 24760
rect 16776 24614 16804 25230
rect 16764 24608 16816 24614
rect 16764 24550 16816 24556
rect 16776 24138 16804 24550
rect 16960 24206 16988 26250
rect 17040 25288 17092 25294
rect 17040 25230 17092 25236
rect 17052 24818 17080 25230
rect 17236 24818 17264 28970
rect 17408 28552 17460 28558
rect 17408 28494 17460 28500
rect 17316 28416 17368 28422
rect 17316 28358 17368 28364
rect 17328 28082 17356 28358
rect 17316 28076 17368 28082
rect 17316 28018 17368 28024
rect 17420 27538 17448 28494
rect 17788 28218 17816 30058
rect 18248 29578 18276 30534
rect 18524 30258 18552 32166
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 19996 31414 20024 32710
rect 20088 32026 20116 32846
rect 20076 32020 20128 32026
rect 20076 31962 20128 31968
rect 20272 31958 20300 32982
rect 20352 32972 20404 32978
rect 20352 32914 20404 32920
rect 20364 32434 20392 32914
rect 20352 32428 20404 32434
rect 20352 32370 20404 32376
rect 20456 32314 20484 36740
rect 20628 34128 20680 34134
rect 20628 34070 20680 34076
rect 20640 33590 20668 34070
rect 20628 33584 20680 33590
rect 20628 33526 20680 33532
rect 20536 33448 20588 33454
rect 20536 33390 20588 33396
rect 20548 33318 20576 33390
rect 20536 33312 20588 33318
rect 20536 33254 20588 33260
rect 20364 32286 20484 32314
rect 20260 31952 20312 31958
rect 20260 31894 20312 31900
rect 20364 31770 20392 32286
rect 20548 31822 20576 33254
rect 20732 32298 20760 37198
rect 20824 36786 20852 37402
rect 21088 36916 21140 36922
rect 21088 36858 21140 36864
rect 20812 36780 20864 36786
rect 20812 36722 20864 36728
rect 21100 36174 21128 36858
rect 21088 36168 21140 36174
rect 21088 36110 21140 36116
rect 20904 34604 20956 34610
rect 20904 34546 20956 34552
rect 20916 33658 20944 34546
rect 21088 34400 21140 34406
rect 21088 34342 21140 34348
rect 21100 33998 21128 34342
rect 21088 33992 21140 33998
rect 21088 33934 21140 33940
rect 20904 33652 20956 33658
rect 20904 33594 20956 33600
rect 21272 33584 21324 33590
rect 21272 33526 21324 33532
rect 20812 33516 20864 33522
rect 20812 33458 20864 33464
rect 20824 33114 20852 33458
rect 20812 33108 20864 33114
rect 20812 33050 20864 33056
rect 20812 32836 20864 32842
rect 20812 32778 20864 32784
rect 20720 32292 20772 32298
rect 20720 32234 20772 32240
rect 20628 31952 20680 31958
rect 20628 31894 20680 31900
rect 20272 31754 20392 31770
rect 20536 31816 20588 31822
rect 20536 31758 20588 31764
rect 20180 31742 20392 31754
rect 20180 31726 20300 31742
rect 19984 31408 20036 31414
rect 19984 31350 20036 31356
rect 19248 30796 19300 30802
rect 19248 30738 19300 30744
rect 18512 30252 18564 30258
rect 18512 30194 18564 30200
rect 18420 30116 18472 30122
rect 18420 30058 18472 30064
rect 18432 29578 18460 30058
rect 18524 30054 18552 30194
rect 18512 30048 18564 30054
rect 18512 29990 18564 29996
rect 18524 29782 18552 29990
rect 18512 29776 18564 29782
rect 18512 29718 18564 29724
rect 19260 29646 19288 30738
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19800 30252 19852 30258
rect 19800 30194 19852 30200
rect 19812 29782 19840 30194
rect 19800 29776 19852 29782
rect 19800 29718 19852 29724
rect 18512 29640 18564 29646
rect 18512 29582 18564 29588
rect 18972 29640 19024 29646
rect 18972 29582 19024 29588
rect 19248 29640 19300 29646
rect 19248 29582 19300 29588
rect 18236 29572 18288 29578
rect 18236 29514 18288 29520
rect 18420 29572 18472 29578
rect 18420 29514 18472 29520
rect 18524 29238 18552 29582
rect 18512 29232 18564 29238
rect 18512 29174 18564 29180
rect 18696 29232 18748 29238
rect 18696 29174 18748 29180
rect 18236 28416 18288 28422
rect 18236 28358 18288 28364
rect 17776 28212 17828 28218
rect 17776 28154 17828 28160
rect 18248 28082 18276 28358
rect 18236 28076 18288 28082
rect 18236 28018 18288 28024
rect 17868 28008 17920 28014
rect 17868 27950 17920 27956
rect 18052 28008 18104 28014
rect 18052 27950 18104 27956
rect 17880 27674 17908 27950
rect 17868 27668 17920 27674
rect 17868 27610 17920 27616
rect 18064 27606 18092 27950
rect 18052 27600 18104 27606
rect 18052 27542 18104 27548
rect 18604 27600 18656 27606
rect 18604 27542 18656 27548
rect 17408 27532 17460 27538
rect 17408 27474 17460 27480
rect 17420 26382 17448 27474
rect 17592 27464 17644 27470
rect 17592 27406 17644 27412
rect 17408 26376 17460 26382
rect 17408 26318 17460 26324
rect 17604 25702 17632 27406
rect 18144 27396 18196 27402
rect 18144 27338 18196 27344
rect 17868 25968 17920 25974
rect 17868 25910 17920 25916
rect 17592 25696 17644 25702
rect 17592 25638 17644 25644
rect 17604 25362 17632 25638
rect 17592 25356 17644 25362
rect 17592 25298 17644 25304
rect 17040 24812 17092 24818
rect 17040 24754 17092 24760
rect 17224 24812 17276 24818
rect 17224 24754 17276 24760
rect 17408 24812 17460 24818
rect 17408 24754 17460 24760
rect 17052 24290 17080 24754
rect 17132 24744 17184 24750
rect 17132 24686 17184 24692
rect 17144 24410 17172 24686
rect 17132 24404 17184 24410
rect 17132 24346 17184 24352
rect 17052 24274 17172 24290
rect 17052 24268 17184 24274
rect 17052 24262 17132 24268
rect 16948 24200 17000 24206
rect 16948 24142 17000 24148
rect 16764 24132 16816 24138
rect 16764 24074 16816 24080
rect 16028 23860 16080 23866
rect 16028 23802 16080 23808
rect 17052 23730 17080 24262
rect 17132 24210 17184 24216
rect 17040 23724 17092 23730
rect 17040 23666 17092 23672
rect 16672 23656 16724 23662
rect 16672 23598 16724 23604
rect 15752 23588 15804 23594
rect 15752 23530 15804 23536
rect 15660 22092 15712 22098
rect 15660 22034 15712 22040
rect 16212 22092 16264 22098
rect 16212 22034 16264 22040
rect 14372 22024 14424 22030
rect 14372 21966 14424 21972
rect 15476 22024 15528 22030
rect 15476 21966 15528 21972
rect 15384 21956 15436 21962
rect 15384 21898 15436 21904
rect 15108 21888 15160 21894
rect 15108 21830 15160 21836
rect 14372 21684 14424 21690
rect 14372 21626 14424 21632
rect 14384 20942 14412 21626
rect 15120 21554 15148 21830
rect 14740 21548 14792 21554
rect 14740 21490 14792 21496
rect 15108 21548 15160 21554
rect 15108 21490 15160 21496
rect 14372 20936 14424 20942
rect 14372 20878 14424 20884
rect 14648 20936 14700 20942
rect 14648 20878 14700 20884
rect 14660 20754 14688 20878
rect 14108 20534 14136 20742
rect 14200 20726 14688 20754
rect 14096 20528 14148 20534
rect 14096 20470 14148 20476
rect 13360 19916 13412 19922
rect 13360 19858 13412 19864
rect 12900 19372 12952 19378
rect 12900 19314 12952 19320
rect 12912 18358 12940 19314
rect 13636 18692 13688 18698
rect 13636 18634 13688 18640
rect 12900 18352 12952 18358
rect 12900 18294 12952 18300
rect 13544 18080 13596 18086
rect 13544 18022 13596 18028
rect 13268 17672 13320 17678
rect 13266 17640 13268 17649
rect 13320 17640 13322 17649
rect 13556 17610 13584 18022
rect 13266 17575 13322 17584
rect 13544 17604 13596 17610
rect 13544 17546 13596 17552
rect 13360 17332 13412 17338
rect 13360 17274 13412 17280
rect 13268 16720 13320 16726
rect 13268 16662 13320 16668
rect 12268 16546 12388 16574
rect 12164 3392 12216 3398
rect 12164 3334 12216 3340
rect 12072 3188 12124 3194
rect 12072 3130 12124 3136
rect 12268 3126 12296 16546
rect 13280 16046 13308 16662
rect 13372 16590 13400 17274
rect 13648 17202 13676 18634
rect 13728 18284 13780 18290
rect 13728 18226 13780 18232
rect 13740 17882 13768 18226
rect 13728 17876 13780 17882
rect 13728 17818 13780 17824
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 13728 17604 13780 17610
rect 13728 17546 13780 17552
rect 13740 17270 13768 17546
rect 14108 17338 14136 17614
rect 14096 17332 14148 17338
rect 14096 17274 14148 17280
rect 13728 17264 13780 17270
rect 13728 17206 13780 17212
rect 13452 17196 13504 17202
rect 13452 17138 13504 17144
rect 13636 17196 13688 17202
rect 13636 17138 13688 17144
rect 13360 16584 13412 16590
rect 13360 16526 13412 16532
rect 13372 16182 13400 16526
rect 13360 16176 13412 16182
rect 13360 16118 13412 16124
rect 13268 16040 13320 16046
rect 13268 15982 13320 15988
rect 13280 15706 13308 15982
rect 13360 15904 13412 15910
rect 13360 15846 13412 15852
rect 13268 15700 13320 15706
rect 13268 15642 13320 15648
rect 13372 15502 13400 15846
rect 13464 15706 13492 17138
rect 13544 16448 13596 16454
rect 13544 16390 13596 16396
rect 13452 15700 13504 15706
rect 13452 15642 13504 15648
rect 13556 15502 13584 16390
rect 13648 15638 13676 17138
rect 13820 16992 13872 16998
rect 13820 16934 13872 16940
rect 13832 16658 13860 16934
rect 13820 16652 13872 16658
rect 13820 16594 13872 16600
rect 13636 15632 13688 15638
rect 13636 15574 13688 15580
rect 14004 15564 14056 15570
rect 14004 15506 14056 15512
rect 13360 15496 13412 15502
rect 13360 15438 13412 15444
rect 13544 15496 13596 15502
rect 13544 15438 13596 15444
rect 13820 15496 13872 15502
rect 13820 15438 13872 15444
rect 14016 15450 14044 15506
rect 13176 15428 13228 15434
rect 13176 15370 13228 15376
rect 13452 15428 13504 15434
rect 13452 15370 13504 15376
rect 13188 15162 13216 15370
rect 13176 15156 13228 15162
rect 13176 15098 13228 15104
rect 13464 15026 13492 15370
rect 13556 15162 13584 15438
rect 13544 15156 13596 15162
rect 13544 15098 13596 15104
rect 13452 15020 13504 15026
rect 13452 14962 13504 14968
rect 13464 14414 13492 14962
rect 13556 14482 13584 15098
rect 13832 14618 13860 15438
rect 14016 15422 14136 15450
rect 14108 14890 14136 15422
rect 14200 15026 14228 20726
rect 14752 20330 14780 21490
rect 14830 20904 14886 20913
rect 14830 20839 14886 20848
rect 15016 20868 15068 20874
rect 14844 20534 14872 20839
rect 15016 20810 15068 20816
rect 14832 20528 14884 20534
rect 14832 20470 14884 20476
rect 14740 20324 14792 20330
rect 14740 20266 14792 20272
rect 15028 19446 15056 20810
rect 15120 20262 15148 21490
rect 15396 21146 15424 21898
rect 15488 21554 15516 21966
rect 15476 21548 15528 21554
rect 15476 21490 15528 21496
rect 15384 21140 15436 21146
rect 15384 21082 15436 21088
rect 15672 20942 15700 22034
rect 15844 22024 15896 22030
rect 15844 21966 15896 21972
rect 15856 21486 15884 21966
rect 16224 21690 16252 22034
rect 16212 21684 16264 21690
rect 16212 21626 16264 21632
rect 16684 21554 16712 23598
rect 16672 21548 16724 21554
rect 16672 21490 16724 21496
rect 17224 21548 17276 21554
rect 17224 21490 17276 21496
rect 15844 21480 15896 21486
rect 15844 21422 15896 21428
rect 15856 21010 15884 21422
rect 16212 21072 16264 21078
rect 16212 21014 16264 21020
rect 15844 21004 15896 21010
rect 15844 20946 15896 20952
rect 15660 20936 15712 20942
rect 15660 20878 15712 20884
rect 15568 20800 15620 20806
rect 15568 20742 15620 20748
rect 15108 20256 15160 20262
rect 15108 20198 15160 20204
rect 15016 19440 15068 19446
rect 15016 19382 15068 19388
rect 14280 19168 14332 19174
rect 14280 19110 14332 19116
rect 14292 18834 14320 19110
rect 15028 18902 15056 19382
rect 14648 18896 14700 18902
rect 14648 18838 14700 18844
rect 15016 18896 15068 18902
rect 15016 18838 15068 18844
rect 14280 18828 14332 18834
rect 14280 18770 14332 18776
rect 14464 17876 14516 17882
rect 14464 17818 14516 17824
rect 14372 17808 14424 17814
rect 14372 17750 14424 17756
rect 14384 17202 14412 17750
rect 14476 17610 14504 17818
rect 14660 17746 14688 18838
rect 14924 18828 14976 18834
rect 14924 18770 14976 18776
rect 14936 18222 14964 18770
rect 15016 18760 15068 18766
rect 15016 18702 15068 18708
rect 15028 18222 15056 18702
rect 14924 18216 14976 18222
rect 14924 18158 14976 18164
rect 15016 18216 15068 18222
rect 15016 18158 15068 18164
rect 15200 18148 15252 18154
rect 15200 18090 15252 18096
rect 14740 18080 14792 18086
rect 14740 18022 14792 18028
rect 15108 18080 15160 18086
rect 15108 18022 15160 18028
rect 14648 17740 14700 17746
rect 14648 17682 14700 17688
rect 14752 17678 14780 18022
rect 14924 17876 14976 17882
rect 14924 17818 14976 17824
rect 14740 17672 14792 17678
rect 14740 17614 14792 17620
rect 14464 17604 14516 17610
rect 14464 17546 14516 17552
rect 14556 17604 14608 17610
rect 14556 17546 14608 17552
rect 14372 17196 14424 17202
rect 14372 17138 14424 17144
rect 14280 17128 14332 17134
rect 14280 17070 14332 17076
rect 14292 16590 14320 17070
rect 14372 17060 14424 17066
rect 14372 17002 14424 17008
rect 14384 16794 14412 17002
rect 14568 16998 14596 17546
rect 14752 17134 14780 17614
rect 14936 17202 14964 17818
rect 14924 17196 14976 17202
rect 14924 17138 14976 17144
rect 14740 17128 14792 17134
rect 14740 17070 14792 17076
rect 15120 17082 15148 18022
rect 15212 17270 15240 18090
rect 15384 17876 15436 17882
rect 15384 17818 15436 17824
rect 15290 17640 15346 17649
rect 15290 17575 15292 17584
rect 15344 17575 15346 17584
rect 15292 17546 15344 17552
rect 15396 17542 15424 17818
rect 15580 17762 15608 20742
rect 15856 20262 15884 20946
rect 16028 20460 16080 20466
rect 16028 20402 16080 20408
rect 15844 20256 15896 20262
rect 15844 20198 15896 20204
rect 16040 19854 16068 20402
rect 16120 20392 16172 20398
rect 16120 20334 16172 20340
rect 15844 19848 15896 19854
rect 15844 19790 15896 19796
rect 16028 19848 16080 19854
rect 16028 19790 16080 19796
rect 15660 19372 15712 19378
rect 15660 19314 15712 19320
rect 15672 18154 15700 19314
rect 15856 19310 15884 19790
rect 16132 19378 16160 20334
rect 16224 19514 16252 21014
rect 16580 20936 16632 20942
rect 16578 20904 16580 20913
rect 16632 20904 16634 20913
rect 16304 20868 16356 20874
rect 16578 20839 16634 20848
rect 16304 20810 16356 20816
rect 16212 19508 16264 19514
rect 16212 19450 16264 19456
rect 16316 19446 16344 20810
rect 16580 20324 16632 20330
rect 16580 20266 16632 20272
rect 16592 19922 16620 20266
rect 16684 19990 16712 21490
rect 17236 21146 17264 21490
rect 17224 21140 17276 21146
rect 17224 21082 17276 21088
rect 16856 21072 16908 21078
rect 16856 21014 16908 21020
rect 16868 20942 16896 21014
rect 16856 20936 16908 20942
rect 16856 20878 16908 20884
rect 17132 20936 17184 20942
rect 17132 20878 17184 20884
rect 17144 20602 17172 20878
rect 17132 20596 17184 20602
rect 17132 20538 17184 20544
rect 17224 20256 17276 20262
rect 17224 20198 17276 20204
rect 16672 19984 16724 19990
rect 16672 19926 16724 19932
rect 16580 19916 16632 19922
rect 16580 19858 16632 19864
rect 16304 19440 16356 19446
rect 16304 19382 16356 19388
rect 16120 19372 16172 19378
rect 16120 19314 16172 19320
rect 15844 19304 15896 19310
rect 15844 19246 15896 19252
rect 15856 18290 15884 19246
rect 16132 18834 16160 19314
rect 16316 18834 16344 19382
rect 16120 18828 16172 18834
rect 16120 18770 16172 18776
rect 16304 18828 16356 18834
rect 16304 18770 16356 18776
rect 15936 18624 15988 18630
rect 15936 18566 15988 18572
rect 15948 18290 15976 18566
rect 16132 18408 16160 18770
rect 16212 18420 16264 18426
rect 16132 18380 16212 18408
rect 16212 18362 16264 18368
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 15936 18284 15988 18290
rect 15936 18226 15988 18232
rect 15660 18148 15712 18154
rect 15660 18090 15712 18096
rect 15580 17734 15700 17762
rect 15384 17536 15436 17542
rect 15384 17478 15436 17484
rect 15200 17264 15252 17270
rect 15200 17206 15252 17212
rect 15476 17196 15528 17202
rect 15476 17138 15528 17144
rect 15120 17054 15240 17082
rect 14556 16992 14608 16998
rect 14556 16934 14608 16940
rect 15108 16992 15160 16998
rect 15108 16934 15160 16940
rect 14372 16788 14424 16794
rect 14372 16730 14424 16736
rect 14464 16788 14516 16794
rect 14464 16730 14516 16736
rect 14476 16658 14504 16730
rect 14464 16652 14516 16658
rect 14464 16594 14516 16600
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 14292 16114 14320 16526
rect 14372 16176 14424 16182
rect 14372 16118 14424 16124
rect 14280 16108 14332 16114
rect 14280 16050 14332 16056
rect 14384 16046 14412 16118
rect 14372 16040 14424 16046
rect 14372 15982 14424 15988
rect 14280 15632 14332 15638
rect 14278 15600 14280 15609
rect 14332 15600 14334 15609
rect 14278 15535 14334 15544
rect 14292 15434 14320 15535
rect 14384 15502 14412 15982
rect 14464 15972 14516 15978
rect 14464 15914 14516 15920
rect 14372 15496 14424 15502
rect 14372 15438 14424 15444
rect 14280 15428 14332 15434
rect 14280 15370 14332 15376
rect 14292 15026 14320 15370
rect 14476 15366 14504 15914
rect 14464 15360 14516 15366
rect 14464 15302 14516 15308
rect 14188 15020 14240 15026
rect 14188 14962 14240 14968
rect 14280 15020 14332 15026
rect 14280 14962 14332 14968
rect 14096 14884 14148 14890
rect 14096 14826 14148 14832
rect 13820 14612 13872 14618
rect 13820 14554 13872 14560
rect 13544 14476 13596 14482
rect 13544 14418 13596 14424
rect 13452 14408 13504 14414
rect 13452 14350 13504 14356
rect 14108 13938 14136 14826
rect 14372 14272 14424 14278
rect 14372 14214 14424 14220
rect 14384 14006 14412 14214
rect 14372 14000 14424 14006
rect 14372 13942 14424 13948
rect 14096 13932 14148 13938
rect 14096 13874 14148 13880
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 12808 13320 12860 13326
rect 12808 13262 12860 13268
rect 12348 13184 12400 13190
rect 12348 13126 12400 13132
rect 12360 12918 12388 13126
rect 12820 12986 12848 13262
rect 12808 12980 12860 12986
rect 12808 12922 12860 12928
rect 12348 12912 12400 12918
rect 12348 12854 12400 12860
rect 12716 12776 12768 12782
rect 12716 12718 12768 12724
rect 12728 12442 12756 12718
rect 12716 12436 12768 12442
rect 12716 12378 12768 12384
rect 13648 6866 13676 13806
rect 13728 12776 13780 12782
rect 13728 12718 13780 12724
rect 13636 6860 13688 6866
rect 13636 6802 13688 6808
rect 12256 3120 12308 3126
rect 12256 3062 12308 3068
rect 13740 2514 13768 12718
rect 13820 12708 13872 12714
rect 13820 12650 13872 12656
rect 13832 12238 13860 12650
rect 14108 12306 14136 13874
rect 14096 12300 14148 12306
rect 14096 12242 14148 12248
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 14108 10674 14136 12242
rect 14568 11014 14596 16934
rect 15120 16794 15148 16934
rect 14924 16788 14976 16794
rect 14924 16730 14976 16736
rect 15108 16788 15160 16794
rect 15108 16730 15160 16736
rect 14936 15910 14964 16730
rect 15108 16584 15160 16590
rect 15212 16572 15240 17054
rect 15488 16726 15516 17138
rect 15476 16720 15528 16726
rect 15476 16662 15528 16668
rect 15160 16544 15240 16572
rect 15108 16526 15160 16532
rect 15476 16448 15528 16454
rect 15476 16390 15528 16396
rect 15488 16250 15516 16390
rect 15476 16244 15528 16250
rect 15476 16186 15528 16192
rect 14924 15904 14976 15910
rect 14924 15846 14976 15852
rect 15108 15904 15160 15910
rect 15108 15846 15160 15852
rect 15568 15904 15620 15910
rect 15568 15846 15620 15852
rect 15120 15706 15148 15846
rect 15108 15700 15160 15706
rect 15108 15642 15160 15648
rect 14648 15360 14700 15366
rect 14648 15302 14700 15308
rect 14660 15094 14688 15302
rect 15016 15156 15068 15162
rect 15016 15098 15068 15104
rect 14648 15088 14700 15094
rect 14648 15030 14700 15036
rect 15028 14414 15056 15098
rect 15120 15026 15148 15642
rect 15580 15586 15608 15846
rect 15396 15570 15608 15586
rect 15384 15564 15608 15570
rect 15436 15558 15608 15564
rect 15384 15506 15436 15512
rect 15200 15496 15252 15502
rect 15200 15438 15252 15444
rect 15212 15094 15240 15438
rect 15476 15360 15528 15366
rect 15476 15302 15528 15308
rect 15200 15088 15252 15094
rect 15200 15030 15252 15036
rect 15108 15020 15160 15026
rect 15108 14962 15160 14968
rect 15120 14414 15148 14962
rect 15212 14618 15240 15030
rect 15488 15026 15516 15302
rect 15476 15020 15528 15026
rect 15476 14962 15528 14968
rect 15200 14612 15252 14618
rect 15200 14554 15252 14560
rect 15580 14550 15608 15558
rect 15672 15502 15700 17734
rect 15856 17649 15884 18226
rect 15948 17814 15976 18226
rect 16120 17876 16172 17882
rect 16120 17818 16172 17824
rect 15936 17808 15988 17814
rect 15936 17750 15988 17756
rect 15842 17640 15898 17649
rect 15752 17604 15804 17610
rect 15842 17575 15898 17584
rect 15752 17546 15804 17552
rect 15764 17202 15792 17546
rect 15752 17196 15804 17202
rect 15752 17138 15804 17144
rect 15936 16584 15988 16590
rect 15936 16526 15988 16532
rect 15752 16448 15804 16454
rect 15752 16390 15804 16396
rect 15764 16114 15792 16390
rect 15752 16108 15804 16114
rect 15752 16050 15804 16056
rect 15764 15502 15792 16050
rect 15660 15496 15712 15502
rect 15660 15438 15712 15444
rect 15752 15496 15804 15502
rect 15752 15438 15804 15444
rect 15672 14550 15700 15438
rect 15948 14958 15976 16526
rect 16132 15609 16160 17818
rect 16118 15600 16174 15609
rect 16118 15535 16120 15544
rect 16172 15535 16174 15544
rect 16120 15506 16172 15512
rect 15936 14952 15988 14958
rect 15936 14894 15988 14900
rect 15568 14544 15620 14550
rect 15568 14486 15620 14492
rect 15660 14544 15712 14550
rect 15660 14486 15712 14492
rect 15016 14408 15068 14414
rect 15016 14350 15068 14356
rect 15108 14408 15160 14414
rect 15108 14350 15160 14356
rect 15672 14006 15700 14486
rect 15948 14414 15976 14894
rect 15936 14408 15988 14414
rect 15936 14350 15988 14356
rect 15948 14074 15976 14350
rect 15936 14068 15988 14074
rect 15936 14010 15988 14016
rect 15660 14000 15712 14006
rect 15660 13942 15712 13948
rect 16316 13462 16344 18770
rect 16592 18290 16620 19858
rect 16948 19168 17000 19174
rect 16948 19110 17000 19116
rect 16960 18766 16988 19110
rect 16948 18760 17000 18766
rect 16948 18702 17000 18708
rect 16672 18692 16724 18698
rect 16672 18634 16724 18640
rect 16580 18284 16632 18290
rect 16580 18226 16632 18232
rect 16488 18080 16540 18086
rect 16488 18022 16540 18028
rect 16500 17610 16528 18022
rect 16684 17610 16712 18634
rect 16960 18290 16988 18702
rect 16948 18284 17000 18290
rect 16948 18226 17000 18232
rect 16488 17604 16540 17610
rect 16488 17546 16540 17552
rect 16672 17604 16724 17610
rect 16672 17546 16724 17552
rect 16500 16794 16528 17546
rect 17132 17536 17184 17542
rect 17132 17478 17184 17484
rect 16948 17128 17000 17134
rect 16948 17070 17000 17076
rect 16580 16992 16632 16998
rect 16580 16934 16632 16940
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 16488 16788 16540 16794
rect 16488 16730 16540 16736
rect 16592 16590 16620 16934
rect 16580 16584 16632 16590
rect 16580 16526 16632 16532
rect 16396 15496 16448 15502
rect 16396 15438 16448 15444
rect 16408 15026 16436 15438
rect 16396 15020 16448 15026
rect 16396 14962 16448 14968
rect 16408 14346 16436 14962
rect 16396 14340 16448 14346
rect 16396 14282 16448 14288
rect 15200 13456 15252 13462
rect 15200 13398 15252 13404
rect 16304 13456 16356 13462
rect 16304 13398 16356 13404
rect 15212 12850 15240 13398
rect 16120 13320 16172 13326
rect 16120 13262 16172 13268
rect 15200 12844 15252 12850
rect 15200 12786 15252 12792
rect 15936 12776 15988 12782
rect 15936 12718 15988 12724
rect 14740 12164 14792 12170
rect 14740 12106 14792 12112
rect 14752 11898 14780 12106
rect 14740 11892 14792 11898
rect 14740 11834 14792 11840
rect 14556 11008 14608 11014
rect 14556 10950 14608 10956
rect 14096 10668 14148 10674
rect 14096 10610 14148 10616
rect 14740 10668 14792 10674
rect 14740 10610 14792 10616
rect 14832 10668 14884 10674
rect 14832 10610 14884 10616
rect 14752 10130 14780 10610
rect 14844 10266 14872 10610
rect 15948 10266 15976 12718
rect 16132 12442 16160 13262
rect 16408 13190 16436 14282
rect 16684 14278 16712 16934
rect 16960 16658 16988 17070
rect 17144 16998 17172 17478
rect 17236 17202 17264 20198
rect 17420 18766 17448 24754
rect 17684 23724 17736 23730
rect 17684 23666 17736 23672
rect 17696 22778 17724 23666
rect 17880 23186 17908 25910
rect 17960 25900 18012 25906
rect 17960 25842 18012 25848
rect 17972 24682 18000 25842
rect 17960 24676 18012 24682
rect 17960 24618 18012 24624
rect 18156 24274 18184 27338
rect 18616 24614 18644 27542
rect 18708 25906 18736 29174
rect 18788 28076 18840 28082
rect 18788 28018 18840 28024
rect 18800 27402 18828 28018
rect 18984 27878 19012 29582
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 19432 29232 19484 29238
rect 19432 29174 19484 29180
rect 19444 28626 19472 29174
rect 19432 28620 19484 28626
rect 19432 28562 19484 28568
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 18972 27872 19024 27878
rect 18972 27814 19024 27820
rect 18788 27396 18840 27402
rect 18788 27338 18840 27344
rect 18696 25900 18748 25906
rect 18696 25842 18748 25848
rect 18708 24818 18736 25842
rect 18696 24812 18748 24818
rect 18696 24754 18748 24760
rect 18604 24608 18656 24614
rect 18604 24550 18656 24556
rect 18144 24268 18196 24274
rect 18144 24210 18196 24216
rect 18052 24064 18104 24070
rect 18052 24006 18104 24012
rect 17868 23180 17920 23186
rect 17868 23122 17920 23128
rect 17684 22772 17736 22778
rect 17684 22714 17736 22720
rect 17880 22166 17908 23122
rect 18064 22642 18092 24006
rect 18156 23118 18184 24210
rect 18144 23112 18196 23118
rect 18144 23054 18196 23060
rect 18052 22636 18104 22642
rect 18052 22578 18104 22584
rect 17868 22160 17920 22166
rect 17868 22102 17920 22108
rect 18156 22030 18184 23054
rect 18604 22636 18656 22642
rect 18604 22578 18656 22584
rect 18616 22234 18644 22578
rect 18604 22228 18656 22234
rect 18604 22170 18656 22176
rect 17960 22024 18012 22030
rect 17960 21966 18012 21972
rect 18144 22024 18196 22030
rect 18144 21966 18196 21972
rect 17592 21344 17644 21350
rect 17592 21286 17644 21292
rect 17604 20913 17632 21286
rect 17684 21072 17736 21078
rect 17684 21014 17736 21020
rect 17590 20904 17646 20913
rect 17590 20839 17592 20848
rect 17644 20839 17646 20848
rect 17592 20810 17644 20816
rect 17604 20398 17632 20810
rect 17696 20466 17724 21014
rect 17972 20942 18000 21966
rect 18788 21548 18840 21554
rect 18788 21490 18840 21496
rect 17960 20936 18012 20942
rect 17960 20878 18012 20884
rect 17684 20460 17736 20466
rect 17684 20402 17736 20408
rect 17592 20392 17644 20398
rect 17592 20334 17644 20340
rect 17960 20392 18012 20398
rect 17960 20334 18012 20340
rect 17776 19984 17828 19990
rect 17776 19926 17828 19932
rect 17788 19378 17816 19926
rect 17776 19372 17828 19378
rect 17776 19314 17828 19320
rect 17408 18760 17460 18766
rect 17408 18702 17460 18708
rect 17592 18692 17644 18698
rect 17592 18634 17644 18640
rect 17604 17882 17632 18634
rect 17592 17876 17644 17882
rect 17592 17818 17644 17824
rect 17972 17746 18000 20334
rect 18800 19990 18828 21490
rect 18880 20256 18932 20262
rect 18880 20198 18932 20204
rect 18788 19984 18840 19990
rect 18788 19926 18840 19932
rect 18892 19378 18920 20198
rect 18052 19372 18104 19378
rect 18052 19314 18104 19320
rect 18880 19372 18932 19378
rect 18880 19314 18932 19320
rect 18064 18970 18092 19314
rect 18696 19168 18748 19174
rect 18696 19110 18748 19116
rect 18052 18964 18104 18970
rect 18052 18906 18104 18912
rect 18708 18290 18736 19110
rect 18880 18692 18932 18698
rect 18880 18634 18932 18640
rect 18892 18290 18920 18634
rect 18052 18284 18104 18290
rect 18052 18226 18104 18232
rect 18696 18284 18748 18290
rect 18696 18226 18748 18232
rect 18880 18284 18932 18290
rect 18880 18226 18932 18232
rect 17960 17740 18012 17746
rect 17960 17682 18012 17688
rect 17868 17672 17920 17678
rect 17868 17614 17920 17620
rect 17880 17270 17908 17614
rect 17960 17332 18012 17338
rect 17960 17274 18012 17280
rect 17868 17264 17920 17270
rect 17868 17206 17920 17212
rect 17224 17196 17276 17202
rect 17224 17138 17276 17144
rect 17132 16992 17184 16998
rect 17132 16934 17184 16940
rect 17972 16810 18000 17274
rect 18064 17218 18092 18226
rect 18328 17672 18380 17678
rect 18328 17614 18380 17620
rect 18064 17202 18276 17218
rect 18064 17196 18288 17202
rect 18064 17190 18236 17196
rect 18064 16998 18092 17190
rect 18236 17138 18288 17144
rect 18052 16992 18104 16998
rect 18052 16934 18104 16940
rect 17972 16782 18092 16810
rect 17960 16720 18012 16726
rect 17960 16662 18012 16668
rect 16948 16652 17000 16658
rect 16948 16594 17000 16600
rect 17684 16652 17736 16658
rect 17684 16594 17736 16600
rect 17040 16516 17092 16522
rect 17040 16458 17092 16464
rect 17052 15502 17080 16458
rect 17696 16046 17724 16594
rect 17972 16114 18000 16662
rect 18064 16590 18092 16782
rect 18052 16584 18104 16590
rect 18052 16526 18104 16532
rect 18144 16244 18196 16250
rect 18144 16186 18196 16192
rect 17960 16108 18012 16114
rect 17960 16050 18012 16056
rect 17684 16040 17736 16046
rect 17684 15982 17736 15988
rect 18156 15706 18184 16186
rect 18144 15700 18196 15706
rect 18144 15642 18196 15648
rect 18340 15502 18368 17614
rect 18892 17218 18920 18226
rect 18984 17898 19012 27814
rect 20180 27606 20208 31726
rect 20352 31340 20404 31346
rect 20352 31282 20404 31288
rect 20364 31142 20392 31282
rect 20352 31136 20404 31142
rect 20352 31078 20404 31084
rect 20260 28484 20312 28490
rect 20260 28426 20312 28432
rect 20272 28218 20300 28426
rect 20260 28212 20312 28218
rect 20260 28154 20312 28160
rect 20364 28150 20392 31078
rect 20548 30598 20576 31758
rect 20640 30734 20668 31894
rect 20628 30728 20680 30734
rect 20628 30670 20680 30676
rect 20536 30592 20588 30598
rect 20536 30534 20588 30540
rect 20444 29640 20496 29646
rect 20444 29582 20496 29588
rect 20456 29238 20484 29582
rect 20548 29578 20576 30534
rect 20536 29572 20588 29578
rect 20536 29514 20588 29520
rect 20640 29510 20668 30670
rect 20732 30190 20760 32234
rect 20824 31822 20852 32778
rect 21284 32570 21312 33526
rect 21272 32564 21324 32570
rect 21272 32506 21324 32512
rect 20812 31816 20864 31822
rect 20864 31764 20944 31770
rect 20812 31758 20944 31764
rect 20824 31754 20944 31758
rect 20824 31742 21036 31754
rect 20916 31726 21036 31742
rect 20812 31680 20864 31686
rect 20812 31622 20864 31628
rect 20824 31346 20852 31622
rect 20812 31340 20864 31346
rect 20812 31282 20864 31288
rect 21008 30870 21036 31726
rect 21364 31272 21416 31278
rect 21364 31214 21416 31220
rect 21548 31272 21600 31278
rect 21548 31214 21600 31220
rect 21376 30938 21404 31214
rect 21364 30932 21416 30938
rect 21364 30874 21416 30880
rect 20996 30864 21048 30870
rect 20996 30806 21048 30812
rect 20812 30796 20864 30802
rect 20812 30738 20864 30744
rect 20720 30184 20772 30190
rect 20720 30126 20772 30132
rect 20824 30054 20852 30738
rect 21008 30734 21036 30806
rect 20996 30728 21048 30734
rect 20996 30670 21048 30676
rect 21376 30394 21404 30874
rect 21560 30734 21588 31214
rect 21548 30728 21600 30734
rect 21548 30670 21600 30676
rect 21364 30388 21416 30394
rect 21364 30330 21416 30336
rect 21560 30326 21588 30670
rect 21548 30320 21600 30326
rect 21548 30262 21600 30268
rect 20812 30048 20864 30054
rect 20812 29990 20864 29996
rect 20996 30048 21048 30054
rect 20996 29990 21048 29996
rect 20812 29572 20864 29578
rect 20812 29514 20864 29520
rect 20628 29504 20680 29510
rect 20628 29446 20680 29452
rect 20824 29306 20852 29514
rect 20812 29300 20864 29306
rect 20812 29242 20864 29248
rect 20444 29232 20496 29238
rect 20444 29174 20496 29180
rect 21008 29170 21036 29990
rect 20904 29164 20956 29170
rect 20904 29106 20956 29112
rect 20996 29164 21048 29170
rect 20996 29106 21048 29112
rect 20916 28762 20944 29106
rect 20904 28756 20956 28762
rect 20904 28698 20956 28704
rect 21180 28416 21232 28422
rect 21180 28358 21232 28364
rect 20352 28144 20404 28150
rect 20352 28086 20404 28092
rect 20444 28076 20496 28082
rect 20444 28018 20496 28024
rect 20456 27674 20484 28018
rect 21192 27674 21220 28358
rect 20444 27668 20496 27674
rect 20444 27610 20496 27616
rect 21180 27668 21232 27674
rect 21180 27610 21232 27616
rect 20168 27600 20220 27606
rect 20168 27542 20220 27548
rect 21192 27470 21220 27610
rect 20812 27464 20864 27470
rect 20812 27406 20864 27412
rect 21180 27464 21232 27470
rect 21180 27406 21232 27412
rect 21456 27464 21508 27470
rect 21456 27406 21508 27412
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 19432 27124 19484 27130
rect 19432 27066 19484 27072
rect 19444 26790 19472 27066
rect 20824 27062 20852 27406
rect 20996 27396 21048 27402
rect 20996 27338 21048 27344
rect 20812 27056 20864 27062
rect 20812 26998 20864 27004
rect 19524 26988 19576 26994
rect 19524 26930 19576 26936
rect 19432 26784 19484 26790
rect 19432 26726 19484 26732
rect 19444 26450 19472 26726
rect 19536 26586 19564 26930
rect 19708 26784 19760 26790
rect 19708 26726 19760 26732
rect 19524 26580 19576 26586
rect 19524 26522 19576 26528
rect 19432 26444 19484 26450
rect 19432 26386 19484 26392
rect 19720 26382 19748 26726
rect 20824 26586 20852 26998
rect 21008 26926 21036 27338
rect 20996 26920 21048 26926
rect 20996 26862 21048 26868
rect 20812 26580 20864 26586
rect 20812 26522 20864 26528
rect 19708 26376 19760 26382
rect 19708 26318 19760 26324
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 20824 26042 20852 26522
rect 21008 26382 21036 26862
rect 20996 26376 21048 26382
rect 20996 26318 21048 26324
rect 20812 26036 20864 26042
rect 20812 25978 20864 25984
rect 21192 25974 21220 27406
rect 21468 26382 21496 27406
rect 21456 26376 21508 26382
rect 21508 26336 21588 26364
rect 21456 26318 21508 26324
rect 21560 26246 21588 26336
rect 21548 26240 21600 26246
rect 21548 26182 21600 26188
rect 21560 26042 21588 26182
rect 21548 26036 21600 26042
rect 21548 25978 21600 25984
rect 21180 25968 21232 25974
rect 21180 25910 21232 25916
rect 21456 25968 21508 25974
rect 21456 25910 21508 25916
rect 20812 25288 20864 25294
rect 20812 25230 20864 25236
rect 20168 25152 20220 25158
rect 20168 25094 20220 25100
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 19616 24812 19668 24818
rect 19616 24754 19668 24760
rect 19628 24410 19656 24754
rect 19616 24404 19668 24410
rect 19616 24346 19668 24352
rect 20180 24274 20208 25094
rect 20824 24410 20852 25230
rect 21272 25220 21324 25226
rect 21272 25162 21324 25168
rect 21284 24750 21312 25162
rect 21272 24744 21324 24750
rect 21272 24686 21324 24692
rect 20904 24608 20956 24614
rect 20904 24550 20956 24556
rect 20812 24404 20864 24410
rect 20812 24346 20864 24352
rect 20168 24268 20220 24274
rect 20168 24210 20220 24216
rect 20628 24268 20680 24274
rect 20628 24210 20680 24216
rect 20076 24200 20128 24206
rect 20076 24142 20128 24148
rect 19432 24132 19484 24138
rect 19432 24074 19484 24080
rect 19444 23322 19472 24074
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 20088 23866 20116 24142
rect 20076 23860 20128 23866
rect 20076 23802 20128 23808
rect 19800 23588 19852 23594
rect 19800 23530 19852 23536
rect 19432 23316 19484 23322
rect 19432 23258 19484 23264
rect 19812 23118 19840 23530
rect 20180 23186 20208 24210
rect 20640 23730 20668 24210
rect 20824 24206 20852 24346
rect 20916 24342 20944 24550
rect 20904 24336 20956 24342
rect 20904 24278 20956 24284
rect 21180 24336 21232 24342
rect 21180 24278 21232 24284
rect 20812 24200 20864 24206
rect 20812 24142 20864 24148
rect 20812 24064 20864 24070
rect 20812 24006 20864 24012
rect 21088 24064 21140 24070
rect 21088 24006 21140 24012
rect 20628 23724 20680 23730
rect 20628 23666 20680 23672
rect 20720 23724 20772 23730
rect 20720 23666 20772 23672
rect 20168 23180 20220 23186
rect 20168 23122 20220 23128
rect 19800 23112 19852 23118
rect 19800 23054 19852 23060
rect 20640 23050 20668 23666
rect 20732 23118 20760 23666
rect 20824 23662 20852 24006
rect 21100 23662 21128 24006
rect 21192 23662 21220 24278
rect 21284 23798 21312 24686
rect 21272 23792 21324 23798
rect 21272 23734 21324 23740
rect 20812 23656 20864 23662
rect 20812 23598 20864 23604
rect 21088 23656 21140 23662
rect 21088 23598 21140 23604
rect 21180 23656 21232 23662
rect 21180 23598 21232 23604
rect 20824 23322 20852 23598
rect 20904 23520 20956 23526
rect 20904 23462 20956 23468
rect 20812 23316 20864 23322
rect 20812 23258 20864 23264
rect 20720 23112 20772 23118
rect 20720 23054 20772 23060
rect 20916 23050 20944 23462
rect 21192 23050 21220 23598
rect 21364 23588 21416 23594
rect 21364 23530 21416 23536
rect 20628 23044 20680 23050
rect 20628 22986 20680 22992
rect 20904 23044 20956 23050
rect 20904 22986 20956 22992
rect 21180 23044 21232 23050
rect 21180 22986 21232 22992
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 20640 22778 20668 22986
rect 20628 22772 20680 22778
rect 20628 22714 20680 22720
rect 20916 22642 20944 22986
rect 20904 22636 20956 22642
rect 20904 22578 20956 22584
rect 19064 22432 19116 22438
rect 19064 22374 19116 22380
rect 19076 21622 19104 22374
rect 20720 22160 20772 22166
rect 20720 22102 20772 22108
rect 19984 21888 20036 21894
rect 19984 21830 20036 21836
rect 20628 21888 20680 21894
rect 20628 21830 20680 21836
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19064 21616 19116 21622
rect 19064 21558 19116 21564
rect 19996 20874 20024 21830
rect 19984 20868 20036 20874
rect 19984 20810 20036 20816
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19340 20392 19392 20398
rect 19340 20334 19392 20340
rect 19996 20346 20024 20810
rect 20076 20800 20128 20806
rect 20076 20742 20128 20748
rect 20088 20534 20116 20742
rect 20076 20528 20128 20534
rect 20076 20470 20128 20476
rect 19352 19854 19380 20334
rect 19996 20318 20116 20346
rect 19996 20262 20024 20318
rect 19984 20256 20036 20262
rect 19984 20198 20036 20204
rect 19340 19848 19392 19854
rect 19340 19790 19392 19796
rect 19432 19780 19484 19786
rect 19432 19722 19484 19728
rect 19340 19712 19392 19718
rect 19340 19654 19392 19660
rect 19352 19514 19380 19654
rect 19340 19508 19392 19514
rect 19340 19450 19392 19456
rect 19444 18970 19472 19722
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 19432 18964 19484 18970
rect 19432 18906 19484 18912
rect 20088 18902 20116 20318
rect 20076 18896 20128 18902
rect 20076 18838 20128 18844
rect 19984 18624 20036 18630
rect 19984 18566 20036 18572
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19996 18290 20024 18566
rect 19984 18284 20036 18290
rect 19984 18226 20036 18232
rect 20088 18154 20116 18838
rect 20076 18148 20128 18154
rect 20076 18090 20128 18096
rect 20168 18080 20220 18086
rect 20168 18022 20220 18028
rect 18984 17870 19104 17898
rect 18972 17740 19024 17746
rect 18972 17682 19024 17688
rect 18984 17338 19012 17682
rect 18972 17332 19024 17338
rect 18972 17274 19024 17280
rect 18892 17202 19012 17218
rect 18892 17196 19024 17202
rect 18892 17190 18972 17196
rect 18972 17138 19024 17144
rect 18420 16992 18472 16998
rect 18420 16934 18472 16940
rect 18432 16794 18460 16934
rect 18420 16788 18472 16794
rect 18420 16730 18472 16736
rect 17040 15496 17092 15502
rect 17040 15438 17092 15444
rect 17408 15496 17460 15502
rect 17408 15438 17460 15444
rect 18052 15496 18104 15502
rect 18052 15438 18104 15444
rect 18328 15496 18380 15502
rect 18328 15438 18380 15444
rect 17420 15162 17448 15438
rect 17408 15156 17460 15162
rect 17408 15098 17460 15104
rect 17420 14482 17448 15098
rect 17960 14816 18012 14822
rect 17960 14758 18012 14764
rect 17408 14476 17460 14482
rect 17408 14418 17460 14424
rect 16672 14272 16724 14278
rect 16672 14214 16724 14220
rect 16580 14000 16632 14006
rect 16580 13942 16632 13948
rect 16592 13326 16620 13942
rect 16948 13864 17000 13870
rect 16948 13806 17000 13812
rect 16856 13728 16908 13734
rect 16856 13670 16908 13676
rect 16868 13394 16896 13670
rect 16672 13388 16724 13394
rect 16856 13388 16908 13394
rect 16724 13348 16856 13376
rect 16672 13330 16724 13336
rect 16856 13330 16908 13336
rect 16580 13320 16632 13326
rect 16580 13262 16632 13268
rect 16488 13252 16540 13258
rect 16488 13194 16540 13200
rect 16396 13184 16448 13190
rect 16396 13126 16448 13132
rect 16304 12844 16356 12850
rect 16304 12786 16356 12792
rect 16316 12714 16344 12786
rect 16408 12730 16436 13126
rect 16500 12850 16528 13194
rect 16488 12844 16540 12850
rect 16488 12786 16540 12792
rect 16304 12708 16356 12714
rect 16408 12702 16528 12730
rect 16304 12650 16356 12656
rect 16120 12436 16172 12442
rect 16120 12378 16172 12384
rect 16316 12238 16344 12650
rect 16304 12232 16356 12238
rect 16304 12174 16356 12180
rect 16304 12096 16356 12102
rect 16304 12038 16356 12044
rect 16316 11762 16344 12038
rect 16500 11762 16528 12702
rect 16592 12442 16620 13262
rect 16684 12646 16712 13330
rect 16960 12782 16988 13806
rect 17868 13728 17920 13734
rect 17868 13670 17920 13676
rect 17880 13462 17908 13670
rect 17868 13456 17920 13462
rect 17868 13398 17920 13404
rect 17224 12912 17276 12918
rect 17224 12854 17276 12860
rect 16948 12776 17000 12782
rect 16948 12718 17000 12724
rect 16672 12640 16724 12646
rect 16672 12582 16724 12588
rect 16580 12436 16632 12442
rect 16580 12378 16632 12384
rect 16960 12238 16988 12718
rect 17236 12442 17264 12854
rect 17224 12436 17276 12442
rect 17224 12378 17276 12384
rect 16948 12232 17000 12238
rect 16948 12174 17000 12180
rect 17236 11898 17264 12378
rect 17880 12374 17908 13398
rect 17972 12850 18000 14758
rect 18064 14482 18092 15438
rect 18340 15026 18368 15438
rect 18420 15360 18472 15366
rect 18420 15302 18472 15308
rect 18328 15020 18380 15026
rect 18328 14962 18380 14968
rect 18432 14890 18460 15302
rect 19076 15094 19104 17870
rect 20076 17672 20128 17678
rect 20076 17614 20128 17620
rect 19984 17604 20036 17610
rect 19984 17546 20036 17552
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 19996 17134 20024 17546
rect 20088 17202 20116 17614
rect 20180 17610 20208 18022
rect 20168 17604 20220 17610
rect 20168 17546 20220 17552
rect 20076 17196 20128 17202
rect 20076 17138 20128 17144
rect 19984 17128 20036 17134
rect 19984 17070 20036 17076
rect 19248 16992 19300 16998
rect 19248 16934 19300 16940
rect 19260 16590 19288 16934
rect 20088 16590 20116 17138
rect 20640 17134 20668 21830
rect 20732 21622 20760 22102
rect 20916 22030 20944 22578
rect 21376 22030 21404 23530
rect 21468 22710 21496 25910
rect 21560 23866 21588 25978
rect 21548 23860 21600 23866
rect 21548 23802 21600 23808
rect 21456 22704 21508 22710
rect 21456 22646 21508 22652
rect 20904 22024 20956 22030
rect 20904 21966 20956 21972
rect 21364 22024 21416 22030
rect 21364 21966 21416 21972
rect 20916 21690 20944 21966
rect 20904 21684 20956 21690
rect 20904 21626 20956 21632
rect 20720 21616 20772 21622
rect 20720 21558 20772 21564
rect 20812 21344 20864 21350
rect 20812 21286 20864 21292
rect 20824 21146 20852 21286
rect 20812 21140 20864 21146
rect 20812 21082 20864 21088
rect 20720 21004 20772 21010
rect 20720 20946 20772 20952
rect 20732 19990 20760 20946
rect 21088 20936 21140 20942
rect 21088 20878 21140 20884
rect 20812 20868 20864 20874
rect 20812 20810 20864 20816
rect 20720 19984 20772 19990
rect 20720 19926 20772 19932
rect 20824 19122 20852 20810
rect 21100 20602 21128 20878
rect 21272 20800 21324 20806
rect 21272 20742 21324 20748
rect 21088 20596 21140 20602
rect 21088 20538 21140 20544
rect 20732 19094 20852 19122
rect 20628 17128 20680 17134
rect 20628 17070 20680 17076
rect 19248 16584 19300 16590
rect 19248 16526 19300 16532
rect 20076 16584 20128 16590
rect 20076 16526 20128 16532
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 19340 16040 19392 16046
rect 19340 15982 19392 15988
rect 19352 15434 19380 15982
rect 19432 15564 19484 15570
rect 19432 15506 19484 15512
rect 19340 15428 19392 15434
rect 19340 15370 19392 15376
rect 19352 15178 19380 15370
rect 19260 15150 19380 15178
rect 19064 15088 19116 15094
rect 19064 15030 19116 15036
rect 18420 14884 18472 14890
rect 18420 14826 18472 14832
rect 18052 14476 18104 14482
rect 18052 14418 18104 14424
rect 18328 13864 18380 13870
rect 18328 13806 18380 13812
rect 18052 13184 18104 13190
rect 18052 13126 18104 13132
rect 18064 12918 18092 13126
rect 18052 12912 18104 12918
rect 18052 12854 18104 12860
rect 17960 12844 18012 12850
rect 17960 12786 18012 12792
rect 17868 12368 17920 12374
rect 17868 12310 17920 12316
rect 18340 12238 18368 13806
rect 18328 12232 18380 12238
rect 18328 12174 18380 12180
rect 17500 12164 17552 12170
rect 17500 12106 17552 12112
rect 17224 11892 17276 11898
rect 17224 11834 17276 11840
rect 16304 11756 16356 11762
rect 16304 11698 16356 11704
rect 16488 11756 16540 11762
rect 16488 11698 16540 11704
rect 17236 11150 17264 11834
rect 17512 11150 17540 12106
rect 19156 12096 19208 12102
rect 19156 12038 19208 12044
rect 18236 11688 18288 11694
rect 18236 11630 18288 11636
rect 17224 11144 17276 11150
rect 17224 11086 17276 11092
rect 17500 11144 17552 11150
rect 17500 11086 17552 11092
rect 17132 11008 17184 11014
rect 17132 10950 17184 10956
rect 17316 11008 17368 11014
rect 17316 10950 17368 10956
rect 16948 10600 17000 10606
rect 16948 10542 17000 10548
rect 16488 10532 16540 10538
rect 16488 10474 16540 10480
rect 16500 10266 16528 10474
rect 14832 10260 14884 10266
rect 14832 10202 14884 10208
rect 15936 10260 15988 10266
rect 15936 10202 15988 10208
rect 16488 10260 16540 10266
rect 16488 10202 16540 10208
rect 14740 10124 14792 10130
rect 14740 10066 14792 10072
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 14752 8498 14780 10066
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 15660 10056 15712 10062
rect 15660 9998 15712 10004
rect 15396 9586 15424 9998
rect 15476 9988 15528 9994
rect 15476 9930 15528 9936
rect 15488 9654 15516 9930
rect 15672 9654 15700 9998
rect 16120 9920 16172 9926
rect 16120 9862 16172 9868
rect 16488 9920 16540 9926
rect 16488 9862 16540 9868
rect 15476 9648 15528 9654
rect 15476 9590 15528 9596
rect 15660 9648 15712 9654
rect 15660 9590 15712 9596
rect 15384 9580 15436 9586
rect 15384 9522 15436 9528
rect 15396 8974 15424 9522
rect 15936 9512 15988 9518
rect 15936 9454 15988 9460
rect 15384 8968 15436 8974
rect 15384 8910 15436 8916
rect 15660 8968 15712 8974
rect 15660 8910 15712 8916
rect 15568 8832 15620 8838
rect 15568 8774 15620 8780
rect 15580 8566 15608 8774
rect 15568 8560 15620 8566
rect 15568 8502 15620 8508
rect 14740 8492 14792 8498
rect 14740 8434 14792 8440
rect 15672 8090 15700 8910
rect 15660 8084 15712 8090
rect 15660 8026 15712 8032
rect 15948 7954 15976 9454
rect 16132 9450 16160 9862
rect 16304 9580 16356 9586
rect 16304 9522 16356 9528
rect 16120 9444 16172 9450
rect 16120 9386 16172 9392
rect 16132 8974 16160 9386
rect 16316 8974 16344 9522
rect 16500 9042 16528 9862
rect 16488 9036 16540 9042
rect 16488 8978 16540 8984
rect 16120 8968 16172 8974
rect 16120 8910 16172 8916
rect 16304 8968 16356 8974
rect 16304 8910 16356 8916
rect 16132 8634 16160 8910
rect 16120 8628 16172 8634
rect 16120 8570 16172 8576
rect 15936 7948 15988 7954
rect 15936 7890 15988 7896
rect 16132 7886 16160 8570
rect 16316 8566 16344 8910
rect 16304 8560 16356 8566
rect 16304 8502 16356 8508
rect 16316 8090 16344 8502
rect 16304 8084 16356 8090
rect 16304 8026 16356 8032
rect 16868 7954 16896 10066
rect 16960 9654 16988 10542
rect 16948 9648 17000 9654
rect 16948 9590 17000 9596
rect 17144 9518 17172 10950
rect 17328 10130 17356 10950
rect 17512 10266 17540 11086
rect 18144 10736 18196 10742
rect 18144 10678 18196 10684
rect 18052 10464 18104 10470
rect 18052 10406 18104 10412
rect 17500 10260 17552 10266
rect 17500 10202 17552 10208
rect 17316 10124 17368 10130
rect 17316 10066 17368 10072
rect 17960 9988 18012 9994
rect 17960 9930 18012 9936
rect 17132 9512 17184 9518
rect 17132 9454 17184 9460
rect 17144 8430 17172 9454
rect 17972 9178 18000 9930
rect 17960 9172 18012 9178
rect 17960 9114 18012 9120
rect 17868 9104 17920 9110
rect 17868 9046 17920 9052
rect 17880 8498 17908 9046
rect 18064 8974 18092 10406
rect 18156 9722 18184 10678
rect 18248 10538 18276 11630
rect 18512 11144 18564 11150
rect 18512 11086 18564 11092
rect 18524 10674 18552 11086
rect 19168 11082 19196 12038
rect 19156 11076 19208 11082
rect 19156 11018 19208 11024
rect 19260 11014 19288 15150
rect 19444 14414 19472 15506
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 20088 15026 20116 16526
rect 20732 16250 20760 19094
rect 20812 18964 20864 18970
rect 20812 18906 20864 18912
rect 20824 18698 20852 18906
rect 20904 18760 20956 18766
rect 20904 18702 20956 18708
rect 20812 18692 20864 18698
rect 20812 18634 20864 18640
rect 20720 16244 20772 16250
rect 20720 16186 20772 16192
rect 20732 15570 20760 16186
rect 20720 15564 20772 15570
rect 20720 15506 20772 15512
rect 20824 15502 20852 18634
rect 20916 17678 20944 18702
rect 20996 18692 21048 18698
rect 20996 18634 21048 18640
rect 20904 17672 20956 17678
rect 20904 17614 20956 17620
rect 20812 15496 20864 15502
rect 20812 15438 20864 15444
rect 20720 15428 20772 15434
rect 20720 15370 20772 15376
rect 20536 15360 20588 15366
rect 20536 15302 20588 15308
rect 20444 15088 20496 15094
rect 20444 15030 20496 15036
rect 20076 15020 20128 15026
rect 20076 14962 20128 14968
rect 19616 14816 19668 14822
rect 19616 14758 19668 14764
rect 19628 14618 19656 14758
rect 19616 14612 19668 14618
rect 19616 14554 19668 14560
rect 20168 14476 20220 14482
rect 20168 14418 20220 14424
rect 19432 14408 19484 14414
rect 19432 14350 19484 14356
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 20180 14006 20208 14418
rect 20456 14414 20484 15030
rect 20548 15026 20576 15302
rect 20536 15020 20588 15026
rect 20536 14962 20588 14968
rect 20260 14408 20312 14414
rect 20260 14350 20312 14356
rect 20444 14408 20496 14414
rect 20444 14350 20496 14356
rect 20272 14074 20300 14350
rect 20444 14272 20496 14278
rect 20444 14214 20496 14220
rect 20260 14068 20312 14074
rect 20260 14010 20312 14016
rect 20168 14000 20220 14006
rect 20168 13942 20220 13948
rect 19984 13932 20036 13938
rect 19984 13874 20036 13880
rect 19996 13734 20024 13874
rect 19984 13728 20036 13734
rect 19984 13670 20036 13676
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 20180 12442 20208 13942
rect 20352 13932 20404 13938
rect 20352 13874 20404 13880
rect 20364 13802 20392 13874
rect 20352 13796 20404 13802
rect 20352 13738 20404 13744
rect 20456 13734 20484 14214
rect 20732 14006 20760 15370
rect 21008 14618 21036 18634
rect 21180 16652 21232 16658
rect 21180 16594 21232 16600
rect 21192 16182 21220 16594
rect 21180 16176 21232 16182
rect 21180 16118 21232 16124
rect 20996 14612 21048 14618
rect 20996 14554 21048 14560
rect 20720 14000 20772 14006
rect 20720 13942 20772 13948
rect 20720 13864 20772 13870
rect 20720 13806 20772 13812
rect 20444 13728 20496 13734
rect 20444 13670 20496 13676
rect 20260 13388 20312 13394
rect 20260 13330 20312 13336
rect 20272 12986 20300 13330
rect 20260 12980 20312 12986
rect 20260 12922 20312 12928
rect 20352 12844 20404 12850
rect 20352 12786 20404 12792
rect 20364 12442 20392 12786
rect 20168 12436 20220 12442
rect 20168 12378 20220 12384
rect 20352 12436 20404 12442
rect 20352 12378 20404 12384
rect 19340 12368 19392 12374
rect 19340 12310 19392 12316
rect 19352 11558 19380 12310
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 20364 11898 20392 12378
rect 20456 12306 20484 13670
rect 20732 13326 20760 13806
rect 20720 13320 20772 13326
rect 20720 13262 20772 13268
rect 20536 13184 20588 13190
rect 20536 13126 20588 13132
rect 20548 12714 20576 13126
rect 21180 12980 21232 12986
rect 21180 12922 21232 12928
rect 21088 12844 21140 12850
rect 21088 12786 21140 12792
rect 20536 12708 20588 12714
rect 20536 12650 20588 12656
rect 20444 12300 20496 12306
rect 20444 12242 20496 12248
rect 20548 12170 20576 12650
rect 20536 12164 20588 12170
rect 20536 12106 20588 12112
rect 20996 12096 21048 12102
rect 20996 12038 21048 12044
rect 20352 11892 20404 11898
rect 20352 11834 20404 11840
rect 19524 11824 19576 11830
rect 19524 11766 19576 11772
rect 19708 11824 19760 11830
rect 19708 11766 19760 11772
rect 19340 11552 19392 11558
rect 19340 11494 19392 11500
rect 19432 11552 19484 11558
rect 19432 11494 19484 11500
rect 19444 11218 19472 11494
rect 19536 11354 19564 11766
rect 19524 11348 19576 11354
rect 19524 11290 19576 11296
rect 19432 11212 19484 11218
rect 19432 11154 19484 11160
rect 19720 11150 19748 11766
rect 21008 11354 21036 12038
rect 20996 11348 21048 11354
rect 20996 11290 21048 11296
rect 19708 11144 19760 11150
rect 19708 11086 19760 11092
rect 21008 11082 21036 11290
rect 21100 11150 21128 12786
rect 21192 12238 21220 12922
rect 21284 12238 21312 20742
rect 21652 19718 21680 39238
rect 22756 38214 22784 39374
rect 23492 39098 23520 39918
rect 24596 39438 24624 40394
rect 24584 39432 24636 39438
rect 24584 39374 24636 39380
rect 23480 39092 23532 39098
rect 23480 39034 23532 39040
rect 22928 38956 22980 38962
rect 22928 38898 22980 38904
rect 22744 38208 22796 38214
rect 22744 38150 22796 38156
rect 21824 37868 21876 37874
rect 21824 37810 21876 37816
rect 21916 37868 21968 37874
rect 21916 37810 21968 37816
rect 21732 36576 21784 36582
rect 21732 36518 21784 36524
rect 21744 36242 21772 36518
rect 21732 36236 21784 36242
rect 21732 36178 21784 36184
rect 21836 35154 21864 37810
rect 21928 36378 21956 37810
rect 22468 37120 22520 37126
rect 22468 37062 22520 37068
rect 22480 36854 22508 37062
rect 22468 36848 22520 36854
rect 22468 36790 22520 36796
rect 22100 36780 22152 36786
rect 22100 36722 22152 36728
rect 22652 36780 22704 36786
rect 22652 36722 22704 36728
rect 21916 36372 21968 36378
rect 21916 36314 21968 36320
rect 21824 35148 21876 35154
rect 21824 35090 21876 35096
rect 22112 34626 22140 36722
rect 22664 36106 22692 36722
rect 22836 36576 22888 36582
rect 22836 36518 22888 36524
rect 22652 36100 22704 36106
rect 22652 36042 22704 36048
rect 22664 35630 22692 36042
rect 22284 35624 22336 35630
rect 22284 35566 22336 35572
rect 22652 35624 22704 35630
rect 22652 35566 22704 35572
rect 22192 35012 22244 35018
rect 22192 34954 22244 34960
rect 22204 34746 22232 34954
rect 22192 34740 22244 34746
rect 22192 34682 22244 34688
rect 22112 34598 22232 34626
rect 22204 33930 22232 34598
rect 22192 33924 22244 33930
rect 22192 33866 22244 33872
rect 22204 33590 22232 33866
rect 22192 33584 22244 33590
rect 22192 33526 22244 33532
rect 22100 31748 22152 31754
rect 22100 31690 22152 31696
rect 22008 31680 22060 31686
rect 22008 31622 22060 31628
rect 22020 31346 22048 31622
rect 22112 31482 22140 31690
rect 22100 31476 22152 31482
rect 22100 31418 22152 31424
rect 22008 31340 22060 31346
rect 22008 31282 22060 31288
rect 22204 30258 22232 33526
rect 22192 30252 22244 30258
rect 22192 30194 22244 30200
rect 22296 30054 22324 35566
rect 22560 35556 22612 35562
rect 22560 35498 22612 35504
rect 22376 35488 22428 35494
rect 22376 35430 22428 35436
rect 22388 34610 22416 35430
rect 22572 34610 22600 35498
rect 22664 35306 22692 35566
rect 22848 35562 22876 36518
rect 22836 35556 22888 35562
rect 22836 35498 22888 35504
rect 22664 35290 22784 35306
rect 22664 35284 22796 35290
rect 22664 35278 22744 35284
rect 22744 35226 22796 35232
rect 22652 35080 22704 35086
rect 22652 35022 22704 35028
rect 22376 34604 22428 34610
rect 22376 34546 22428 34552
rect 22560 34604 22612 34610
rect 22560 34546 22612 34552
rect 22664 33998 22692 35022
rect 22756 34610 22784 35226
rect 22940 34678 22968 38898
rect 24964 38350 24992 40870
rect 26436 40662 26464 43200
rect 26700 40928 26752 40934
rect 26700 40870 26752 40876
rect 26976 40928 27028 40934
rect 26976 40870 27028 40876
rect 26424 40656 26476 40662
rect 26424 40598 26476 40604
rect 26712 40594 26740 40870
rect 26700 40588 26752 40594
rect 26700 40530 26752 40536
rect 26332 40452 26384 40458
rect 26332 40394 26384 40400
rect 26344 40050 26372 40394
rect 26988 40050 27016 40870
rect 25964 40044 26016 40050
rect 25964 39986 26016 39992
rect 26332 40044 26384 40050
rect 26332 39986 26384 39992
rect 26976 40044 27028 40050
rect 26976 39986 27028 39992
rect 25976 39098 26004 39986
rect 27356 39982 27384 43302
rect 27710 43200 27766 44000
rect 28354 43200 28410 44000
rect 29642 43330 29698 44000
rect 29642 43302 30052 43330
rect 29642 43200 29698 43302
rect 29552 40928 29604 40934
rect 29552 40870 29604 40876
rect 29564 40594 29592 40870
rect 30024 40594 30052 43302
rect 30286 43200 30342 44000
rect 30930 43200 30986 44000
rect 32218 43330 32274 44000
rect 32218 43302 32444 43330
rect 32218 43200 32274 43302
rect 32128 40928 32180 40934
rect 32128 40870 32180 40876
rect 32312 40928 32364 40934
rect 32312 40870 32364 40876
rect 29552 40588 29604 40594
rect 29552 40530 29604 40536
rect 30012 40588 30064 40594
rect 30012 40530 30064 40536
rect 29736 40452 29788 40458
rect 29736 40394 29788 40400
rect 29748 40186 29776 40394
rect 29736 40180 29788 40186
rect 29736 40122 29788 40128
rect 32140 40050 32168 40870
rect 32324 40594 32352 40870
rect 32312 40588 32364 40594
rect 32312 40530 32364 40536
rect 29276 40044 29328 40050
rect 29276 39986 29328 39992
rect 31392 40044 31444 40050
rect 31392 39986 31444 39992
rect 32128 40044 32180 40050
rect 32128 39986 32180 39992
rect 27160 39976 27212 39982
rect 27160 39918 27212 39924
rect 27344 39976 27396 39982
rect 27344 39918 27396 39924
rect 27172 39642 27200 39918
rect 27160 39636 27212 39642
rect 27160 39578 27212 39584
rect 26608 39432 26660 39438
rect 26608 39374 26660 39380
rect 25964 39092 26016 39098
rect 25964 39034 26016 39040
rect 26620 38865 26648 39374
rect 29288 39302 29316 39986
rect 31404 39370 31432 39986
rect 32416 39982 32444 43302
rect 32862 43200 32918 44000
rect 33506 43200 33562 44000
rect 34150 43200 34206 44000
rect 35438 43200 35494 44000
rect 36082 43200 36138 44000
rect 36726 43200 36782 44000
rect 37370 43200 37426 44000
rect 38658 43200 38714 44000
rect 39302 43200 39358 44000
rect 39946 43200 40002 44000
rect 40590 43330 40646 44000
rect 40420 43302 40646 43330
rect 32876 40594 32904 43200
rect 34164 41002 34192 43200
rect 34520 41200 34572 41206
rect 34520 41142 34572 41148
rect 34152 40996 34204 41002
rect 34152 40938 34204 40944
rect 32864 40588 32916 40594
rect 32864 40530 32916 40536
rect 32496 40452 32548 40458
rect 32496 40394 32548 40400
rect 32404 39976 32456 39982
rect 32404 39918 32456 39924
rect 32508 39642 32536 40394
rect 34532 39642 34560 41142
rect 34934 40828 35242 40848
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40752 35242 40772
rect 36096 40594 36124 43200
rect 36084 40588 36136 40594
rect 36084 40530 36136 40536
rect 35900 40452 35952 40458
rect 35900 40394 35952 40400
rect 34796 40112 34848 40118
rect 34796 40054 34848 40060
rect 34808 39642 34836 40054
rect 35348 39976 35400 39982
rect 35348 39918 35400 39924
rect 34934 39740 35242 39760
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39664 35242 39684
rect 32496 39636 32548 39642
rect 32496 39578 32548 39584
rect 34520 39636 34572 39642
rect 34520 39578 34572 39584
rect 34796 39636 34848 39642
rect 34796 39578 34848 39584
rect 32862 39536 32918 39545
rect 32862 39471 32918 39480
rect 32876 39438 32904 39471
rect 32864 39432 32916 39438
rect 32864 39374 32916 39380
rect 31392 39364 31444 39370
rect 31392 39306 31444 39312
rect 29276 39296 29328 39302
rect 29276 39238 29328 39244
rect 29288 39001 29316 39238
rect 29274 38992 29330 39001
rect 35360 38962 35388 39918
rect 35912 39642 35940 40394
rect 35900 39636 35952 39642
rect 35900 39578 35952 39584
rect 36740 39574 36768 43200
rect 39302 41576 39358 41585
rect 39302 41511 39358 41520
rect 37464 40928 37516 40934
rect 37464 40870 37516 40876
rect 37476 40594 37504 40870
rect 39316 40594 39344 41511
rect 40132 40996 40184 41002
rect 40132 40938 40184 40944
rect 40040 40928 40092 40934
rect 40040 40870 40092 40876
rect 37464 40588 37516 40594
rect 37464 40530 37516 40536
rect 39304 40588 39356 40594
rect 39304 40530 39356 40536
rect 37004 40520 37056 40526
rect 37004 40462 37056 40468
rect 37016 39642 37044 40462
rect 37648 40452 37700 40458
rect 37648 40394 37700 40400
rect 37660 40186 37688 40394
rect 39302 40216 39358 40225
rect 37648 40180 37700 40186
rect 39302 40151 39358 40160
rect 37648 40122 37700 40128
rect 39316 40118 39344 40151
rect 39304 40112 39356 40118
rect 39304 40054 39356 40060
rect 40052 40050 40080 40870
rect 38200 40044 38252 40050
rect 38200 39986 38252 39992
rect 40040 40044 40092 40050
rect 40040 39986 40092 39992
rect 37004 39636 37056 39642
rect 37004 39578 37056 39584
rect 36728 39568 36780 39574
rect 36728 39510 36780 39516
rect 35900 39432 35952 39438
rect 35900 39374 35952 39380
rect 29274 38927 29330 38936
rect 32680 38956 32732 38962
rect 32680 38898 32732 38904
rect 32864 38956 32916 38962
rect 32864 38898 32916 38904
rect 33508 38956 33560 38962
rect 33508 38898 33560 38904
rect 35348 38956 35400 38962
rect 35348 38898 35400 38904
rect 26606 38856 26662 38865
rect 26606 38791 26662 38800
rect 25964 38412 26016 38418
rect 25964 38354 26016 38360
rect 24952 38344 25004 38350
rect 24952 38286 25004 38292
rect 25872 38344 25924 38350
rect 25872 38286 25924 38292
rect 23388 38208 23440 38214
rect 23388 38150 23440 38156
rect 24768 38208 24820 38214
rect 24768 38150 24820 38156
rect 23296 37664 23348 37670
rect 23296 37606 23348 37612
rect 23308 37262 23336 37606
rect 23204 37256 23256 37262
rect 23124 37204 23204 37210
rect 23124 37198 23256 37204
rect 23296 37256 23348 37262
rect 23296 37198 23348 37204
rect 23124 37182 23244 37198
rect 23124 36786 23152 37182
rect 23204 37120 23256 37126
rect 23204 37062 23256 37068
rect 23216 36922 23244 37062
rect 23204 36916 23256 36922
rect 23204 36858 23256 36864
rect 23112 36780 23164 36786
rect 23112 36722 23164 36728
rect 23308 36718 23336 37198
rect 23296 36712 23348 36718
rect 23296 36654 23348 36660
rect 23308 36174 23336 36654
rect 23296 36168 23348 36174
rect 23296 36110 23348 36116
rect 23400 35086 23428 38150
rect 23848 37868 23900 37874
rect 23848 37810 23900 37816
rect 24124 37868 24176 37874
rect 24124 37810 24176 37816
rect 23860 36854 23888 37810
rect 23848 36848 23900 36854
rect 23848 36790 23900 36796
rect 23480 36576 23532 36582
rect 23480 36518 23532 36524
rect 23492 35698 23520 36518
rect 23860 36378 23888 36790
rect 24136 36718 24164 37810
rect 24308 37664 24360 37670
rect 24308 37606 24360 37612
rect 24320 37330 24348 37606
rect 24308 37324 24360 37330
rect 24308 37266 24360 37272
rect 24124 36712 24176 36718
rect 24124 36654 24176 36660
rect 23848 36372 23900 36378
rect 23848 36314 23900 36320
rect 24136 35834 24164 36654
rect 24320 36242 24348 37266
rect 24780 36378 24808 38150
rect 24964 38010 24992 38286
rect 25228 38276 25280 38282
rect 25228 38218 25280 38224
rect 24952 38004 25004 38010
rect 24952 37946 25004 37952
rect 24860 37120 24912 37126
rect 24860 37062 24912 37068
rect 24872 36378 24900 37062
rect 24768 36372 24820 36378
rect 24768 36314 24820 36320
rect 24860 36372 24912 36378
rect 24860 36314 24912 36320
rect 24308 36236 24360 36242
rect 24308 36178 24360 36184
rect 24124 35828 24176 35834
rect 24124 35770 24176 35776
rect 24964 35766 24992 37946
rect 25136 37868 25188 37874
rect 25136 37810 25188 37816
rect 25148 37466 25176 37810
rect 25136 37460 25188 37466
rect 25136 37402 25188 37408
rect 25136 37188 25188 37194
rect 25136 37130 25188 37136
rect 25148 35766 25176 37130
rect 25240 36922 25268 38218
rect 25320 37256 25372 37262
rect 25320 37198 25372 37204
rect 25332 36922 25360 37198
rect 25884 37194 25912 38286
rect 25976 37670 26004 38354
rect 26056 38344 26108 38350
rect 26056 38286 26108 38292
rect 25964 37664 26016 37670
rect 25964 37606 26016 37612
rect 25976 37262 26004 37606
rect 25964 37256 26016 37262
rect 25964 37198 26016 37204
rect 25872 37188 25924 37194
rect 25872 37130 25924 37136
rect 25228 36916 25280 36922
rect 25228 36858 25280 36864
rect 25320 36916 25372 36922
rect 25320 36858 25372 36864
rect 25240 36718 25268 36858
rect 25320 36780 25372 36786
rect 25320 36722 25372 36728
rect 25228 36712 25280 36718
rect 25228 36654 25280 36660
rect 25332 36564 25360 36722
rect 25688 36712 25740 36718
rect 25688 36654 25740 36660
rect 25596 36576 25648 36582
rect 25332 36536 25596 36564
rect 25596 36518 25648 36524
rect 25320 36168 25372 36174
rect 25320 36110 25372 36116
rect 24952 35760 25004 35766
rect 24952 35702 25004 35708
rect 25136 35760 25188 35766
rect 25136 35702 25188 35708
rect 23480 35692 23532 35698
rect 23480 35634 23532 35640
rect 24400 35692 24452 35698
rect 24400 35634 24452 35640
rect 24768 35692 24820 35698
rect 24768 35634 24820 35640
rect 23756 35624 23808 35630
rect 23756 35566 23808 35572
rect 23388 35080 23440 35086
rect 23388 35022 23440 35028
rect 22928 34672 22980 34678
rect 22928 34614 22980 34620
rect 22744 34604 22796 34610
rect 22940 34586 23152 34614
rect 22744 34546 22796 34552
rect 22928 34536 22980 34542
rect 22928 34478 22980 34484
rect 22652 33992 22704 33998
rect 22652 33934 22704 33940
rect 22664 33318 22692 33934
rect 22652 33312 22704 33318
rect 22652 33254 22704 33260
rect 22560 32904 22612 32910
rect 22664 32858 22692 33254
rect 22612 32852 22692 32858
rect 22560 32846 22692 32852
rect 22572 32830 22692 32846
rect 22560 32496 22612 32502
rect 22560 32438 22612 32444
rect 22468 32020 22520 32026
rect 22468 31962 22520 31968
rect 22480 30410 22508 31962
rect 22572 30938 22600 32438
rect 22664 31822 22692 32830
rect 22652 31816 22704 31822
rect 22652 31758 22704 31764
rect 22560 30932 22612 30938
rect 22560 30874 22612 30880
rect 22652 30660 22704 30666
rect 22652 30602 22704 30608
rect 22480 30382 22600 30410
rect 22468 30252 22520 30258
rect 22468 30194 22520 30200
rect 22284 30048 22336 30054
rect 22284 29990 22336 29996
rect 22296 29102 22324 29990
rect 22480 29850 22508 30194
rect 22468 29844 22520 29850
rect 22468 29786 22520 29792
rect 22376 29776 22428 29782
rect 22376 29718 22428 29724
rect 22284 29096 22336 29102
rect 22284 29038 22336 29044
rect 22388 29034 22416 29718
rect 22376 29028 22428 29034
rect 22376 28970 22428 28976
rect 21732 28756 21784 28762
rect 21732 28698 21784 28704
rect 21744 28150 21772 28698
rect 22480 28626 22508 29786
rect 22572 29034 22600 30382
rect 22560 29028 22612 29034
rect 22560 28970 22612 28976
rect 22572 28694 22600 28970
rect 22664 28762 22692 30602
rect 22940 29850 22968 34478
rect 23020 33516 23072 33522
rect 23020 33458 23072 33464
rect 23032 32502 23060 33458
rect 23020 32496 23072 32502
rect 23020 32438 23072 32444
rect 22928 29844 22980 29850
rect 22928 29786 22980 29792
rect 22652 28756 22704 28762
rect 22652 28698 22704 28704
rect 22560 28688 22612 28694
rect 22560 28630 22612 28636
rect 22468 28620 22520 28626
rect 22468 28562 22520 28568
rect 22376 28552 22428 28558
rect 22376 28494 22428 28500
rect 21732 28144 21784 28150
rect 21732 28086 21784 28092
rect 22388 27606 22416 28494
rect 22376 27600 22428 27606
rect 22376 27542 22428 27548
rect 21732 27328 21784 27334
rect 21732 27270 21784 27276
rect 22560 27328 22612 27334
rect 22560 27270 22612 27276
rect 21744 26382 21772 27270
rect 21916 26988 21968 26994
rect 21916 26930 21968 26936
rect 21928 26586 21956 26930
rect 21916 26580 21968 26586
rect 21916 26522 21968 26528
rect 22572 26518 22600 27270
rect 22560 26512 22612 26518
rect 22560 26454 22612 26460
rect 23020 26512 23072 26518
rect 23020 26454 23072 26460
rect 21732 26376 21784 26382
rect 21732 26318 21784 26324
rect 21744 25702 21772 26318
rect 23032 25906 23060 26454
rect 23020 25900 23072 25906
rect 23020 25842 23072 25848
rect 21732 25696 21784 25702
rect 21732 25638 21784 25644
rect 22008 24812 22060 24818
rect 22008 24754 22060 24760
rect 22020 24138 22048 24754
rect 22468 24744 22520 24750
rect 22468 24686 22520 24692
rect 22376 24200 22428 24206
rect 22376 24142 22428 24148
rect 22008 24132 22060 24138
rect 22008 24074 22060 24080
rect 22020 23662 22048 24074
rect 22388 23866 22416 24142
rect 22376 23860 22428 23866
rect 22376 23802 22428 23808
rect 22480 23662 22508 24686
rect 22560 24608 22612 24614
rect 22560 24550 22612 24556
rect 22572 24206 22600 24550
rect 22560 24200 22612 24206
rect 22560 24142 22612 24148
rect 22008 23656 22060 23662
rect 22008 23598 22060 23604
rect 22468 23656 22520 23662
rect 22468 23598 22520 23604
rect 21916 23520 21968 23526
rect 21916 23462 21968 23468
rect 21928 22250 21956 23462
rect 22020 23254 22048 23598
rect 22008 23248 22060 23254
rect 22008 23190 22060 23196
rect 22744 22568 22796 22574
rect 22744 22510 22796 22516
rect 21744 22234 21956 22250
rect 22756 22234 22784 22510
rect 21732 22228 21956 22234
rect 21784 22222 21956 22228
rect 21732 22170 21784 22176
rect 21824 21956 21876 21962
rect 21824 21898 21876 21904
rect 21836 21418 21864 21898
rect 21928 21622 21956 22222
rect 22744 22228 22796 22234
rect 22744 22170 22796 22176
rect 22008 22024 22060 22030
rect 22008 21966 22060 21972
rect 21916 21616 21968 21622
rect 21916 21558 21968 21564
rect 21824 21412 21876 21418
rect 21824 21354 21876 21360
rect 21824 21072 21876 21078
rect 21824 21014 21876 21020
rect 21836 20806 21864 21014
rect 21824 20800 21876 20806
rect 21824 20742 21876 20748
rect 21640 19712 21692 19718
rect 21640 19654 21692 19660
rect 21640 18216 21692 18222
rect 21640 18158 21692 18164
rect 21364 17196 21416 17202
rect 21364 17138 21416 17144
rect 21376 16794 21404 17138
rect 21364 16788 21416 16794
rect 21364 16730 21416 16736
rect 21364 15496 21416 15502
rect 21364 15438 21416 15444
rect 21376 13938 21404 15438
rect 21364 13932 21416 13938
rect 21364 13874 21416 13880
rect 21548 13320 21600 13326
rect 21548 13262 21600 13268
rect 21560 12986 21588 13262
rect 21548 12980 21600 12986
rect 21548 12922 21600 12928
rect 21180 12232 21232 12238
rect 21180 12174 21232 12180
rect 21272 12232 21324 12238
rect 21272 12174 21324 12180
rect 21652 12102 21680 18158
rect 21732 16448 21784 16454
rect 21732 16390 21784 16396
rect 21744 15638 21772 16390
rect 21836 15910 21864 20742
rect 22020 19786 22048 21966
rect 22928 21888 22980 21894
rect 22928 21830 22980 21836
rect 22940 21690 22968 21830
rect 22928 21684 22980 21690
rect 22928 21626 22980 21632
rect 22008 19780 22060 19786
rect 22008 19722 22060 19728
rect 22744 19780 22796 19786
rect 22744 19722 22796 19728
rect 22020 19378 22048 19722
rect 22008 19372 22060 19378
rect 22008 19314 22060 19320
rect 22468 19372 22520 19378
rect 22468 19314 22520 19320
rect 22020 18766 22048 19314
rect 22008 18760 22060 18766
rect 22008 18702 22060 18708
rect 22284 18760 22336 18766
rect 22284 18702 22336 18708
rect 22296 18426 22324 18702
rect 22284 18420 22336 18426
rect 22284 18362 22336 18368
rect 22100 17128 22152 17134
rect 22100 17070 22152 17076
rect 22112 16114 22140 17070
rect 22192 16992 22244 16998
rect 22192 16934 22244 16940
rect 22204 16658 22232 16934
rect 22192 16652 22244 16658
rect 22192 16594 22244 16600
rect 22100 16108 22152 16114
rect 22100 16050 22152 16056
rect 21824 15904 21876 15910
rect 21824 15846 21876 15852
rect 21732 15632 21784 15638
rect 21732 15574 21784 15580
rect 21744 14346 21772 15574
rect 21836 15502 21864 15846
rect 21824 15496 21876 15502
rect 21824 15438 21876 15444
rect 21732 14340 21784 14346
rect 21732 14282 21784 14288
rect 22112 14006 22140 16050
rect 22480 15706 22508 19314
rect 22756 18902 22784 19722
rect 22744 18896 22796 18902
rect 22744 18838 22796 18844
rect 22468 15700 22520 15706
rect 22468 15642 22520 15648
rect 22652 15428 22704 15434
rect 22652 15370 22704 15376
rect 22284 14884 22336 14890
rect 22284 14826 22336 14832
rect 22192 14612 22244 14618
rect 22192 14554 22244 14560
rect 22100 14000 22152 14006
rect 22100 13942 22152 13948
rect 22204 12646 22232 14554
rect 22296 14006 22324 14826
rect 22664 14822 22692 15370
rect 22744 15088 22796 15094
rect 22744 15030 22796 15036
rect 22376 14816 22428 14822
rect 22376 14758 22428 14764
rect 22652 14816 22704 14822
rect 22652 14758 22704 14764
rect 22284 14000 22336 14006
rect 22284 13942 22336 13948
rect 22388 13326 22416 14758
rect 22468 13932 22520 13938
rect 22468 13874 22520 13880
rect 22480 13394 22508 13874
rect 22664 13530 22692 14758
rect 22756 14618 22784 15030
rect 22744 14612 22796 14618
rect 22744 14554 22796 14560
rect 23124 14006 23152 34586
rect 23768 34542 23796 35566
rect 23940 35488 23992 35494
rect 23940 35430 23992 35436
rect 23756 34536 23808 34542
rect 23756 34478 23808 34484
rect 23664 33312 23716 33318
rect 23664 33254 23716 33260
rect 23676 32910 23704 33254
rect 23664 32904 23716 32910
rect 23664 32846 23716 32852
rect 23768 32722 23796 34478
rect 23848 33516 23900 33522
rect 23848 33458 23900 33464
rect 23676 32694 23796 32722
rect 23388 31340 23440 31346
rect 23388 31282 23440 31288
rect 23572 31340 23624 31346
rect 23572 31282 23624 31288
rect 23296 31136 23348 31142
rect 23296 31078 23348 31084
rect 23308 30938 23336 31078
rect 23296 30932 23348 30938
rect 23296 30874 23348 30880
rect 23400 30190 23428 31282
rect 23584 30734 23612 31282
rect 23572 30728 23624 30734
rect 23572 30670 23624 30676
rect 23584 30394 23612 30670
rect 23572 30388 23624 30394
rect 23572 30330 23624 30336
rect 23388 30184 23440 30190
rect 23388 30126 23440 30132
rect 23400 29782 23428 30126
rect 23388 29776 23440 29782
rect 23388 29718 23440 29724
rect 23400 29238 23428 29718
rect 23388 29232 23440 29238
rect 23388 29174 23440 29180
rect 23676 28694 23704 32694
rect 23860 32570 23888 33458
rect 23848 32564 23900 32570
rect 23848 32506 23900 32512
rect 23952 32434 23980 35430
rect 24412 34542 24440 35634
rect 24780 35290 24808 35634
rect 24768 35284 24820 35290
rect 24768 35226 24820 35232
rect 24964 35222 24992 35702
rect 25228 35692 25280 35698
rect 25228 35634 25280 35640
rect 24952 35216 25004 35222
rect 25004 35164 25084 35170
rect 24952 35158 25084 35164
rect 24964 35142 25084 35158
rect 24952 35080 25004 35086
rect 24952 35022 25004 35028
rect 24400 34536 24452 34542
rect 24400 34478 24452 34484
rect 24860 33448 24912 33454
rect 24860 33390 24912 33396
rect 24768 33312 24820 33318
rect 24768 33254 24820 33260
rect 24780 32910 24808 33254
rect 24872 33114 24900 33390
rect 24860 33108 24912 33114
rect 24860 33050 24912 33056
rect 24872 32910 24900 33050
rect 24768 32904 24820 32910
rect 24768 32846 24820 32852
rect 24860 32904 24912 32910
rect 24860 32846 24912 32852
rect 24400 32768 24452 32774
rect 24400 32710 24452 32716
rect 24412 32502 24440 32710
rect 24400 32496 24452 32502
rect 24400 32438 24452 32444
rect 23940 32428 23992 32434
rect 23940 32370 23992 32376
rect 24216 32428 24268 32434
rect 24216 32370 24268 32376
rect 23756 32360 23808 32366
rect 23756 32302 23808 32308
rect 23664 28688 23716 28694
rect 23664 28630 23716 28636
rect 23676 28490 23704 28630
rect 23664 28484 23716 28490
rect 23664 28426 23716 28432
rect 23664 28008 23716 28014
rect 23664 27950 23716 27956
rect 23296 27532 23348 27538
rect 23296 27474 23348 27480
rect 23204 27464 23256 27470
rect 23204 27406 23256 27412
rect 23216 27130 23244 27406
rect 23308 27130 23336 27474
rect 23204 27124 23256 27130
rect 23204 27066 23256 27072
rect 23296 27124 23348 27130
rect 23296 27066 23348 27072
rect 23216 26450 23244 27066
rect 23572 27056 23624 27062
rect 23676 27010 23704 27950
rect 23624 27004 23704 27010
rect 23572 26998 23704 27004
rect 23584 26982 23704 26998
rect 23676 26450 23704 26982
rect 23204 26444 23256 26450
rect 23204 26386 23256 26392
rect 23664 26444 23716 26450
rect 23664 26386 23716 26392
rect 23676 25906 23704 26386
rect 23664 25900 23716 25906
rect 23664 25842 23716 25848
rect 23296 25696 23348 25702
rect 23296 25638 23348 25644
rect 23204 24608 23256 24614
rect 23204 24550 23256 24556
rect 23216 23798 23244 24550
rect 23204 23792 23256 23798
rect 23204 23734 23256 23740
rect 23308 23118 23336 25638
rect 23480 25152 23532 25158
rect 23480 25094 23532 25100
rect 23388 24812 23440 24818
rect 23388 24754 23440 24760
rect 23400 24410 23428 24754
rect 23388 24404 23440 24410
rect 23388 24346 23440 24352
rect 23388 23180 23440 23186
rect 23388 23122 23440 23128
rect 23296 23112 23348 23118
rect 23296 23054 23348 23060
rect 23400 22506 23428 23122
rect 23388 22500 23440 22506
rect 23388 22442 23440 22448
rect 23400 22166 23428 22442
rect 23388 22160 23440 22166
rect 23388 22102 23440 22108
rect 23492 21554 23520 25094
rect 23768 24274 23796 32302
rect 24228 31346 24256 32370
rect 24780 32366 24808 32846
rect 24768 32360 24820 32366
rect 24768 32302 24820 32308
rect 24872 32026 24900 32846
rect 24964 32570 24992 35022
rect 25056 34678 25084 35142
rect 25044 34672 25096 34678
rect 25044 34614 25096 34620
rect 25136 34604 25188 34610
rect 25136 34546 25188 34552
rect 25148 33522 25176 34546
rect 25240 34474 25268 35634
rect 25228 34468 25280 34474
rect 25228 34410 25280 34416
rect 25332 34354 25360 36110
rect 25504 35828 25556 35834
rect 25504 35770 25556 35776
rect 25412 34536 25464 34542
rect 25412 34478 25464 34484
rect 25240 34326 25360 34354
rect 25044 33516 25096 33522
rect 25044 33458 25096 33464
rect 25136 33516 25188 33522
rect 25136 33458 25188 33464
rect 25056 33046 25084 33458
rect 25044 33040 25096 33046
rect 25044 32982 25096 32988
rect 25056 32910 25084 32982
rect 25044 32904 25096 32910
rect 25044 32846 25096 32852
rect 24952 32564 25004 32570
rect 24952 32506 25004 32512
rect 24964 32434 24992 32506
rect 24952 32428 25004 32434
rect 24952 32370 25004 32376
rect 24860 32020 24912 32026
rect 24860 31962 24912 31968
rect 24676 31816 24728 31822
rect 24676 31758 24728 31764
rect 24768 31816 24820 31822
rect 24768 31758 24820 31764
rect 24216 31340 24268 31346
rect 24216 31282 24268 31288
rect 23848 29572 23900 29578
rect 23848 29514 23900 29520
rect 23860 28558 23888 29514
rect 23848 28552 23900 28558
rect 23848 28494 23900 28500
rect 23860 27062 23888 28494
rect 23848 27056 23900 27062
rect 23900 27004 24072 27010
rect 23848 26998 24072 27004
rect 23860 26982 24072 26998
rect 24044 26976 24072 26982
rect 24044 26948 24164 26976
rect 23848 26376 23900 26382
rect 23848 26318 23900 26324
rect 23756 24268 23808 24274
rect 23756 24210 23808 24216
rect 23860 23730 23888 26318
rect 24032 24268 24084 24274
rect 24032 24210 24084 24216
rect 23848 23724 23900 23730
rect 23848 23666 23900 23672
rect 23848 23112 23900 23118
rect 23848 23054 23900 23060
rect 23860 22642 23888 23054
rect 23848 22636 23900 22642
rect 23848 22578 23900 22584
rect 23480 21548 23532 21554
rect 23480 21490 23532 21496
rect 23492 20942 23520 21490
rect 23480 20936 23532 20942
rect 23480 20878 23532 20884
rect 23492 14822 23520 20878
rect 23940 20460 23992 20466
rect 23940 20402 23992 20408
rect 23952 19786 23980 20402
rect 23940 19780 23992 19786
rect 23940 19722 23992 19728
rect 23572 18692 23624 18698
rect 23572 18634 23624 18640
rect 23480 14816 23532 14822
rect 23480 14758 23532 14764
rect 23112 14000 23164 14006
rect 23112 13942 23164 13948
rect 22652 13524 22704 13530
rect 22652 13466 22704 13472
rect 22468 13388 22520 13394
rect 22468 13330 22520 13336
rect 22376 13320 22428 13326
rect 22376 13262 22428 13268
rect 22192 12640 22244 12646
rect 22192 12582 22244 12588
rect 21640 12096 21692 12102
rect 21640 12038 21692 12044
rect 22480 11762 22508 13330
rect 23492 12434 23520 14758
rect 23584 14550 23612 18634
rect 23664 17536 23716 17542
rect 23664 17478 23716 17484
rect 23848 17536 23900 17542
rect 23848 17478 23900 17484
rect 23676 16590 23704 17478
rect 23860 16794 23888 17478
rect 23848 16788 23900 16794
rect 23848 16730 23900 16736
rect 23664 16584 23716 16590
rect 23664 16526 23716 16532
rect 23676 16114 23704 16526
rect 23756 16516 23808 16522
rect 23756 16458 23808 16464
rect 23664 16108 23716 16114
rect 23664 16050 23716 16056
rect 23768 15978 23796 16458
rect 23756 15972 23808 15978
rect 23756 15914 23808 15920
rect 23572 14544 23624 14550
rect 23572 14486 23624 14492
rect 23940 12844 23992 12850
rect 23940 12786 23992 12792
rect 23400 12406 23520 12434
rect 21180 11756 21232 11762
rect 21180 11698 21232 11704
rect 22468 11756 22520 11762
rect 22468 11698 22520 11704
rect 22560 11756 22612 11762
rect 22560 11698 22612 11704
rect 21192 11354 21220 11698
rect 21180 11348 21232 11354
rect 21180 11290 21232 11296
rect 21088 11144 21140 11150
rect 21088 11086 21140 11092
rect 22192 11144 22244 11150
rect 22192 11086 22244 11092
rect 20996 11076 21048 11082
rect 20996 11018 21048 11024
rect 19248 11008 19300 11014
rect 19248 10950 19300 10956
rect 19432 11008 19484 11014
rect 19432 10950 19484 10956
rect 18696 10804 18748 10810
rect 18696 10746 18748 10752
rect 18512 10668 18564 10674
rect 18512 10610 18564 10616
rect 18236 10532 18288 10538
rect 18236 10474 18288 10480
rect 18708 10266 18736 10746
rect 19260 10742 19288 10950
rect 19248 10736 19300 10742
rect 19248 10678 19300 10684
rect 19444 10674 19472 10950
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 21100 10810 21128 11086
rect 21088 10804 21140 10810
rect 21088 10746 21140 10752
rect 19064 10668 19116 10674
rect 19064 10610 19116 10616
rect 19432 10668 19484 10674
rect 19432 10610 19484 10616
rect 19984 10668 20036 10674
rect 19984 10610 20036 10616
rect 18236 10260 18288 10266
rect 18236 10202 18288 10208
rect 18696 10260 18748 10266
rect 18696 10202 18748 10208
rect 18248 9926 18276 10202
rect 19076 10130 19104 10610
rect 19156 10600 19208 10606
rect 19156 10542 19208 10548
rect 19064 10124 19116 10130
rect 19064 10066 19116 10072
rect 18236 9920 18288 9926
rect 18236 9862 18288 9868
rect 18144 9716 18196 9722
rect 18144 9658 18196 9664
rect 18144 9512 18196 9518
rect 18248 9500 18276 9862
rect 18788 9648 18840 9654
rect 18788 9590 18840 9596
rect 18196 9472 18276 9500
rect 18512 9512 18564 9518
rect 18144 9454 18196 9460
rect 18696 9512 18748 9518
rect 18564 9472 18696 9500
rect 18512 9454 18564 9460
rect 18696 9454 18748 9460
rect 18800 9450 18828 9590
rect 18788 9444 18840 9450
rect 18788 9386 18840 9392
rect 18052 8968 18104 8974
rect 18052 8910 18104 8916
rect 17868 8492 17920 8498
rect 17868 8434 17920 8440
rect 17132 8424 17184 8430
rect 17132 8366 17184 8372
rect 17408 8424 17460 8430
rect 17408 8366 17460 8372
rect 17224 8288 17276 8294
rect 17224 8230 17276 8236
rect 16856 7948 16908 7954
rect 16856 7890 16908 7896
rect 16120 7880 16172 7886
rect 16120 7822 16172 7828
rect 17132 7812 17184 7818
rect 17132 7754 17184 7760
rect 17144 7274 17172 7754
rect 17236 7478 17264 8230
rect 17224 7472 17276 7478
rect 17224 7414 17276 7420
rect 17420 7410 17448 8366
rect 17880 8090 17908 8434
rect 19168 8294 19196 10542
rect 19248 10464 19300 10470
rect 19248 10406 19300 10412
rect 19260 10062 19288 10406
rect 19248 10056 19300 10062
rect 19248 9998 19300 10004
rect 19444 9994 19472 10610
rect 19996 10266 20024 10610
rect 19984 10260 20036 10266
rect 19984 10202 20036 10208
rect 22204 10062 22232 11086
rect 22192 10056 22244 10062
rect 22192 9998 22244 10004
rect 22376 10056 22428 10062
rect 22376 9998 22428 10004
rect 19432 9988 19484 9994
rect 19432 9930 19484 9936
rect 21732 9920 21784 9926
rect 21732 9862 21784 9868
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 21744 9586 21772 9862
rect 21732 9580 21784 9586
rect 21732 9522 21784 9528
rect 22192 9580 22244 9586
rect 22192 9522 22244 9528
rect 21548 9172 21600 9178
rect 21548 9114 21600 9120
rect 21560 8974 21588 9114
rect 21744 9042 21772 9522
rect 21732 9036 21784 9042
rect 21732 8978 21784 8984
rect 20996 8968 21048 8974
rect 20996 8910 21048 8916
rect 21548 8968 21600 8974
rect 21548 8910 21600 8916
rect 20720 8900 20772 8906
rect 20720 8842 20772 8848
rect 19432 8832 19484 8838
rect 19432 8774 19484 8780
rect 20628 8832 20680 8838
rect 20628 8774 20680 8780
rect 19444 8566 19472 8774
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 19432 8560 19484 8566
rect 19432 8502 19484 8508
rect 20260 8356 20312 8362
rect 20260 8298 20312 8304
rect 18604 8288 18656 8294
rect 18604 8230 18656 8236
rect 19156 8288 19208 8294
rect 19156 8230 19208 8236
rect 17868 8084 17920 8090
rect 17868 8026 17920 8032
rect 17880 7546 17908 8026
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 18616 7410 18644 8230
rect 18788 7812 18840 7818
rect 18788 7754 18840 7760
rect 18800 7546 18828 7754
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 18788 7540 18840 7546
rect 18788 7482 18840 7488
rect 17408 7404 17460 7410
rect 17408 7346 17460 7352
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 17132 7268 17184 7274
rect 17132 7210 17184 7216
rect 20272 6798 20300 8298
rect 20640 8090 20668 8774
rect 20732 8498 20760 8842
rect 21008 8498 21036 8910
rect 21560 8634 21588 8910
rect 21548 8628 21600 8634
rect 21548 8570 21600 8576
rect 21744 8498 21772 8978
rect 22204 8634 22232 9522
rect 22388 9178 22416 9998
rect 22480 9518 22508 11698
rect 22572 10266 22600 11698
rect 22836 11348 22888 11354
rect 22836 11290 22888 11296
rect 22848 10606 22876 11290
rect 23400 11150 23428 12406
rect 23952 11898 23980 12786
rect 23940 11892 23992 11898
rect 23940 11834 23992 11840
rect 23480 11756 23532 11762
rect 23480 11698 23532 11704
rect 23388 11144 23440 11150
rect 23388 11086 23440 11092
rect 22836 10600 22888 10606
rect 22836 10542 22888 10548
rect 23492 10266 23520 11698
rect 24044 11354 24072 24210
rect 24136 21690 24164 26948
rect 24228 23050 24256 31282
rect 24400 30592 24452 30598
rect 24400 30534 24452 30540
rect 24412 30326 24440 30534
rect 24400 30320 24452 30326
rect 24400 30262 24452 30268
rect 24688 30258 24716 31758
rect 24780 31346 24808 31758
rect 25044 31476 25096 31482
rect 25044 31418 25096 31424
rect 24768 31340 24820 31346
rect 24768 31282 24820 31288
rect 24860 31136 24912 31142
rect 24860 31078 24912 31084
rect 24872 30734 24900 31078
rect 25056 30938 25084 31418
rect 25044 30932 25096 30938
rect 25044 30874 25096 30880
rect 25056 30734 25084 30874
rect 25148 30870 25176 33458
rect 25136 30864 25188 30870
rect 25136 30806 25188 30812
rect 24872 30728 24938 30734
rect 24872 30688 24886 30728
rect 24886 30670 24938 30676
rect 25044 30728 25096 30734
rect 25044 30670 25096 30676
rect 24676 30252 24728 30258
rect 24676 30194 24728 30200
rect 25136 29708 25188 29714
rect 25136 29650 25188 29656
rect 25148 29578 25176 29650
rect 25136 29572 25188 29578
rect 25136 29514 25188 29520
rect 24952 29504 25004 29510
rect 24952 29446 25004 29452
rect 24860 29232 24912 29238
rect 24860 29174 24912 29180
rect 24584 29028 24636 29034
rect 24584 28970 24636 28976
rect 24308 28960 24360 28966
rect 24308 28902 24360 28908
rect 24320 25906 24348 28902
rect 24400 28076 24452 28082
rect 24400 28018 24452 28024
rect 24412 27674 24440 28018
rect 24400 27668 24452 27674
rect 24400 27610 24452 27616
rect 24492 27600 24544 27606
rect 24492 27542 24544 27548
rect 24400 26240 24452 26246
rect 24400 26182 24452 26188
rect 24412 25974 24440 26182
rect 24400 25968 24452 25974
rect 24400 25910 24452 25916
rect 24308 25900 24360 25906
rect 24308 25842 24360 25848
rect 24320 25362 24348 25842
rect 24308 25356 24360 25362
rect 24308 25298 24360 25304
rect 24504 25242 24532 27542
rect 24596 27470 24624 28970
rect 24872 28694 24900 29174
rect 24860 28688 24912 28694
rect 24860 28630 24912 28636
rect 24584 27464 24636 27470
rect 24584 27406 24636 27412
rect 24584 26376 24636 26382
rect 24584 26318 24636 26324
rect 24596 25498 24624 26318
rect 24964 26042 24992 29446
rect 25148 27606 25176 29514
rect 25240 29510 25268 34326
rect 25424 32910 25452 34478
rect 25412 32904 25464 32910
rect 25412 32846 25464 32852
rect 25516 32230 25544 35770
rect 25608 35086 25636 36518
rect 25700 36174 25728 36654
rect 25884 36242 25912 37130
rect 25976 36938 26004 37198
rect 26068 37126 26096 38286
rect 26424 38208 26476 38214
rect 26424 38150 26476 38156
rect 26332 37936 26384 37942
rect 26332 37878 26384 37884
rect 26344 37262 26372 37878
rect 26332 37256 26384 37262
rect 26332 37198 26384 37204
rect 26056 37120 26108 37126
rect 26056 37062 26108 37068
rect 25976 36910 26096 36938
rect 25872 36236 25924 36242
rect 25792 36196 25872 36224
rect 25688 36168 25740 36174
rect 25688 36110 25740 36116
rect 25688 36032 25740 36038
rect 25688 35974 25740 35980
rect 25700 35290 25728 35974
rect 25792 35494 25820 36196
rect 25872 36178 25924 36184
rect 26068 36174 26096 36910
rect 26436 36174 26464 38150
rect 26620 37670 26648 38791
rect 30656 38548 30708 38554
rect 30656 38490 30708 38496
rect 30196 38344 30248 38350
rect 30196 38286 30248 38292
rect 30104 38208 30156 38214
rect 30104 38150 30156 38156
rect 28448 37936 28500 37942
rect 28448 37878 28500 37884
rect 28264 37868 28316 37874
rect 28264 37810 28316 37816
rect 26608 37664 26660 37670
rect 26608 37606 26660 37612
rect 26608 37188 26660 37194
rect 26608 37130 26660 37136
rect 26620 36378 26648 37130
rect 28276 36922 28304 37810
rect 28264 36916 28316 36922
rect 28264 36858 28316 36864
rect 26884 36780 26936 36786
rect 26884 36722 26936 36728
rect 26608 36372 26660 36378
rect 26608 36314 26660 36320
rect 26056 36168 26108 36174
rect 26056 36110 26108 36116
rect 26424 36168 26476 36174
rect 26424 36110 26476 36116
rect 25872 35760 25924 35766
rect 25872 35702 25924 35708
rect 25780 35488 25832 35494
rect 25780 35430 25832 35436
rect 25688 35284 25740 35290
rect 25688 35226 25740 35232
rect 25792 35154 25820 35430
rect 25780 35148 25832 35154
rect 25780 35090 25832 35096
rect 25884 35086 25912 35702
rect 26068 35630 26096 36110
rect 25964 35624 26016 35630
rect 25964 35566 26016 35572
rect 26056 35624 26108 35630
rect 26056 35566 26108 35572
rect 25976 35086 26004 35566
rect 26608 35556 26660 35562
rect 26608 35498 26660 35504
rect 26148 35488 26200 35494
rect 26148 35430 26200 35436
rect 26160 35086 26188 35430
rect 26620 35086 26648 35498
rect 25596 35080 25648 35086
rect 25596 35022 25648 35028
rect 25872 35080 25924 35086
rect 25872 35022 25924 35028
rect 25964 35080 26016 35086
rect 25964 35022 26016 35028
rect 26148 35080 26200 35086
rect 26148 35022 26200 35028
rect 26608 35080 26660 35086
rect 26608 35022 26660 35028
rect 25688 34944 25740 34950
rect 25688 34886 25740 34892
rect 25700 34610 25728 34886
rect 25688 34604 25740 34610
rect 25688 34546 25740 34552
rect 25976 33658 26004 35022
rect 26896 35018 26924 36722
rect 28460 35698 28488 37878
rect 30116 37874 30144 38150
rect 30104 37868 30156 37874
rect 30104 37810 30156 37816
rect 30208 37466 30236 38286
rect 30288 38276 30340 38282
rect 30288 38218 30340 38224
rect 30300 38010 30328 38218
rect 30288 38004 30340 38010
rect 30288 37946 30340 37952
rect 29736 37460 29788 37466
rect 29736 37402 29788 37408
rect 30196 37460 30248 37466
rect 30196 37402 30248 37408
rect 29748 37194 29776 37402
rect 29920 37392 29972 37398
rect 29920 37334 29972 37340
rect 29000 37188 29052 37194
rect 29000 37130 29052 37136
rect 29736 37188 29788 37194
rect 29736 37130 29788 37136
rect 28632 37120 28684 37126
rect 28632 37062 28684 37068
rect 28908 37120 28960 37126
rect 28908 37062 28960 37068
rect 28644 36786 28672 37062
rect 28920 36922 28948 37062
rect 28908 36916 28960 36922
rect 28908 36858 28960 36864
rect 28632 36780 28684 36786
rect 28632 36722 28684 36728
rect 26976 35692 27028 35698
rect 26976 35634 27028 35640
rect 28448 35692 28500 35698
rect 28448 35634 28500 35640
rect 26988 35018 27016 35634
rect 28460 35154 28488 35634
rect 28448 35148 28500 35154
rect 28448 35090 28500 35096
rect 28908 35148 28960 35154
rect 28908 35090 28960 35096
rect 26424 35012 26476 35018
rect 26424 34954 26476 34960
rect 26516 35012 26568 35018
rect 26516 34954 26568 34960
rect 26884 35012 26936 35018
rect 26884 34954 26936 34960
rect 26976 35012 27028 35018
rect 26976 34954 27028 34960
rect 26436 34610 26464 34954
rect 26424 34604 26476 34610
rect 26424 34546 26476 34552
rect 26528 34406 26556 34954
rect 26516 34400 26568 34406
rect 26516 34342 26568 34348
rect 26528 33998 26556 34342
rect 26148 33992 26200 33998
rect 26148 33934 26200 33940
rect 26516 33992 26568 33998
rect 26516 33934 26568 33940
rect 25964 33652 26016 33658
rect 25964 33594 26016 33600
rect 26160 33454 26188 33934
rect 26528 33522 26556 33934
rect 26516 33516 26568 33522
rect 26516 33458 26568 33464
rect 26148 33448 26200 33454
rect 26148 33390 26200 33396
rect 25688 33312 25740 33318
rect 25688 33254 25740 33260
rect 26332 33312 26384 33318
rect 26332 33254 26384 33260
rect 25700 32978 25728 33254
rect 26148 33108 26200 33114
rect 26148 33050 26200 33056
rect 25688 32972 25740 32978
rect 25688 32914 25740 32920
rect 26160 32910 26188 33050
rect 26148 32904 26200 32910
rect 26148 32846 26200 32852
rect 26240 32836 26292 32842
rect 26240 32778 26292 32784
rect 25320 32224 25372 32230
rect 25320 32166 25372 32172
rect 25504 32224 25556 32230
rect 25504 32166 25556 32172
rect 25872 32224 25924 32230
rect 25872 32166 25924 32172
rect 25228 29504 25280 29510
rect 25228 29446 25280 29452
rect 25136 27600 25188 27606
rect 25136 27542 25188 27548
rect 25044 27464 25096 27470
rect 25044 27406 25096 27412
rect 25056 26382 25084 27406
rect 25044 26376 25096 26382
rect 25044 26318 25096 26324
rect 24952 26036 25004 26042
rect 24952 25978 25004 25984
rect 24584 25492 24636 25498
rect 24584 25434 24636 25440
rect 24320 25214 24532 25242
rect 24216 23044 24268 23050
rect 24216 22986 24268 22992
rect 24216 22024 24268 22030
rect 24216 21966 24268 21972
rect 24124 21684 24176 21690
rect 24124 21626 24176 21632
rect 24228 20602 24256 21966
rect 24216 20596 24268 20602
rect 24320 20584 24348 25214
rect 25056 24682 25084 26318
rect 25136 25696 25188 25702
rect 25136 25638 25188 25644
rect 25148 25430 25176 25638
rect 25136 25424 25188 25430
rect 25136 25366 25188 25372
rect 25332 24750 25360 32166
rect 25504 31884 25556 31890
rect 25504 31826 25556 31832
rect 25516 30394 25544 31826
rect 25688 31408 25740 31414
rect 25688 31350 25740 31356
rect 25504 30388 25556 30394
rect 25504 30330 25556 30336
rect 25516 29510 25544 30330
rect 25700 30258 25728 31350
rect 25884 31346 25912 32166
rect 25964 31816 26016 31822
rect 25964 31758 26016 31764
rect 25976 31686 26004 31758
rect 25964 31680 26016 31686
rect 25964 31622 26016 31628
rect 25976 31482 26004 31622
rect 26252 31482 26280 32778
rect 26344 32774 26372 33254
rect 26332 32768 26384 32774
rect 26332 32710 26384 32716
rect 25964 31476 26016 31482
rect 25964 31418 26016 31424
rect 26240 31476 26292 31482
rect 26240 31418 26292 31424
rect 25872 31340 25924 31346
rect 25872 31282 25924 31288
rect 25884 31226 25912 31282
rect 25792 31198 26004 31226
rect 25792 30938 25820 31198
rect 25976 31142 26004 31198
rect 25872 31136 25924 31142
rect 25872 31078 25924 31084
rect 25964 31136 26016 31142
rect 25964 31078 26016 31084
rect 25780 30932 25832 30938
rect 25780 30874 25832 30880
rect 25792 30326 25820 30874
rect 25780 30320 25832 30326
rect 25780 30262 25832 30268
rect 25688 30252 25740 30258
rect 25688 30194 25740 30200
rect 25884 29850 25912 31078
rect 26252 30666 26280 31418
rect 26344 31278 26372 32710
rect 26988 32570 27016 34954
rect 27252 34944 27304 34950
rect 27252 34886 27304 34892
rect 27264 34678 27292 34886
rect 27252 34672 27304 34678
rect 27252 34614 27304 34620
rect 27528 34604 27580 34610
rect 27528 34546 27580 34552
rect 27160 34196 27212 34202
rect 27160 34138 27212 34144
rect 27068 33652 27120 33658
rect 27068 33594 27120 33600
rect 27080 32910 27108 33594
rect 27172 33114 27200 34138
rect 27540 33658 27568 34546
rect 28448 33924 28500 33930
rect 28448 33866 28500 33872
rect 27988 33856 28040 33862
rect 27988 33798 28040 33804
rect 27528 33652 27580 33658
rect 27528 33594 27580 33600
rect 28000 33590 28028 33798
rect 27988 33584 28040 33590
rect 27988 33526 28040 33532
rect 27160 33108 27212 33114
rect 27160 33050 27212 33056
rect 27068 32904 27120 32910
rect 27068 32846 27120 32852
rect 26424 32564 26476 32570
rect 26424 32506 26476 32512
rect 26976 32564 27028 32570
rect 26976 32506 27028 32512
rect 26436 31822 26464 32506
rect 27080 32366 27108 32846
rect 27160 32428 27212 32434
rect 27160 32370 27212 32376
rect 27068 32360 27120 32366
rect 27068 32302 27120 32308
rect 27172 32026 27200 32370
rect 27160 32020 27212 32026
rect 27160 31962 27212 31968
rect 26424 31816 26476 31822
rect 26424 31758 26476 31764
rect 27172 31754 27200 31962
rect 26976 31748 27028 31754
rect 27172 31726 27384 31754
rect 26976 31690 27028 31696
rect 26988 31482 27016 31690
rect 26976 31476 27028 31482
rect 26976 31418 27028 31424
rect 27356 31414 27384 31726
rect 28460 31414 28488 33866
rect 28920 33522 28948 35090
rect 29012 33930 29040 37130
rect 29748 36922 29776 37130
rect 29736 36916 29788 36922
rect 29736 36858 29788 36864
rect 29736 36168 29788 36174
rect 29736 36110 29788 36116
rect 29552 36032 29604 36038
rect 29552 35974 29604 35980
rect 29564 35766 29592 35974
rect 29748 35834 29776 36110
rect 29736 35828 29788 35834
rect 29736 35770 29788 35776
rect 29552 35760 29604 35766
rect 29552 35702 29604 35708
rect 29828 35012 29880 35018
rect 29828 34954 29880 34960
rect 29840 34202 29868 34954
rect 29932 34610 29960 37334
rect 30300 37126 30328 37946
rect 30668 37262 30696 38490
rect 32692 38486 32720 38898
rect 32680 38480 32732 38486
rect 32680 38422 32732 38428
rect 31668 38276 31720 38282
rect 31668 38218 31720 38224
rect 31208 38208 31260 38214
rect 31208 38150 31260 38156
rect 31220 38010 31248 38150
rect 31208 38004 31260 38010
rect 31208 37946 31260 37952
rect 30656 37256 30708 37262
rect 30656 37198 30708 37204
rect 30288 37120 30340 37126
rect 30288 37062 30340 37068
rect 30300 36786 30328 37062
rect 30668 36922 30696 37198
rect 30656 36916 30708 36922
rect 30656 36858 30708 36864
rect 31220 36786 31248 37946
rect 31300 37664 31352 37670
rect 31300 37606 31352 37612
rect 31312 37466 31340 37606
rect 31680 37466 31708 38218
rect 32128 38208 32180 38214
rect 32128 38150 32180 38156
rect 31300 37460 31352 37466
rect 31300 37402 31352 37408
rect 31668 37460 31720 37466
rect 31668 37402 31720 37408
rect 31680 37262 31708 37402
rect 31668 37256 31720 37262
rect 31668 37198 31720 37204
rect 31760 37188 31812 37194
rect 31760 37130 31812 37136
rect 30288 36780 30340 36786
rect 30288 36722 30340 36728
rect 31208 36780 31260 36786
rect 31208 36722 31260 36728
rect 30656 36168 30708 36174
rect 30656 36110 30708 36116
rect 30748 36168 30800 36174
rect 30748 36110 30800 36116
rect 30668 35562 30696 36110
rect 30656 35556 30708 35562
rect 30656 35498 30708 35504
rect 30564 35284 30616 35290
rect 30564 35226 30616 35232
rect 30576 34746 30604 35226
rect 30288 34740 30340 34746
rect 30288 34682 30340 34688
rect 30564 34740 30616 34746
rect 30564 34682 30616 34688
rect 29920 34604 29972 34610
rect 29920 34546 29972 34552
rect 29828 34196 29880 34202
rect 29828 34138 29880 34144
rect 29000 33924 29052 33930
rect 29000 33866 29052 33872
rect 28908 33516 28960 33522
rect 28908 33458 28960 33464
rect 28920 32434 28948 33458
rect 29932 33114 29960 34546
rect 30012 34400 30064 34406
rect 30012 34342 30064 34348
rect 30024 33998 30052 34342
rect 30300 34066 30328 34682
rect 30668 34610 30696 35498
rect 30760 35290 30788 36110
rect 31772 36038 31800 37130
rect 32140 36786 32168 38150
rect 32692 37874 32720 38422
rect 32876 38350 32904 38898
rect 33324 38752 33376 38758
rect 33324 38694 33376 38700
rect 32864 38344 32916 38350
rect 32864 38286 32916 38292
rect 32772 37936 32824 37942
rect 32772 37878 32824 37884
rect 32680 37868 32732 37874
rect 32680 37810 32732 37816
rect 32220 37120 32272 37126
rect 32220 37062 32272 37068
rect 32784 37074 32812 37878
rect 32876 37670 32904 38286
rect 32864 37664 32916 37670
rect 32864 37606 32916 37612
rect 32876 37262 32904 37606
rect 33336 37466 33364 38694
rect 33520 38010 33548 38898
rect 33784 38752 33836 38758
rect 33784 38694 33836 38700
rect 33796 38350 33824 38694
rect 34934 38652 35242 38672
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38576 35242 38596
rect 33784 38344 33836 38350
rect 33784 38286 33836 38292
rect 34796 38344 34848 38350
rect 34796 38286 34848 38292
rect 33508 38004 33560 38010
rect 33508 37946 33560 37952
rect 34520 37868 34572 37874
rect 34520 37810 34572 37816
rect 33324 37460 33376 37466
rect 33324 37402 33376 37408
rect 32864 37256 32916 37262
rect 32864 37198 32916 37204
rect 32956 37256 33008 37262
rect 32956 37198 33008 37204
rect 32864 37120 32916 37126
rect 32784 37068 32864 37074
rect 32784 37062 32916 37068
rect 32128 36780 32180 36786
rect 32128 36722 32180 36728
rect 31760 36032 31812 36038
rect 31760 35974 31812 35980
rect 32140 35834 32168 36722
rect 32128 35828 32180 35834
rect 32128 35770 32180 35776
rect 30840 35760 30892 35766
rect 30840 35702 30892 35708
rect 30748 35284 30800 35290
rect 30748 35226 30800 35232
rect 30852 34746 30880 35702
rect 32036 35692 32088 35698
rect 32036 35634 32088 35640
rect 31392 35556 31444 35562
rect 31392 35498 31444 35504
rect 30932 35488 30984 35494
rect 30932 35430 30984 35436
rect 30840 34740 30892 34746
rect 30840 34682 30892 34688
rect 30380 34604 30432 34610
rect 30380 34546 30432 34552
rect 30656 34604 30708 34610
rect 30656 34546 30708 34552
rect 30392 34202 30420 34546
rect 30380 34196 30432 34202
rect 30380 34138 30432 34144
rect 30288 34060 30340 34066
rect 30288 34002 30340 34008
rect 30012 33992 30064 33998
rect 30012 33934 30064 33940
rect 29920 33108 29972 33114
rect 29920 33050 29972 33056
rect 30944 33046 30972 35430
rect 31208 35284 31260 35290
rect 31208 35226 31260 35232
rect 31220 34746 31248 35226
rect 31208 34740 31260 34746
rect 31208 34682 31260 34688
rect 30932 33040 30984 33046
rect 30932 32982 30984 32988
rect 29920 32904 29972 32910
rect 29920 32846 29972 32852
rect 29932 32570 29960 32846
rect 30944 32570 30972 32982
rect 31208 32768 31260 32774
rect 31208 32710 31260 32716
rect 29920 32564 29972 32570
rect 29920 32506 29972 32512
rect 30932 32564 30984 32570
rect 30932 32506 30984 32512
rect 28632 32428 28684 32434
rect 28632 32370 28684 32376
rect 28908 32428 28960 32434
rect 28908 32370 28960 32376
rect 29644 32428 29696 32434
rect 29644 32370 29696 32376
rect 31116 32428 31168 32434
rect 31116 32370 31168 32376
rect 28540 31884 28592 31890
rect 28540 31826 28592 31832
rect 27344 31408 27396 31414
rect 27344 31350 27396 31356
rect 28448 31408 28500 31414
rect 28448 31350 28500 31356
rect 26332 31272 26384 31278
rect 26332 31214 26384 31220
rect 27160 31272 27212 31278
rect 27160 31214 27212 31220
rect 26884 31204 26936 31210
rect 26884 31146 26936 31152
rect 26896 30938 26924 31146
rect 26884 30932 26936 30938
rect 26884 30874 26936 30880
rect 27068 30728 27120 30734
rect 27068 30670 27120 30676
rect 26240 30660 26292 30666
rect 26240 30602 26292 30608
rect 26252 30394 26280 30602
rect 26240 30388 26292 30394
rect 26240 30330 26292 30336
rect 27080 29850 27108 30670
rect 27172 30258 27200 31214
rect 28552 30802 28580 31826
rect 28540 30796 28592 30802
rect 28540 30738 28592 30744
rect 28448 30660 28500 30666
rect 28448 30602 28500 30608
rect 27160 30252 27212 30258
rect 27160 30194 27212 30200
rect 27804 30252 27856 30258
rect 27804 30194 27856 30200
rect 27816 29850 27844 30194
rect 25872 29844 25924 29850
rect 25872 29786 25924 29792
rect 27068 29844 27120 29850
rect 27068 29786 27120 29792
rect 27804 29844 27856 29850
rect 27804 29786 27856 29792
rect 28460 29714 28488 30602
rect 28552 30258 28580 30738
rect 28644 30666 28672 32370
rect 28920 31890 28948 32370
rect 28908 31884 28960 31890
rect 28908 31826 28960 31832
rect 29184 31680 29236 31686
rect 29184 31622 29236 31628
rect 29000 31340 29052 31346
rect 29000 31282 29052 31288
rect 29012 30870 29040 31282
rect 29000 30864 29052 30870
rect 29000 30806 29052 30812
rect 28632 30660 28684 30666
rect 28632 30602 28684 30608
rect 28540 30252 28592 30258
rect 28540 30194 28592 30200
rect 28632 30048 28684 30054
rect 28552 29996 28632 30002
rect 28552 29990 28684 29996
rect 28552 29974 28672 29990
rect 28448 29708 28500 29714
rect 28448 29650 28500 29656
rect 25780 29572 25832 29578
rect 25780 29514 25832 29520
rect 25504 29504 25556 29510
rect 25504 29446 25556 29452
rect 25792 29238 25820 29514
rect 26608 29300 26660 29306
rect 26608 29242 26660 29248
rect 25780 29232 25832 29238
rect 25780 29174 25832 29180
rect 25964 29232 26016 29238
rect 25964 29174 26016 29180
rect 25976 28626 26004 29174
rect 26332 28960 26384 28966
rect 26332 28902 26384 28908
rect 25964 28620 26016 28626
rect 25964 28562 26016 28568
rect 25688 28416 25740 28422
rect 25688 28358 25740 28364
rect 25872 28416 25924 28422
rect 25872 28358 25924 28364
rect 25596 26988 25648 26994
rect 25596 26930 25648 26936
rect 25608 26586 25636 26930
rect 25596 26580 25648 26586
rect 25596 26522 25648 26528
rect 25412 26240 25464 26246
rect 25412 26182 25464 26188
rect 25424 26042 25452 26182
rect 25412 26036 25464 26042
rect 25412 25978 25464 25984
rect 25504 25900 25556 25906
rect 25504 25842 25556 25848
rect 25516 25498 25544 25842
rect 25504 25492 25556 25498
rect 25504 25434 25556 25440
rect 25700 25294 25728 28358
rect 25884 28150 25912 28358
rect 25872 28144 25924 28150
rect 25872 28086 25924 28092
rect 25780 28076 25832 28082
rect 25780 28018 25832 28024
rect 25792 27470 25820 28018
rect 25976 27674 26004 28562
rect 26240 28552 26292 28558
rect 26240 28494 26292 28500
rect 26056 28144 26108 28150
rect 26056 28086 26108 28092
rect 25964 27668 26016 27674
rect 25964 27610 26016 27616
rect 26068 27470 26096 28086
rect 26252 27878 26280 28494
rect 26344 28218 26372 28902
rect 26332 28212 26384 28218
rect 26332 28154 26384 28160
rect 26240 27872 26292 27878
rect 26240 27814 26292 27820
rect 25780 27464 25832 27470
rect 25780 27406 25832 27412
rect 26056 27464 26108 27470
rect 26056 27406 26108 27412
rect 26332 26784 26384 26790
rect 26332 26726 26384 26732
rect 26344 26382 26372 26726
rect 26332 26376 26384 26382
rect 26332 26318 26384 26324
rect 26332 25900 26384 25906
rect 26332 25842 26384 25848
rect 26240 25764 26292 25770
rect 26240 25706 26292 25712
rect 26252 25362 26280 25706
rect 26240 25356 26292 25362
rect 26240 25298 26292 25304
rect 25688 25288 25740 25294
rect 25688 25230 25740 25236
rect 25700 24954 25728 25230
rect 25688 24948 25740 24954
rect 25688 24890 25740 24896
rect 25320 24744 25372 24750
rect 25320 24686 25372 24692
rect 25044 24676 25096 24682
rect 25044 24618 25096 24624
rect 25596 24268 25648 24274
rect 25596 24210 25648 24216
rect 24400 24200 24452 24206
rect 24400 24142 24452 24148
rect 24492 24200 24544 24206
rect 24492 24142 24544 24148
rect 24412 23866 24440 24142
rect 24400 23860 24452 23866
rect 24400 23802 24452 23808
rect 24412 23186 24440 23802
rect 24400 23180 24452 23186
rect 24400 23122 24452 23128
rect 24504 23118 24532 24142
rect 24676 24064 24728 24070
rect 24676 24006 24728 24012
rect 24688 23798 24716 24006
rect 25608 23866 25636 24210
rect 25700 24206 25728 24890
rect 26252 24614 26280 25298
rect 26240 24608 26292 24614
rect 26240 24550 26292 24556
rect 26252 24206 26280 24550
rect 26344 24342 26372 25842
rect 26620 25362 26648 29242
rect 28552 29170 28580 29974
rect 29012 29714 29040 30806
rect 29000 29708 29052 29714
rect 29000 29650 29052 29656
rect 29000 29504 29052 29510
rect 29000 29446 29052 29452
rect 28356 29164 28408 29170
rect 28356 29106 28408 29112
rect 28540 29164 28592 29170
rect 28540 29106 28592 29112
rect 27160 28960 27212 28966
rect 27160 28902 27212 28908
rect 26884 28756 26936 28762
rect 26884 28698 26936 28704
rect 26700 27328 26752 27334
rect 26700 27270 26752 27276
rect 26608 25356 26660 25362
rect 26608 25298 26660 25304
rect 26620 24750 26648 25298
rect 26712 24954 26740 27270
rect 26700 24948 26752 24954
rect 26700 24890 26752 24896
rect 26608 24744 26660 24750
rect 26608 24686 26660 24692
rect 26332 24336 26384 24342
rect 26332 24278 26384 24284
rect 25688 24200 25740 24206
rect 25688 24142 25740 24148
rect 26240 24200 26292 24206
rect 26240 24142 26292 24148
rect 25596 23860 25648 23866
rect 25596 23802 25648 23808
rect 24676 23792 24728 23798
rect 24676 23734 24728 23740
rect 25136 23724 25188 23730
rect 25136 23666 25188 23672
rect 24860 23656 24912 23662
rect 24860 23598 24912 23604
rect 24872 23322 24900 23598
rect 24860 23316 24912 23322
rect 24860 23258 24912 23264
rect 24492 23112 24544 23118
rect 24492 23054 24544 23060
rect 24400 23044 24452 23050
rect 24400 22986 24452 22992
rect 24412 21690 24440 22986
rect 24504 22234 24532 23054
rect 25148 22574 25176 23666
rect 26240 23316 26292 23322
rect 26240 23258 26292 23264
rect 25136 22568 25188 22574
rect 25136 22510 25188 22516
rect 24492 22228 24544 22234
rect 24492 22170 24544 22176
rect 25148 22166 25176 22510
rect 25136 22160 25188 22166
rect 25136 22102 25188 22108
rect 26056 22024 26108 22030
rect 26056 21966 26108 21972
rect 25964 21956 26016 21962
rect 25964 21898 26016 21904
rect 24400 21684 24452 21690
rect 24400 21626 24452 21632
rect 24400 21548 24452 21554
rect 24400 21490 24452 21496
rect 24676 21548 24728 21554
rect 24676 21490 24728 21496
rect 24412 21146 24440 21490
rect 24584 21412 24636 21418
rect 24584 21354 24636 21360
rect 24400 21140 24452 21146
rect 24400 21082 24452 21088
rect 24596 20942 24624 21354
rect 24688 21350 24716 21490
rect 24768 21480 24820 21486
rect 24768 21422 24820 21428
rect 24676 21344 24728 21350
rect 24676 21286 24728 21292
rect 24584 20936 24636 20942
rect 24584 20878 24636 20884
rect 24320 20556 24440 20584
rect 24216 20538 24268 20544
rect 24124 20460 24176 20466
rect 24124 20402 24176 20408
rect 24308 20460 24360 20466
rect 24308 20402 24360 20408
rect 24136 19990 24164 20402
rect 24124 19984 24176 19990
rect 24124 19926 24176 19932
rect 24320 19514 24348 20402
rect 24308 19508 24360 19514
rect 24308 19450 24360 19456
rect 24308 19236 24360 19242
rect 24308 19178 24360 19184
rect 24320 13954 24348 19178
rect 24412 15094 24440 20556
rect 24596 19854 24624 20878
rect 24584 19848 24636 19854
rect 24584 19790 24636 19796
rect 24596 19718 24624 19790
rect 24584 19712 24636 19718
rect 24584 19654 24636 19660
rect 24492 19372 24544 19378
rect 24492 19314 24544 19320
rect 24504 18630 24532 19314
rect 24596 19310 24624 19654
rect 24584 19304 24636 19310
rect 24584 19246 24636 19252
rect 24688 19242 24716 21286
rect 24780 20602 24808 21422
rect 25136 21344 25188 21350
rect 25136 21286 25188 21292
rect 25148 21146 25176 21286
rect 25136 21140 25188 21146
rect 25136 21082 25188 21088
rect 25044 20936 25096 20942
rect 25044 20878 25096 20884
rect 24860 20868 24912 20874
rect 24860 20810 24912 20816
rect 24768 20596 24820 20602
rect 24768 20538 24820 20544
rect 24872 20466 24900 20810
rect 25056 20534 25084 20878
rect 25044 20528 25096 20534
rect 24964 20488 25044 20516
rect 24860 20460 24912 20466
rect 24860 20402 24912 20408
rect 24860 20324 24912 20330
rect 24860 20266 24912 20272
rect 24768 19848 24820 19854
rect 24768 19790 24820 19796
rect 24780 19378 24808 19790
rect 24768 19372 24820 19378
rect 24768 19314 24820 19320
rect 24676 19236 24728 19242
rect 24676 19178 24728 19184
rect 24872 19174 24900 20266
rect 24964 19854 24992 20488
rect 25044 20470 25096 20476
rect 24952 19848 25004 19854
rect 24952 19790 25004 19796
rect 24964 19514 24992 19790
rect 24952 19508 25004 19514
rect 24952 19450 25004 19456
rect 24860 19168 24912 19174
rect 24860 19110 24912 19116
rect 24492 18624 24544 18630
rect 24492 18566 24544 18572
rect 24768 17196 24820 17202
rect 24768 17138 24820 17144
rect 24492 16992 24544 16998
rect 24492 16934 24544 16940
rect 24504 16658 24532 16934
rect 24780 16794 24808 17138
rect 24768 16788 24820 16794
rect 24768 16730 24820 16736
rect 24492 16652 24544 16658
rect 24492 16594 24544 16600
rect 24504 16114 24532 16594
rect 24780 16538 24808 16730
rect 24860 16652 24912 16658
rect 24860 16594 24912 16600
rect 24596 16522 24808 16538
rect 24596 16516 24820 16522
rect 24596 16510 24768 16516
rect 24492 16108 24544 16114
rect 24492 16050 24544 16056
rect 24596 15910 24624 16510
rect 24768 16458 24820 16464
rect 24676 16448 24728 16454
rect 24676 16390 24728 16396
rect 24688 16114 24716 16390
rect 24676 16108 24728 16114
rect 24676 16050 24728 16056
rect 24584 15904 24636 15910
rect 24584 15846 24636 15852
rect 24400 15088 24452 15094
rect 24400 15030 24452 15036
rect 24412 14074 24440 15030
rect 24688 14822 24716 16050
rect 24780 15978 24808 16458
rect 24768 15972 24820 15978
rect 24768 15914 24820 15920
rect 24872 15910 24900 16594
rect 25148 16454 25176 21082
rect 25976 21010 26004 21898
rect 26068 21690 26096 21966
rect 26056 21684 26108 21690
rect 26056 21626 26108 21632
rect 25964 21004 26016 21010
rect 25964 20946 26016 20952
rect 25780 20324 25832 20330
rect 25780 20266 25832 20272
rect 25228 20256 25280 20262
rect 25228 20198 25280 20204
rect 25240 19854 25268 20198
rect 25792 19922 25820 20266
rect 25504 19916 25556 19922
rect 25504 19858 25556 19864
rect 25780 19916 25832 19922
rect 25780 19858 25832 19864
rect 25228 19848 25280 19854
rect 25228 19790 25280 19796
rect 25240 19514 25268 19790
rect 25228 19508 25280 19514
rect 25228 19450 25280 19456
rect 25516 19378 25544 19858
rect 25504 19372 25556 19378
rect 25504 19314 25556 19320
rect 25516 18902 25544 19314
rect 26252 18970 26280 23258
rect 26344 23254 26372 24278
rect 26712 23730 26740 24890
rect 26700 23724 26752 23730
rect 26700 23666 26752 23672
rect 26896 23322 26924 28698
rect 27172 28558 27200 28902
rect 28368 28558 28396 29106
rect 27160 28552 27212 28558
rect 27160 28494 27212 28500
rect 27896 28552 27948 28558
rect 27896 28494 27948 28500
rect 28356 28552 28408 28558
rect 28356 28494 28408 28500
rect 27908 28218 27936 28494
rect 27896 28212 27948 28218
rect 27896 28154 27948 28160
rect 27436 27872 27488 27878
rect 27436 27814 27488 27820
rect 27160 25696 27212 25702
rect 27160 25638 27212 25644
rect 27172 25362 27200 25638
rect 27160 25356 27212 25362
rect 27160 25298 27212 25304
rect 27160 24812 27212 24818
rect 27160 24754 27212 24760
rect 27172 24274 27200 24754
rect 27448 24682 27476 27814
rect 27804 27464 27856 27470
rect 27804 27406 27856 27412
rect 27816 27130 27844 27406
rect 27908 27402 27936 28154
rect 28172 27872 28224 27878
rect 28172 27814 28224 27820
rect 28184 27674 28212 27814
rect 28172 27668 28224 27674
rect 28172 27610 28224 27616
rect 27896 27396 27948 27402
rect 27896 27338 27948 27344
rect 27908 27130 27936 27338
rect 27804 27124 27856 27130
rect 27804 27066 27856 27072
rect 27896 27124 27948 27130
rect 27896 27066 27948 27072
rect 27528 26240 27580 26246
rect 27528 26182 27580 26188
rect 27540 25974 27568 26182
rect 27528 25968 27580 25974
rect 27528 25910 27580 25916
rect 27540 24886 27568 25910
rect 27816 25226 27844 27066
rect 27908 25906 27936 27066
rect 28368 26994 28396 28494
rect 28448 28212 28500 28218
rect 28448 28154 28500 28160
rect 28460 28082 28488 28154
rect 28448 28076 28500 28082
rect 28448 28018 28500 28024
rect 28552 27554 28580 29106
rect 28816 28688 28868 28694
rect 28816 28630 28868 28636
rect 28632 28552 28684 28558
rect 28632 28494 28684 28500
rect 28644 27878 28672 28494
rect 28828 27946 28856 28630
rect 29012 28422 29040 29446
rect 29196 29170 29224 31622
rect 29656 31482 29684 32370
rect 30380 32292 30432 32298
rect 30380 32234 30432 32240
rect 29644 31476 29696 31482
rect 29644 31418 29696 31424
rect 30392 31414 30420 32234
rect 31128 32230 31156 32370
rect 31220 32366 31248 32710
rect 31208 32360 31260 32366
rect 31208 32302 31260 32308
rect 31404 32298 31432 35498
rect 32048 35086 32076 35634
rect 32036 35080 32088 35086
rect 32036 35022 32088 35028
rect 31852 34944 31904 34950
rect 31852 34886 31904 34892
rect 31864 34406 31892 34886
rect 32048 34474 32076 35022
rect 32036 34468 32088 34474
rect 32036 34410 32088 34416
rect 31852 34400 31904 34406
rect 31852 34342 31904 34348
rect 32048 34202 32076 34410
rect 32036 34196 32088 34202
rect 32036 34138 32088 34144
rect 32048 33590 32076 34138
rect 32036 33584 32088 33590
rect 32036 33526 32088 33532
rect 32232 32978 32260 37062
rect 32784 37046 32904 37062
rect 32404 36032 32456 36038
rect 32404 35974 32456 35980
rect 32416 35834 32444 35974
rect 32404 35828 32456 35834
rect 32404 35770 32456 35776
rect 32772 35556 32824 35562
rect 32772 35498 32824 35504
rect 32784 35154 32812 35498
rect 32772 35148 32824 35154
rect 32772 35090 32824 35096
rect 32496 34944 32548 34950
rect 32496 34886 32548 34892
rect 32404 33516 32456 33522
rect 32404 33458 32456 33464
rect 32312 33108 32364 33114
rect 32312 33050 32364 33056
rect 32220 32972 32272 32978
rect 32220 32914 32272 32920
rect 32324 32434 32352 33050
rect 32312 32428 32364 32434
rect 32312 32370 32364 32376
rect 31576 32360 31628 32366
rect 31576 32302 31628 32308
rect 31392 32292 31444 32298
rect 31392 32234 31444 32240
rect 31116 32224 31168 32230
rect 31116 32166 31168 32172
rect 31128 31822 31156 32166
rect 31404 31906 31432 32234
rect 31312 31878 31432 31906
rect 31116 31816 31168 31822
rect 31116 31758 31168 31764
rect 31312 31754 31340 31878
rect 31404 31754 31432 31878
rect 31300 31748 31352 31754
rect 31300 31690 31352 31696
rect 31392 31748 31444 31754
rect 31392 31690 31444 31696
rect 30840 31680 30892 31686
rect 30840 31622 30892 31628
rect 30852 31482 30880 31622
rect 30840 31476 30892 31482
rect 30840 31418 30892 31424
rect 30380 31408 30432 31414
rect 30380 31350 30432 31356
rect 30852 31346 30880 31418
rect 30840 31340 30892 31346
rect 30840 31282 30892 31288
rect 31588 31278 31616 32302
rect 32324 31958 32352 32370
rect 32312 31952 32364 31958
rect 32312 31894 32364 31900
rect 31668 31816 31720 31822
rect 31668 31758 31720 31764
rect 31576 31272 31628 31278
rect 31576 31214 31628 31220
rect 30840 31136 30892 31142
rect 30840 31078 30892 31084
rect 30852 30734 30880 31078
rect 31588 30734 31616 31214
rect 30380 30728 30432 30734
rect 30380 30670 30432 30676
rect 30840 30728 30892 30734
rect 30840 30670 30892 30676
rect 31576 30728 31628 30734
rect 31576 30670 31628 30676
rect 29736 29844 29788 29850
rect 29736 29786 29788 29792
rect 29748 29306 29776 29786
rect 30392 29646 30420 30670
rect 30656 29844 30708 29850
rect 30656 29786 30708 29792
rect 30380 29640 30432 29646
rect 30380 29582 30432 29588
rect 30012 29572 30064 29578
rect 30012 29514 30064 29520
rect 30024 29306 30052 29514
rect 29736 29300 29788 29306
rect 29736 29242 29788 29248
rect 30012 29300 30064 29306
rect 30012 29242 30064 29248
rect 29184 29164 29236 29170
rect 29184 29106 29236 29112
rect 29368 29164 29420 29170
rect 29368 29106 29420 29112
rect 29092 29096 29144 29102
rect 29092 29038 29144 29044
rect 29104 28506 29132 29038
rect 29196 28665 29224 29106
rect 29380 28694 29408 29106
rect 29368 28688 29420 28694
rect 29182 28656 29238 28665
rect 29368 28630 29420 28636
rect 29182 28591 29238 28600
rect 30392 28558 30420 29582
rect 29184 28552 29236 28558
rect 29104 28500 29184 28506
rect 29104 28494 29236 28500
rect 29644 28552 29696 28558
rect 29644 28494 29696 28500
rect 30380 28552 30432 28558
rect 30380 28494 30432 28500
rect 29104 28478 29224 28494
rect 29000 28416 29052 28422
rect 29000 28358 29052 28364
rect 29090 28384 29146 28393
rect 29090 28319 29146 28328
rect 29104 28082 29132 28319
rect 29092 28076 29144 28082
rect 29092 28018 29144 28024
rect 29000 28008 29052 28014
rect 29000 27950 29052 27956
rect 28816 27940 28868 27946
rect 28816 27882 28868 27888
rect 28632 27872 28684 27878
rect 28632 27814 28684 27820
rect 28816 27668 28868 27674
rect 28816 27610 28868 27616
rect 28460 27526 28580 27554
rect 28356 26988 28408 26994
rect 28356 26930 28408 26936
rect 27896 25900 27948 25906
rect 27896 25842 27948 25848
rect 27804 25220 27856 25226
rect 27804 25162 27856 25168
rect 27528 24880 27580 24886
rect 27528 24822 27580 24828
rect 27436 24676 27488 24682
rect 27436 24618 27488 24624
rect 27160 24268 27212 24274
rect 27160 24210 27212 24216
rect 26976 24132 27028 24138
rect 26976 24074 27028 24080
rect 26988 23730 27016 24074
rect 27344 23860 27396 23866
rect 27344 23802 27396 23808
rect 26976 23724 27028 23730
rect 26976 23666 27028 23672
rect 27160 23724 27212 23730
rect 27160 23666 27212 23672
rect 26884 23316 26936 23322
rect 26884 23258 26936 23264
rect 26332 23248 26384 23254
rect 26332 23190 26384 23196
rect 26976 23044 27028 23050
rect 26976 22986 27028 22992
rect 26332 22704 26384 22710
rect 26332 22646 26384 22652
rect 26344 20262 26372 22646
rect 26988 22642 27016 22986
rect 27172 22642 27200 23666
rect 27356 23662 27384 23802
rect 27448 23730 27476 24618
rect 27436 23724 27488 23730
rect 27436 23666 27488 23672
rect 27252 23656 27304 23662
rect 27252 23598 27304 23604
rect 27344 23656 27396 23662
rect 27344 23598 27396 23604
rect 27264 22778 27292 23598
rect 27356 23526 27384 23598
rect 27344 23520 27396 23526
rect 27344 23462 27396 23468
rect 27252 22772 27304 22778
rect 27252 22714 27304 22720
rect 26976 22636 27028 22642
rect 26976 22578 27028 22584
rect 27160 22636 27212 22642
rect 27160 22578 27212 22584
rect 26988 22234 27016 22578
rect 27172 22438 27200 22578
rect 27356 22574 27384 23462
rect 27540 22642 27568 24822
rect 28264 24200 28316 24206
rect 28264 24142 28316 24148
rect 28172 24132 28224 24138
rect 28172 24074 28224 24080
rect 28184 23730 28212 24074
rect 28172 23724 28224 23730
rect 28172 23666 28224 23672
rect 27528 22636 27580 22642
rect 27528 22578 27580 22584
rect 27344 22568 27396 22574
rect 27344 22510 27396 22516
rect 27160 22432 27212 22438
rect 27160 22374 27212 22380
rect 26976 22228 27028 22234
rect 26976 22170 27028 22176
rect 27356 21078 27384 22510
rect 27802 22128 27858 22137
rect 27802 22063 27804 22072
rect 27856 22063 27858 22072
rect 28172 22092 28224 22098
rect 27804 22034 27856 22040
rect 28172 22034 28224 22040
rect 28184 21894 28212 22034
rect 28172 21888 28224 21894
rect 28172 21830 28224 21836
rect 27620 21616 27672 21622
rect 27620 21558 27672 21564
rect 27528 21548 27580 21554
rect 27528 21490 27580 21496
rect 27344 21072 27396 21078
rect 27344 21014 27396 21020
rect 27068 20936 27120 20942
rect 27068 20878 27120 20884
rect 26700 20868 26752 20874
rect 26700 20810 26752 20816
rect 26712 20466 26740 20810
rect 26700 20460 26752 20466
rect 26700 20402 26752 20408
rect 26332 20256 26384 20262
rect 26332 20198 26384 20204
rect 26884 19984 26936 19990
rect 26884 19926 26936 19932
rect 26332 19916 26384 19922
rect 26332 19858 26384 19864
rect 26344 19242 26372 19858
rect 26896 19446 26924 19926
rect 27080 19514 27108 20878
rect 27540 20602 27568 21490
rect 27632 20942 27660 21558
rect 28184 21554 28212 21830
rect 28172 21548 28224 21554
rect 28172 21490 28224 21496
rect 27896 21412 27948 21418
rect 27896 21354 27948 21360
rect 27908 20942 27936 21354
rect 27620 20936 27672 20942
rect 27620 20878 27672 20884
rect 27896 20936 27948 20942
rect 27896 20878 27948 20884
rect 27620 20800 27672 20806
rect 27620 20742 27672 20748
rect 27528 20596 27580 20602
rect 27528 20538 27580 20544
rect 27632 20534 27660 20742
rect 27620 20528 27672 20534
rect 27620 20470 27672 20476
rect 27252 20392 27304 20398
rect 27252 20334 27304 20340
rect 27160 20256 27212 20262
rect 27160 20198 27212 20204
rect 27068 19508 27120 19514
rect 27068 19450 27120 19456
rect 26884 19440 26936 19446
rect 26884 19382 26936 19388
rect 26332 19236 26384 19242
rect 26332 19178 26384 19184
rect 26240 18964 26292 18970
rect 26240 18906 26292 18912
rect 25504 18896 25556 18902
rect 25504 18838 25556 18844
rect 26252 17882 26280 18906
rect 26240 17876 26292 17882
rect 26240 17818 26292 17824
rect 26884 17604 26936 17610
rect 26884 17546 26936 17552
rect 25596 17196 25648 17202
rect 25596 17138 25648 17144
rect 25608 16590 25636 17138
rect 26896 17134 26924 17546
rect 26884 17128 26936 17134
rect 26884 17070 26936 17076
rect 26240 16720 26292 16726
rect 26240 16662 26292 16668
rect 25596 16584 25648 16590
rect 25596 16526 25648 16532
rect 25136 16448 25188 16454
rect 25136 16390 25188 16396
rect 25608 16046 25636 16526
rect 26148 16448 26200 16454
rect 26148 16390 26200 16396
rect 26160 16182 26188 16390
rect 26148 16176 26200 16182
rect 26148 16118 26200 16124
rect 25596 16040 25648 16046
rect 25596 15982 25648 15988
rect 26160 15910 26188 16118
rect 26252 16114 26280 16662
rect 26240 16108 26292 16114
rect 26240 16050 26292 16056
rect 26700 16108 26752 16114
rect 26700 16050 26752 16056
rect 24860 15904 24912 15910
rect 24860 15846 24912 15852
rect 25596 15904 25648 15910
rect 25596 15846 25648 15852
rect 26148 15904 26200 15910
rect 26148 15846 26200 15852
rect 24872 15570 24900 15846
rect 24860 15564 24912 15570
rect 24860 15506 24912 15512
rect 24768 15496 24820 15502
rect 24768 15438 24820 15444
rect 24780 15094 24808 15438
rect 25608 15162 25636 15846
rect 26712 15502 26740 16050
rect 26700 15496 26752 15502
rect 26700 15438 26752 15444
rect 25596 15156 25648 15162
rect 25596 15098 25648 15104
rect 24768 15088 24820 15094
rect 24768 15030 24820 15036
rect 24676 14816 24728 14822
rect 24676 14758 24728 14764
rect 25228 14816 25280 14822
rect 25228 14758 25280 14764
rect 24400 14068 24452 14074
rect 24400 14010 24452 14016
rect 24504 14028 24808 14056
rect 24504 13954 24532 14028
rect 24320 13926 24532 13954
rect 24584 13932 24636 13938
rect 24584 13874 24636 13880
rect 24216 13184 24268 13190
rect 24216 13126 24268 13132
rect 24228 12850 24256 13126
rect 24216 12844 24268 12850
rect 24216 12786 24268 12792
rect 24124 12776 24176 12782
rect 24124 12718 24176 12724
rect 24136 11898 24164 12718
rect 24400 12640 24452 12646
rect 24400 12582 24452 12588
rect 24412 12442 24440 12582
rect 24400 12436 24452 12442
rect 24400 12378 24452 12384
rect 24124 11892 24176 11898
rect 24124 11834 24176 11840
rect 24596 11558 24624 13874
rect 24676 13864 24728 13870
rect 24676 13806 24728 13812
rect 24688 13326 24716 13806
rect 24676 13320 24728 13326
rect 24676 13262 24728 13268
rect 24688 12714 24716 13262
rect 24676 12708 24728 12714
rect 24676 12650 24728 12656
rect 24780 12442 24808 14028
rect 25240 13938 25268 14758
rect 26712 14414 26740 15438
rect 26884 15360 26936 15366
rect 26884 15302 26936 15308
rect 26896 15026 26924 15302
rect 26884 15020 26936 15026
rect 26884 14962 26936 14968
rect 26240 14408 26292 14414
rect 26240 14350 26292 14356
rect 26700 14408 26752 14414
rect 26700 14350 26752 14356
rect 26148 14340 26200 14346
rect 26148 14282 26200 14288
rect 26160 14074 26188 14282
rect 26148 14068 26200 14074
rect 26148 14010 26200 14016
rect 25228 13932 25280 13938
rect 25228 13874 25280 13880
rect 25136 13524 25188 13530
rect 25136 13466 25188 13472
rect 25148 12782 25176 13466
rect 25240 13394 25268 13874
rect 25320 13728 25372 13734
rect 25320 13670 25372 13676
rect 25228 13388 25280 13394
rect 25228 13330 25280 13336
rect 25332 13326 25360 13670
rect 25320 13320 25372 13326
rect 25320 13262 25372 13268
rect 25136 12776 25188 12782
rect 25136 12718 25188 12724
rect 26252 12714 26280 14350
rect 26896 14346 26924 14962
rect 26884 14340 26936 14346
rect 26884 14282 26936 14288
rect 26976 12776 27028 12782
rect 26976 12718 27028 12724
rect 26056 12708 26108 12714
rect 26056 12650 26108 12656
rect 26240 12708 26292 12714
rect 26240 12650 26292 12656
rect 24768 12436 24820 12442
rect 24768 12378 24820 12384
rect 26068 12238 26096 12650
rect 26988 12646 27016 12718
rect 26332 12640 26384 12646
rect 26332 12582 26384 12588
rect 26976 12640 27028 12646
rect 26976 12582 27028 12588
rect 26344 12238 26372 12582
rect 25136 12232 25188 12238
rect 25136 12174 25188 12180
rect 26056 12232 26108 12238
rect 26056 12174 26108 12180
rect 26332 12232 26384 12238
rect 26332 12174 26384 12180
rect 24584 11552 24636 11558
rect 24584 11494 24636 11500
rect 24032 11348 24084 11354
rect 24032 11290 24084 11296
rect 22560 10260 22612 10266
rect 22560 10202 22612 10208
rect 23480 10260 23532 10266
rect 23480 10202 23532 10208
rect 22560 10056 22612 10062
rect 22560 9998 22612 10004
rect 22468 9512 22520 9518
rect 22468 9454 22520 9460
rect 22572 9178 22600 9998
rect 23572 9580 23624 9586
rect 23572 9522 23624 9528
rect 23020 9512 23072 9518
rect 23020 9454 23072 9460
rect 22928 9444 22980 9450
rect 22928 9386 22980 9392
rect 22652 9376 22704 9382
rect 22652 9318 22704 9324
rect 22836 9376 22888 9382
rect 22836 9318 22888 9324
rect 22376 9172 22428 9178
rect 22376 9114 22428 9120
rect 22560 9172 22612 9178
rect 22560 9114 22612 9120
rect 22664 8974 22692 9318
rect 22652 8968 22704 8974
rect 22652 8910 22704 8916
rect 22192 8628 22244 8634
rect 22192 8570 22244 8576
rect 22848 8566 22876 9318
rect 22836 8560 22888 8566
rect 22836 8502 22888 8508
rect 20720 8492 20772 8498
rect 20720 8434 20772 8440
rect 20996 8492 21048 8498
rect 20996 8434 21048 8440
rect 21732 8492 21784 8498
rect 21732 8434 21784 8440
rect 22008 8492 22060 8498
rect 22008 8434 22060 8440
rect 20628 8084 20680 8090
rect 20628 8026 20680 8032
rect 20640 7410 20668 8026
rect 20720 7812 20772 7818
rect 20720 7754 20772 7760
rect 20628 7404 20680 7410
rect 20628 7346 20680 7352
rect 20260 6792 20312 6798
rect 20260 6734 20312 6740
rect 20732 6662 20760 7754
rect 21008 7342 21036 8434
rect 22020 8090 22048 8434
rect 22008 8084 22060 8090
rect 22008 8026 22060 8032
rect 22940 7886 22968 9386
rect 23032 8498 23060 9454
rect 23020 8492 23072 8498
rect 23020 8434 23072 8440
rect 23032 7954 23060 8434
rect 23584 8090 23612 9522
rect 23756 8832 23808 8838
rect 23756 8774 23808 8780
rect 23572 8084 23624 8090
rect 23572 8026 23624 8032
rect 23020 7948 23072 7954
rect 23020 7890 23072 7896
rect 22928 7880 22980 7886
rect 22928 7822 22980 7828
rect 23032 7410 23060 7890
rect 23768 7886 23796 8774
rect 23756 7880 23808 7886
rect 23756 7822 23808 7828
rect 23572 7744 23624 7750
rect 23572 7686 23624 7692
rect 23584 7478 23612 7686
rect 23572 7472 23624 7478
rect 23572 7414 23624 7420
rect 23020 7404 23072 7410
rect 23020 7346 23072 7352
rect 20996 7336 21048 7342
rect 20996 7278 21048 7284
rect 24596 7274 24624 11494
rect 25148 9450 25176 12174
rect 26068 11694 26096 12174
rect 26988 11762 27016 12582
rect 27172 11830 27200 20198
rect 27264 19854 27292 20334
rect 27908 20330 27936 20878
rect 28172 20868 28224 20874
rect 28172 20810 28224 20816
rect 28184 20466 28212 20810
rect 28172 20460 28224 20466
rect 28172 20402 28224 20408
rect 27896 20324 27948 20330
rect 27896 20266 27948 20272
rect 28276 19990 28304 24142
rect 28368 24070 28396 26930
rect 28460 26926 28488 27526
rect 28540 27464 28592 27470
rect 28540 27406 28592 27412
rect 28632 27464 28684 27470
rect 28632 27406 28684 27412
rect 28448 26920 28500 26926
rect 28448 26862 28500 26868
rect 28448 26376 28500 26382
rect 28448 26318 28500 26324
rect 28460 24954 28488 26318
rect 28552 26314 28580 27406
rect 28644 27334 28672 27406
rect 28632 27328 28684 27334
rect 28632 27270 28684 27276
rect 28828 26994 28856 27610
rect 29012 27538 29040 27950
rect 29092 27940 29144 27946
rect 29092 27882 29144 27888
rect 29104 27674 29132 27882
rect 29092 27668 29144 27674
rect 29092 27610 29144 27616
rect 28908 27532 28960 27538
rect 28908 27474 28960 27480
rect 29000 27532 29052 27538
rect 29000 27474 29052 27480
rect 28920 27334 28948 27474
rect 29012 27402 29040 27474
rect 29092 27464 29144 27470
rect 29092 27406 29144 27412
rect 29000 27396 29052 27402
rect 29000 27338 29052 27344
rect 28908 27328 28960 27334
rect 28908 27270 28960 27276
rect 28816 26988 28868 26994
rect 28816 26930 28868 26936
rect 28828 26586 28856 26930
rect 28816 26580 28868 26586
rect 28816 26522 28868 26528
rect 28540 26308 28592 26314
rect 28540 26250 28592 26256
rect 28552 25294 28580 26250
rect 28724 26240 28776 26246
rect 28724 26182 28776 26188
rect 28736 25498 28764 26182
rect 28828 26042 28856 26522
rect 29012 26466 29040 27338
rect 28920 26438 29040 26466
rect 29104 26450 29132 27406
rect 29196 26994 29224 28478
rect 29276 28416 29328 28422
rect 29276 28358 29328 28364
rect 29288 27946 29316 28358
rect 29656 28218 29684 28494
rect 29644 28212 29696 28218
rect 29644 28154 29696 28160
rect 29276 27940 29328 27946
rect 29276 27882 29328 27888
rect 29368 27940 29420 27946
rect 29368 27882 29420 27888
rect 29380 27470 29408 27882
rect 30392 27878 30420 28494
rect 30472 28484 30524 28490
rect 30472 28426 30524 28432
rect 30484 28218 30512 28426
rect 30472 28212 30524 28218
rect 30472 28154 30524 28160
rect 30380 27872 30432 27878
rect 30380 27814 30432 27820
rect 30104 27600 30156 27606
rect 30104 27542 30156 27548
rect 29368 27464 29420 27470
rect 29368 27406 29420 27412
rect 29828 27328 29880 27334
rect 29828 27270 29880 27276
rect 29184 26988 29236 26994
rect 29184 26930 29236 26936
rect 29368 26512 29420 26518
rect 29368 26454 29420 26460
rect 29092 26444 29144 26450
rect 28816 26036 28868 26042
rect 28816 25978 28868 25984
rect 28920 25906 28948 26438
rect 29092 26386 29144 26392
rect 29000 26376 29052 26382
rect 29000 26318 29052 26324
rect 29012 26042 29040 26318
rect 29000 26036 29052 26042
rect 29000 25978 29052 25984
rect 28908 25900 28960 25906
rect 28908 25842 28960 25848
rect 29184 25900 29236 25906
rect 29184 25842 29236 25848
rect 28724 25492 28776 25498
rect 28724 25434 28776 25440
rect 28540 25288 28592 25294
rect 28540 25230 28592 25236
rect 28448 24948 28500 24954
rect 28448 24890 28500 24896
rect 28356 24064 28408 24070
rect 28356 24006 28408 24012
rect 28460 22760 28488 24890
rect 28540 24268 28592 24274
rect 28540 24210 28592 24216
rect 28552 23730 28580 24210
rect 28724 24200 28776 24206
rect 28724 24142 28776 24148
rect 28736 23798 28764 24142
rect 29196 24138 29224 25842
rect 29380 24818 29408 26454
rect 29840 26450 29868 27270
rect 30012 26784 30064 26790
rect 30012 26726 30064 26732
rect 29828 26444 29880 26450
rect 29828 26386 29880 26392
rect 29552 25900 29604 25906
rect 29552 25842 29604 25848
rect 29564 24954 29592 25842
rect 30024 25378 30052 26726
rect 30116 25498 30144 27542
rect 30196 27532 30248 27538
rect 30196 27474 30248 27480
rect 30208 26450 30236 27474
rect 30288 27328 30340 27334
rect 30288 27270 30340 27276
rect 30300 26790 30328 27270
rect 30288 26784 30340 26790
rect 30288 26726 30340 26732
rect 30288 26580 30340 26586
rect 30288 26522 30340 26528
rect 30196 26444 30248 26450
rect 30196 26386 30248 26392
rect 30104 25492 30156 25498
rect 30104 25434 30156 25440
rect 30024 25350 30236 25378
rect 29552 24948 29604 24954
rect 29552 24890 29604 24896
rect 29368 24812 29420 24818
rect 29368 24754 29420 24760
rect 29644 24404 29696 24410
rect 29644 24346 29696 24352
rect 29276 24336 29328 24342
rect 29276 24278 29328 24284
rect 28908 24132 28960 24138
rect 28908 24074 28960 24080
rect 29184 24132 29236 24138
rect 29184 24074 29236 24080
rect 28724 23792 28776 23798
rect 28724 23734 28776 23740
rect 28540 23724 28592 23730
rect 28540 23666 28592 23672
rect 28816 23180 28868 23186
rect 28920 23168 28948 24074
rect 29288 23730 29316 24278
rect 29368 24064 29420 24070
rect 29368 24006 29420 24012
rect 29460 24064 29512 24070
rect 29460 24006 29512 24012
rect 29380 23730 29408 24006
rect 29472 23866 29500 24006
rect 29460 23860 29512 23866
rect 29460 23802 29512 23808
rect 29276 23724 29328 23730
rect 29276 23666 29328 23672
rect 29368 23724 29420 23730
rect 29368 23666 29420 23672
rect 29184 23656 29236 23662
rect 29184 23598 29236 23604
rect 28868 23140 28948 23168
rect 28816 23122 28868 23128
rect 28828 22982 28856 23122
rect 28816 22976 28868 22982
rect 28816 22918 28868 22924
rect 28460 22732 28580 22760
rect 28356 22636 28408 22642
rect 28356 22578 28408 22584
rect 28448 22636 28500 22642
rect 28448 22578 28500 22584
rect 28368 22166 28396 22578
rect 28356 22160 28408 22166
rect 28356 22102 28408 22108
rect 28368 21622 28396 22102
rect 28460 22030 28488 22578
rect 28448 22024 28500 22030
rect 28448 21966 28500 21972
rect 28356 21616 28408 21622
rect 28356 21558 28408 21564
rect 28264 19984 28316 19990
rect 28264 19926 28316 19932
rect 28368 19922 28396 21558
rect 28460 21486 28488 21966
rect 28552 21672 28580 22732
rect 28724 22432 28776 22438
rect 28724 22374 28776 22380
rect 28552 21644 28672 21672
rect 28540 21548 28592 21554
rect 28540 21490 28592 21496
rect 28448 21480 28500 21486
rect 28448 21422 28500 21428
rect 28448 21072 28500 21078
rect 28448 21014 28500 21020
rect 27344 19916 27396 19922
rect 27344 19858 27396 19864
rect 28356 19916 28408 19922
rect 28356 19858 28408 19864
rect 27252 19848 27304 19854
rect 27252 19790 27304 19796
rect 27356 19378 27384 19858
rect 27344 19372 27396 19378
rect 27344 19314 27396 19320
rect 27804 17672 27856 17678
rect 27804 17614 27856 17620
rect 27816 16794 27844 17614
rect 27712 16788 27764 16794
rect 27712 16730 27764 16736
rect 27804 16788 27856 16794
rect 27804 16730 27856 16736
rect 27724 15502 27752 16730
rect 28460 15706 28488 21014
rect 28552 20262 28580 21490
rect 28644 21146 28672 21644
rect 28632 21140 28684 21146
rect 28632 21082 28684 21088
rect 28736 21026 28764 22374
rect 28644 20998 28764 21026
rect 28540 20256 28592 20262
rect 28540 20198 28592 20204
rect 28644 18290 28672 20998
rect 28828 20942 28856 22918
rect 29196 22642 29224 23598
rect 29092 22636 29144 22642
rect 29092 22578 29144 22584
rect 29184 22636 29236 22642
rect 29184 22578 29236 22584
rect 28954 22160 29006 22166
rect 28906 22128 28954 22137
rect 28962 22102 29006 22108
rect 28962 22086 28994 22102
rect 28906 22063 28962 22072
rect 29000 22024 29052 22030
rect 28908 22002 28960 22008
rect 29000 21966 29052 21972
rect 28908 21944 28960 21950
rect 28724 20936 28776 20942
rect 28724 20878 28776 20884
rect 28816 20936 28868 20942
rect 28816 20878 28868 20884
rect 28736 20788 28764 20878
rect 28920 20788 28948 21944
rect 29012 21690 29040 21966
rect 29000 21684 29052 21690
rect 29000 21626 29052 21632
rect 29104 21146 29132 22578
rect 29472 21894 29500 23802
rect 29656 23594 29684 24346
rect 29552 23588 29604 23594
rect 29552 23530 29604 23536
rect 29644 23588 29696 23594
rect 29644 23530 29696 23536
rect 29564 23186 29592 23530
rect 29552 23180 29604 23186
rect 29552 23122 29604 23128
rect 29656 23066 29684 23530
rect 30104 23520 30156 23526
rect 30104 23462 30156 23468
rect 29564 23038 29684 23066
rect 29564 22574 29592 23038
rect 29828 22636 29880 22642
rect 29828 22578 29880 22584
rect 29552 22568 29604 22574
rect 29552 22510 29604 22516
rect 29564 22166 29592 22510
rect 29736 22500 29788 22506
rect 29736 22442 29788 22448
rect 29644 22228 29696 22234
rect 29644 22170 29696 22176
rect 29552 22160 29604 22166
rect 29552 22102 29604 22108
rect 29460 21888 29512 21894
rect 29460 21830 29512 21836
rect 29276 21548 29328 21554
rect 29276 21490 29328 21496
rect 29288 21350 29316 21490
rect 29276 21344 29328 21350
rect 29276 21286 29328 21292
rect 29092 21140 29144 21146
rect 29092 21082 29144 21088
rect 28736 20760 28948 20788
rect 28736 20466 28764 20760
rect 29656 20602 29684 22170
rect 29748 22098 29776 22442
rect 29840 22234 29868 22578
rect 29828 22228 29880 22234
rect 29828 22170 29880 22176
rect 29736 22092 29788 22098
rect 29736 22034 29788 22040
rect 29736 21956 29788 21962
rect 29736 21898 29788 21904
rect 29748 21690 29776 21898
rect 29736 21684 29788 21690
rect 29736 21626 29788 21632
rect 29644 20596 29696 20602
rect 29644 20538 29696 20544
rect 30012 20596 30064 20602
rect 30012 20538 30064 20544
rect 28724 20460 28776 20466
rect 28724 20402 28776 20408
rect 29552 20256 29604 20262
rect 29552 20198 29604 20204
rect 29564 19378 29592 20198
rect 28724 19372 28776 19378
rect 28724 19314 28776 19320
rect 29552 19372 29604 19378
rect 29552 19314 29604 19320
rect 29920 19372 29972 19378
rect 29920 19314 29972 19320
rect 28736 18426 28764 19314
rect 29000 19236 29052 19242
rect 29000 19178 29052 19184
rect 28816 19168 28868 19174
rect 28816 19110 28868 19116
rect 28828 18834 28856 19110
rect 28816 18828 28868 18834
rect 28816 18770 28868 18776
rect 28724 18420 28776 18426
rect 28724 18362 28776 18368
rect 28632 18284 28684 18290
rect 28632 18226 28684 18232
rect 28828 17762 28856 18770
rect 29012 18766 29040 19178
rect 29828 19168 29880 19174
rect 29828 19110 29880 19116
rect 29840 18766 29868 19110
rect 29000 18760 29052 18766
rect 29000 18702 29052 18708
rect 29828 18760 29880 18766
rect 29828 18702 29880 18708
rect 29932 18698 29960 19314
rect 30024 18834 30052 20538
rect 30116 19854 30144 23462
rect 30208 22030 30236 25350
rect 30300 25158 30328 26522
rect 30392 25702 30420 27814
rect 30380 25696 30432 25702
rect 30380 25638 30432 25644
rect 30668 25514 30696 29786
rect 30748 29504 30800 29510
rect 30748 29446 30800 29452
rect 30760 29170 30788 29446
rect 30748 29164 30800 29170
rect 30748 29106 30800 29112
rect 30760 27402 30788 29106
rect 31680 28762 31708 31758
rect 32324 31754 32352 31894
rect 32232 31726 32352 31754
rect 32232 31414 32260 31726
rect 32416 31686 32444 33458
rect 32508 32910 32536 34886
rect 32876 34678 32904 37046
rect 32968 36718 32996 37198
rect 34532 37126 34560 37810
rect 34808 37806 34836 38286
rect 34796 37800 34848 37806
rect 34796 37742 34848 37748
rect 34520 37120 34572 37126
rect 34520 37062 34572 37068
rect 34808 36718 34836 37742
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 35912 37210 35940 39374
rect 36084 38956 36136 38962
rect 36084 38898 36136 38904
rect 36452 38956 36504 38962
rect 36452 38898 36504 38904
rect 38108 38956 38160 38962
rect 38108 38898 38160 38904
rect 35992 38752 36044 38758
rect 35992 38694 36044 38700
rect 36004 38282 36032 38694
rect 35992 38276 36044 38282
rect 35992 38218 36044 38224
rect 36096 38010 36124 38898
rect 36084 38004 36136 38010
rect 36084 37946 36136 37952
rect 36464 37806 36492 38898
rect 36912 38888 36964 38894
rect 36912 38830 36964 38836
rect 36924 38554 36952 38830
rect 36912 38548 36964 38554
rect 36912 38490 36964 38496
rect 36924 37874 36952 38490
rect 37556 38208 37608 38214
rect 37556 38150 37608 38156
rect 37568 37874 37596 38150
rect 38120 38010 38148 38898
rect 38212 38826 38240 39986
rect 40144 39574 40172 40938
rect 40316 40520 40368 40526
rect 40316 40462 40368 40468
rect 40328 39846 40356 40462
rect 40316 39840 40368 39846
rect 40316 39782 40368 39788
rect 40132 39568 40184 39574
rect 40132 39510 40184 39516
rect 39764 39432 39816 39438
rect 39764 39374 39816 39380
rect 39776 39098 39804 39374
rect 40224 39296 40276 39302
rect 40224 39238 40276 39244
rect 39764 39092 39816 39098
rect 39764 39034 39816 39040
rect 38200 38820 38252 38826
rect 38200 38762 38252 38768
rect 38660 38752 38712 38758
rect 38660 38694 38712 38700
rect 38672 38350 38700 38694
rect 38660 38344 38712 38350
rect 38660 38286 38712 38292
rect 38936 38344 38988 38350
rect 38936 38286 38988 38292
rect 38108 38004 38160 38010
rect 38108 37946 38160 37952
rect 38844 38004 38896 38010
rect 38844 37946 38896 37952
rect 36912 37868 36964 37874
rect 36912 37810 36964 37816
rect 37556 37868 37608 37874
rect 37556 37810 37608 37816
rect 38660 37868 38712 37874
rect 38660 37810 38712 37816
rect 36452 37800 36504 37806
rect 36452 37742 36504 37748
rect 36360 37732 36412 37738
rect 36360 37674 36412 37680
rect 35912 37182 36032 37210
rect 35900 37120 35952 37126
rect 35900 37062 35952 37068
rect 35440 36780 35492 36786
rect 35440 36722 35492 36728
rect 32956 36712 33008 36718
rect 32956 36654 33008 36660
rect 34796 36712 34848 36718
rect 34796 36654 34848 36660
rect 32968 36242 32996 36654
rect 33784 36576 33836 36582
rect 33784 36518 33836 36524
rect 33796 36310 33824 36518
rect 33784 36304 33836 36310
rect 33784 36246 33836 36252
rect 34520 36304 34572 36310
rect 34520 36246 34572 36252
rect 32956 36236 33008 36242
rect 32956 36178 33008 36184
rect 32968 35086 32996 36178
rect 33140 36168 33192 36174
rect 33140 36110 33192 36116
rect 33152 36038 33180 36110
rect 33140 36032 33192 36038
rect 33140 35974 33192 35980
rect 32956 35080 33008 35086
rect 32956 35022 33008 35028
rect 32968 34678 32996 35022
rect 33152 35018 33180 35974
rect 34532 35766 34560 36246
rect 34520 35760 34572 35766
rect 34520 35702 34572 35708
rect 34808 35630 34836 36654
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 35348 36236 35400 36242
rect 35348 36178 35400 36184
rect 34796 35624 34848 35630
rect 34796 35566 34848 35572
rect 34808 35154 34836 35566
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 34796 35148 34848 35154
rect 34796 35090 34848 35096
rect 33140 35012 33192 35018
rect 33140 34954 33192 34960
rect 33508 35012 33560 35018
rect 33508 34954 33560 34960
rect 33520 34678 33548 34954
rect 32864 34672 32916 34678
rect 32864 34614 32916 34620
rect 32956 34672 33008 34678
rect 32956 34614 33008 34620
rect 33508 34672 33560 34678
rect 33508 34614 33560 34620
rect 32680 33516 32732 33522
rect 32680 33458 32732 33464
rect 32496 32904 32548 32910
rect 32496 32846 32548 32852
rect 32496 32768 32548 32774
rect 32692 32756 32720 33458
rect 32548 32728 32720 32756
rect 32496 32710 32548 32716
rect 32692 32434 32720 32728
rect 32680 32428 32732 32434
rect 32680 32370 32732 32376
rect 32876 32366 32904 34614
rect 34808 34542 34836 35090
rect 34520 34536 34572 34542
rect 34520 34478 34572 34484
rect 34796 34536 34848 34542
rect 34796 34478 34848 34484
rect 33968 34400 34020 34406
rect 33968 34342 34020 34348
rect 33876 33992 33928 33998
rect 33876 33934 33928 33940
rect 33232 33380 33284 33386
rect 33232 33322 33284 33328
rect 32956 33040 33008 33046
rect 32956 32982 33008 32988
rect 32968 32842 32996 32982
rect 33244 32910 33272 33322
rect 33232 32904 33284 32910
rect 33232 32846 33284 32852
rect 32956 32836 33008 32842
rect 32956 32778 33008 32784
rect 33416 32768 33468 32774
rect 33416 32710 33468 32716
rect 33428 32502 33456 32710
rect 33416 32496 33468 32502
rect 33416 32438 33468 32444
rect 33888 32366 33916 33934
rect 33980 33930 34008 34342
rect 33968 33924 34020 33930
rect 33968 33866 34020 33872
rect 34060 32972 34112 32978
rect 34060 32914 34112 32920
rect 32864 32360 32916 32366
rect 32864 32302 32916 32308
rect 33876 32360 33928 32366
rect 33876 32302 33928 32308
rect 33888 32026 33916 32302
rect 33876 32020 33928 32026
rect 33876 31962 33928 31968
rect 33140 31884 33192 31890
rect 33140 31826 33192 31832
rect 32312 31680 32364 31686
rect 32312 31622 32364 31628
rect 32404 31680 32456 31686
rect 32404 31622 32456 31628
rect 32324 31482 32352 31622
rect 32312 31476 32364 31482
rect 32312 31418 32364 31424
rect 32220 31408 32272 31414
rect 32220 31350 32272 31356
rect 32416 31142 32444 31622
rect 33152 31414 33180 31826
rect 33324 31816 33376 31822
rect 33324 31758 33376 31764
rect 33336 31686 33364 31758
rect 33232 31680 33284 31686
rect 33232 31622 33284 31628
rect 33324 31680 33376 31686
rect 33324 31622 33376 31628
rect 33140 31408 33192 31414
rect 33140 31350 33192 31356
rect 32772 31204 32824 31210
rect 32772 31146 32824 31152
rect 32404 31136 32456 31142
rect 32404 31078 32456 31084
rect 32416 30938 32444 31078
rect 32784 30938 32812 31146
rect 32404 30932 32456 30938
rect 32404 30874 32456 30880
rect 32772 30932 32824 30938
rect 32772 30874 32824 30880
rect 33244 30734 33272 31622
rect 34072 31482 34100 32914
rect 34152 32836 34204 32842
rect 34152 32778 34204 32784
rect 34164 31890 34192 32778
rect 34428 32564 34480 32570
rect 34428 32506 34480 32512
rect 34152 31884 34204 31890
rect 34152 31826 34204 31832
rect 34060 31476 34112 31482
rect 34060 31418 34112 31424
rect 33232 30728 33284 30734
rect 33232 30670 33284 30676
rect 33968 30728 34020 30734
rect 33968 30670 34020 30676
rect 33416 30660 33468 30666
rect 33416 30602 33468 30608
rect 32680 30592 32732 30598
rect 32680 30534 32732 30540
rect 32692 30258 32720 30534
rect 33428 30326 33456 30602
rect 33416 30320 33468 30326
rect 33416 30262 33468 30268
rect 32680 30252 32732 30258
rect 32680 30194 32732 30200
rect 32680 30048 32732 30054
rect 32680 29990 32732 29996
rect 32692 29646 32720 29990
rect 33980 29850 34008 30670
rect 34164 30598 34192 31826
rect 34440 31754 34468 32506
rect 34532 32502 34560 34478
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 35360 34134 35388 36178
rect 35452 35834 35480 36722
rect 35912 36378 35940 37062
rect 35900 36372 35952 36378
rect 35900 36314 35952 36320
rect 35716 36032 35768 36038
rect 35716 35974 35768 35980
rect 35440 35828 35492 35834
rect 35440 35770 35492 35776
rect 35728 35698 35756 35974
rect 35716 35692 35768 35698
rect 35716 35634 35768 35640
rect 35532 35080 35584 35086
rect 35532 35022 35584 35028
rect 35900 35080 35952 35086
rect 35900 35022 35952 35028
rect 35544 34202 35572 35022
rect 35624 34944 35676 34950
rect 35624 34886 35676 34892
rect 35636 34678 35664 34886
rect 35624 34672 35676 34678
rect 35624 34614 35676 34620
rect 35912 34202 35940 35022
rect 35532 34196 35584 34202
rect 35532 34138 35584 34144
rect 35900 34196 35952 34202
rect 35900 34138 35952 34144
rect 35348 34128 35400 34134
rect 35348 34070 35400 34076
rect 35360 33590 35388 34070
rect 35624 34060 35676 34066
rect 35624 34002 35676 34008
rect 35348 33584 35400 33590
rect 35348 33526 35400 33532
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 35360 32978 35388 33526
rect 35348 32972 35400 32978
rect 35348 32914 35400 32920
rect 34704 32904 34756 32910
rect 34704 32846 34756 32852
rect 34716 32570 34744 32846
rect 34704 32564 34756 32570
rect 34704 32506 34756 32512
rect 34520 32496 34572 32502
rect 34520 32438 34572 32444
rect 34256 31726 34468 31754
rect 34152 30592 34204 30598
rect 34152 30534 34204 30540
rect 34164 30394 34192 30534
rect 34152 30388 34204 30394
rect 34152 30330 34204 30336
rect 34256 30138 34284 31726
rect 34428 31680 34480 31686
rect 34428 31622 34480 31628
rect 34440 31482 34468 31622
rect 34428 31476 34480 31482
rect 34428 31418 34480 31424
rect 34532 31414 34560 32438
rect 34520 31408 34572 31414
rect 34520 31350 34572 31356
rect 34428 31340 34480 31346
rect 34428 31282 34480 31288
rect 34336 31136 34388 31142
rect 34336 31078 34388 31084
rect 34348 30938 34376 31078
rect 34336 30932 34388 30938
rect 34336 30874 34388 30880
rect 34348 30190 34376 30874
rect 34440 30734 34468 31282
rect 34428 30728 34480 30734
rect 34428 30670 34480 30676
rect 34532 30326 34560 31350
rect 34716 31142 34744 32506
rect 34796 32224 34848 32230
rect 34796 32166 34848 32172
rect 34808 31890 34836 32166
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 34796 31884 34848 31890
rect 34796 31826 34848 31832
rect 34980 31884 35032 31890
rect 34980 31826 35032 31832
rect 34808 31210 34836 31826
rect 34992 31210 35020 31826
rect 35532 31408 35584 31414
rect 35532 31350 35584 31356
rect 35440 31340 35492 31346
rect 35440 31282 35492 31288
rect 34796 31204 34848 31210
rect 34796 31146 34848 31152
rect 34980 31204 35032 31210
rect 34980 31146 35032 31152
rect 34704 31136 34756 31142
rect 34704 31078 34756 31084
rect 34716 30666 34744 31078
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 35348 30932 35400 30938
rect 35348 30874 35400 30880
rect 34796 30864 34848 30870
rect 35164 30864 35216 30870
rect 34848 30812 35164 30818
rect 34796 30806 35216 30812
rect 34808 30790 35204 30806
rect 34704 30660 34756 30666
rect 34704 30602 34756 30608
rect 34520 30320 34572 30326
rect 34520 30262 34572 30268
rect 35360 30258 35388 30874
rect 35452 30802 35480 31282
rect 35440 30796 35492 30802
rect 35440 30738 35492 30744
rect 35348 30252 35400 30258
rect 35348 30194 35400 30200
rect 34164 30122 34284 30138
rect 34336 30184 34388 30190
rect 34336 30126 34388 30132
rect 34152 30116 34284 30122
rect 34204 30110 34284 30116
rect 34152 30058 34204 30064
rect 34244 30048 34296 30054
rect 34244 29990 34296 29996
rect 33968 29844 34020 29850
rect 33968 29786 34020 29792
rect 32680 29640 32732 29646
rect 32680 29582 32732 29588
rect 34256 29170 34284 29990
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 35452 29850 35480 30738
rect 35544 30734 35572 31350
rect 35636 30802 35664 34002
rect 35808 32904 35860 32910
rect 35808 32846 35860 32852
rect 35716 32768 35768 32774
rect 35716 32710 35768 32716
rect 35728 32434 35756 32710
rect 35820 32434 35848 32846
rect 35716 32428 35768 32434
rect 35716 32370 35768 32376
rect 35808 32428 35860 32434
rect 35808 32370 35860 32376
rect 35624 30796 35676 30802
rect 35624 30738 35676 30744
rect 35532 30728 35584 30734
rect 35532 30670 35584 30676
rect 35544 30394 35572 30670
rect 35532 30388 35584 30394
rect 35532 30330 35584 30336
rect 35440 29844 35492 29850
rect 35440 29786 35492 29792
rect 34704 29640 34756 29646
rect 34704 29582 34756 29588
rect 34244 29164 34296 29170
rect 34244 29106 34296 29112
rect 31668 28756 31720 28762
rect 31668 28698 31720 28704
rect 31392 28416 31444 28422
rect 31392 28358 31444 28364
rect 31300 28076 31352 28082
rect 31404 28064 31432 28358
rect 31680 28098 31708 28698
rect 31496 28082 31708 28098
rect 32772 28144 32824 28150
rect 32772 28086 32824 28092
rect 33232 28144 33284 28150
rect 33232 28086 33284 28092
rect 31352 28036 31432 28064
rect 31300 28018 31352 28024
rect 30748 27396 30800 27402
rect 30748 27338 30800 27344
rect 30760 27146 30788 27338
rect 31404 27334 31432 28036
rect 31484 28076 31708 28082
rect 31536 28070 31708 28076
rect 32588 28076 32640 28082
rect 31484 28018 31536 28024
rect 32588 28018 32640 28024
rect 32496 27940 32548 27946
rect 32496 27882 32548 27888
rect 31668 27872 31720 27878
rect 31668 27814 31720 27820
rect 31680 27538 31708 27814
rect 31668 27532 31720 27538
rect 31668 27474 31720 27480
rect 31392 27328 31444 27334
rect 31392 27270 31444 27276
rect 30760 27118 30880 27146
rect 30748 26988 30800 26994
rect 30748 26930 30800 26936
rect 30760 26382 30788 26930
rect 30852 26926 30880 27118
rect 31404 26994 31432 27270
rect 31392 26988 31444 26994
rect 31392 26930 31444 26936
rect 30840 26920 30892 26926
rect 30840 26862 30892 26868
rect 30748 26376 30800 26382
rect 30748 26318 30800 26324
rect 30760 26042 30788 26318
rect 30748 26036 30800 26042
rect 30748 25978 30800 25984
rect 30840 25696 30892 25702
rect 30840 25638 30892 25644
rect 30472 25492 30524 25498
rect 30668 25486 30788 25514
rect 30472 25434 30524 25440
rect 30484 25294 30512 25434
rect 30656 25356 30708 25362
rect 30656 25298 30708 25304
rect 30472 25288 30524 25294
rect 30472 25230 30524 25236
rect 30288 25152 30340 25158
rect 30288 25094 30340 25100
rect 30380 24200 30432 24206
rect 30484 24188 30512 25230
rect 30564 24880 30616 24886
rect 30564 24822 30616 24828
rect 30576 24206 30604 24822
rect 30668 24410 30696 25298
rect 30760 25158 30788 25486
rect 30748 25152 30800 25158
rect 30748 25094 30800 25100
rect 30760 24750 30788 25094
rect 30748 24744 30800 24750
rect 30748 24686 30800 24692
rect 30656 24404 30708 24410
rect 30656 24346 30708 24352
rect 30432 24160 30512 24188
rect 30564 24200 30616 24206
rect 30380 24142 30432 24148
rect 30616 24160 30696 24188
rect 30564 24142 30616 24148
rect 30564 23656 30616 23662
rect 30564 23598 30616 23604
rect 30380 23520 30432 23526
rect 30380 23462 30432 23468
rect 30392 23186 30420 23462
rect 30380 23180 30432 23186
rect 30380 23122 30432 23128
rect 30472 23044 30524 23050
rect 30472 22986 30524 22992
rect 30196 22024 30248 22030
rect 30196 21966 30248 21972
rect 30288 22024 30340 22030
rect 30288 21966 30340 21972
rect 30300 21894 30328 21966
rect 30288 21888 30340 21894
rect 30288 21830 30340 21836
rect 30288 21412 30340 21418
rect 30288 21354 30340 21360
rect 30300 20806 30328 21354
rect 30288 20800 30340 20806
rect 30288 20742 30340 20748
rect 30300 20398 30328 20742
rect 30196 20392 30248 20398
rect 30196 20334 30248 20340
rect 30288 20392 30340 20398
rect 30288 20334 30340 20340
rect 30208 19854 30236 20334
rect 30380 20256 30432 20262
rect 30380 20198 30432 20204
rect 30392 19854 30420 20198
rect 30104 19848 30156 19854
rect 30104 19790 30156 19796
rect 30196 19848 30248 19854
rect 30196 19790 30248 19796
rect 30380 19848 30432 19854
rect 30380 19790 30432 19796
rect 30116 19310 30144 19790
rect 30484 19378 30512 22986
rect 30576 21622 30604 23598
rect 30564 21616 30616 21622
rect 30564 21558 30616 21564
rect 30668 21554 30696 24160
rect 30852 23186 30880 25638
rect 31116 25424 31168 25430
rect 31116 25366 31168 25372
rect 31128 24954 31156 25366
rect 31300 25288 31352 25294
rect 31300 25230 31352 25236
rect 31116 24948 31168 24954
rect 31116 24890 31168 24896
rect 31312 24614 31340 25230
rect 31300 24608 31352 24614
rect 31300 24550 31352 24556
rect 31300 24200 31352 24206
rect 31300 24142 31352 24148
rect 30932 24064 30984 24070
rect 30932 24006 30984 24012
rect 31116 24064 31168 24070
rect 31116 24006 31168 24012
rect 30944 23662 30972 24006
rect 30932 23656 30984 23662
rect 30932 23598 30984 23604
rect 30840 23180 30892 23186
rect 30840 23122 30892 23128
rect 31128 23118 31156 24006
rect 31312 23866 31340 24142
rect 31300 23860 31352 23866
rect 31300 23802 31352 23808
rect 31116 23112 31168 23118
rect 31116 23054 31168 23060
rect 31404 22642 31432 26930
rect 32036 26784 32088 26790
rect 32036 26726 32088 26732
rect 31852 26580 31904 26586
rect 31852 26522 31904 26528
rect 31576 25832 31628 25838
rect 31576 25774 31628 25780
rect 31588 25294 31616 25774
rect 31576 25288 31628 25294
rect 31576 25230 31628 25236
rect 31588 25158 31616 25230
rect 31576 25152 31628 25158
rect 31576 25094 31628 25100
rect 31760 25152 31812 25158
rect 31760 25094 31812 25100
rect 31576 24948 31628 24954
rect 31576 24890 31628 24896
rect 31588 24750 31616 24890
rect 31772 24818 31800 25094
rect 31760 24812 31812 24818
rect 31760 24754 31812 24760
rect 31576 24744 31628 24750
rect 31576 24686 31628 24692
rect 31484 24608 31536 24614
rect 31484 24550 31536 24556
rect 31496 24410 31524 24550
rect 31484 24404 31536 24410
rect 31484 24346 31536 24352
rect 31496 23730 31524 24346
rect 31760 24200 31812 24206
rect 31760 24142 31812 24148
rect 31484 23724 31536 23730
rect 31484 23666 31536 23672
rect 31772 23662 31800 24142
rect 31760 23656 31812 23662
rect 31760 23598 31812 23604
rect 31392 22636 31444 22642
rect 31392 22578 31444 22584
rect 30656 21548 30708 21554
rect 30656 21490 30708 21496
rect 31576 20868 31628 20874
rect 31576 20810 31628 20816
rect 31392 20800 31444 20806
rect 31392 20742 31444 20748
rect 31404 20466 31432 20742
rect 31588 20602 31616 20810
rect 31576 20596 31628 20602
rect 31576 20538 31628 20544
rect 31864 20534 31892 26522
rect 32048 26382 32076 26726
rect 32312 26512 32364 26518
rect 32312 26454 32364 26460
rect 32036 26376 32088 26382
rect 32036 26318 32088 26324
rect 32324 25906 32352 26454
rect 32508 26382 32536 27882
rect 32600 27674 32628 28018
rect 32588 27668 32640 27674
rect 32588 27610 32640 27616
rect 32600 26450 32628 27610
rect 32784 27334 32812 28086
rect 32864 28076 32916 28082
rect 32864 28018 32916 28024
rect 32772 27328 32824 27334
rect 32772 27270 32824 27276
rect 32784 26586 32812 27270
rect 32876 26994 32904 28018
rect 33244 27062 33272 28086
rect 33416 27872 33468 27878
rect 33416 27814 33468 27820
rect 33428 27470 33456 27814
rect 33416 27464 33468 27470
rect 33416 27406 33468 27412
rect 34152 27328 34204 27334
rect 34152 27270 34204 27276
rect 33232 27056 33284 27062
rect 33232 26998 33284 27004
rect 32864 26988 32916 26994
rect 32864 26930 32916 26936
rect 32772 26580 32824 26586
rect 32772 26522 32824 26528
rect 32588 26444 32640 26450
rect 32588 26386 32640 26392
rect 32496 26376 32548 26382
rect 32496 26318 32548 26324
rect 32876 26042 32904 26930
rect 33244 26586 33272 26998
rect 33784 26988 33836 26994
rect 33836 26948 33916 26976
rect 33784 26930 33836 26936
rect 33324 26920 33376 26926
rect 33324 26862 33376 26868
rect 33232 26580 33284 26586
rect 33232 26522 33284 26528
rect 33336 26042 33364 26862
rect 33888 26314 33916 26948
rect 34060 26580 34112 26586
rect 34060 26522 34112 26528
rect 33876 26308 33928 26314
rect 33876 26250 33928 26256
rect 32864 26036 32916 26042
rect 32864 25978 32916 25984
rect 33324 26036 33376 26042
rect 33324 25978 33376 25984
rect 33888 25906 33916 26250
rect 34072 25906 34100 26522
rect 34164 26382 34192 27270
rect 34716 27062 34744 29582
rect 34796 29572 34848 29578
rect 34796 29514 34848 29520
rect 34808 29306 34836 29514
rect 34796 29300 34848 29306
rect 34796 29242 34848 29248
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 35624 27872 35676 27878
rect 35624 27814 35676 27820
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 34704 27056 34756 27062
rect 34704 26998 34756 27004
rect 34716 26518 34744 26998
rect 35348 26784 35400 26790
rect 35348 26726 35400 26732
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 34704 26512 34756 26518
rect 34704 26454 34756 26460
rect 34152 26376 34204 26382
rect 34152 26318 34204 26324
rect 32312 25900 32364 25906
rect 32312 25842 32364 25848
rect 33876 25900 33928 25906
rect 33876 25842 33928 25848
rect 34060 25900 34112 25906
rect 34060 25842 34112 25848
rect 33232 25492 33284 25498
rect 33232 25434 33284 25440
rect 32404 25288 32456 25294
rect 32404 25230 32456 25236
rect 33048 25288 33100 25294
rect 33048 25230 33100 25236
rect 32312 24812 32364 24818
rect 32312 24754 32364 24760
rect 32324 24138 32352 24754
rect 32416 24750 32444 25230
rect 32772 25220 32824 25226
rect 32772 25162 32824 25168
rect 32680 25152 32732 25158
rect 32680 25094 32732 25100
rect 32404 24744 32456 24750
rect 32404 24686 32456 24692
rect 32692 24410 32720 25094
rect 32784 24750 32812 25162
rect 33060 24954 33088 25230
rect 33048 24948 33100 24954
rect 33048 24890 33100 24896
rect 33060 24750 33088 24890
rect 32772 24744 32824 24750
rect 32772 24686 32824 24692
rect 33048 24744 33100 24750
rect 33048 24686 33100 24692
rect 33244 24614 33272 25434
rect 33416 25288 33468 25294
rect 33416 25230 33468 25236
rect 33324 25152 33376 25158
rect 33324 25094 33376 25100
rect 33336 24886 33364 25094
rect 33324 24880 33376 24886
rect 33324 24822 33376 24828
rect 33232 24608 33284 24614
rect 33232 24550 33284 24556
rect 32680 24404 32732 24410
rect 32680 24346 32732 24352
rect 33244 24206 33272 24550
rect 33428 24410 33456 25230
rect 33416 24404 33468 24410
rect 33416 24346 33468 24352
rect 33232 24200 33284 24206
rect 33232 24142 33284 24148
rect 32312 24132 32364 24138
rect 32312 24074 32364 24080
rect 32220 23724 32272 23730
rect 32220 23666 32272 23672
rect 32232 23322 32260 23666
rect 32324 23662 32352 24074
rect 32312 23656 32364 23662
rect 32312 23598 32364 23604
rect 32220 23316 32272 23322
rect 32220 23258 32272 23264
rect 32404 23248 32456 23254
rect 32404 23190 32456 23196
rect 32416 22642 32444 23190
rect 32128 22636 32180 22642
rect 32128 22578 32180 22584
rect 32220 22636 32272 22642
rect 32220 22578 32272 22584
rect 32404 22636 32456 22642
rect 32404 22578 32456 22584
rect 32140 22234 32168 22578
rect 32128 22228 32180 22234
rect 32128 22170 32180 22176
rect 32232 22030 32260 22578
rect 32416 22166 32444 22578
rect 32864 22432 32916 22438
rect 32864 22374 32916 22380
rect 32404 22160 32456 22166
rect 32404 22102 32456 22108
rect 32220 22024 32272 22030
rect 32220 21966 32272 21972
rect 32312 22024 32364 22030
rect 32312 21966 32364 21972
rect 32232 21350 32260 21966
rect 32220 21344 32272 21350
rect 32220 21286 32272 21292
rect 32128 20800 32180 20806
rect 32128 20742 32180 20748
rect 32140 20602 32168 20742
rect 32232 20602 32260 21286
rect 32324 20942 32352 21966
rect 32416 21690 32444 22102
rect 32876 22030 32904 22374
rect 32864 22024 32916 22030
rect 32864 21966 32916 21972
rect 32404 21684 32456 21690
rect 32404 21626 32456 21632
rect 32588 21684 32640 21690
rect 32588 21626 32640 21632
rect 32496 21412 32548 21418
rect 32496 21354 32548 21360
rect 32404 21140 32456 21146
rect 32508 21128 32536 21354
rect 32456 21100 32536 21128
rect 32404 21082 32456 21088
rect 32312 20936 32364 20942
rect 32312 20878 32364 20884
rect 32128 20596 32180 20602
rect 32128 20538 32180 20544
rect 32220 20596 32272 20602
rect 32220 20538 32272 20544
rect 31852 20528 31904 20534
rect 31852 20470 31904 20476
rect 31392 20460 31444 20466
rect 31392 20402 31444 20408
rect 32220 20256 32272 20262
rect 32220 20198 32272 20204
rect 30656 19984 30708 19990
rect 30656 19926 30708 19932
rect 30472 19372 30524 19378
rect 30472 19314 30524 19320
rect 30104 19304 30156 19310
rect 30104 19246 30156 19252
rect 30012 18828 30064 18834
rect 30012 18770 30064 18776
rect 30484 18766 30512 19314
rect 30472 18760 30524 18766
rect 30472 18702 30524 18708
rect 29920 18692 29972 18698
rect 29920 18634 29972 18640
rect 30012 18692 30064 18698
rect 30012 18634 30064 18640
rect 29092 18624 29144 18630
rect 29092 18566 29144 18572
rect 29644 18624 29696 18630
rect 29644 18566 29696 18572
rect 29104 18358 29132 18566
rect 29092 18352 29144 18358
rect 29092 18294 29144 18300
rect 29460 18352 29512 18358
rect 29460 18294 29512 18300
rect 29472 17814 29500 18294
rect 28736 17734 28856 17762
rect 29460 17808 29512 17814
rect 29460 17750 29512 17756
rect 29368 17740 29420 17746
rect 28736 17678 28764 17734
rect 29368 17682 29420 17688
rect 28724 17672 28776 17678
rect 28724 17614 28776 17620
rect 28632 17536 28684 17542
rect 28632 17478 28684 17484
rect 29000 17536 29052 17542
rect 29000 17478 29052 17484
rect 28448 15700 28500 15706
rect 28448 15642 28500 15648
rect 27712 15496 27764 15502
rect 27712 15438 27764 15444
rect 28172 13932 28224 13938
rect 28172 13874 28224 13880
rect 27528 13796 27580 13802
rect 27528 13738 27580 13744
rect 27252 13252 27304 13258
rect 27252 13194 27304 13200
rect 27264 12850 27292 13194
rect 27540 12918 27568 13738
rect 28184 13530 28212 13874
rect 28172 13524 28224 13530
rect 28172 13466 28224 13472
rect 28356 13184 28408 13190
rect 28356 13126 28408 13132
rect 28448 13184 28500 13190
rect 28448 13126 28500 13132
rect 27528 12912 27580 12918
rect 27528 12854 27580 12860
rect 27252 12844 27304 12850
rect 27252 12786 27304 12792
rect 27160 11824 27212 11830
rect 27160 11766 27212 11772
rect 26976 11756 27028 11762
rect 26976 11698 27028 11704
rect 26056 11688 26108 11694
rect 26056 11630 26108 11636
rect 25320 11552 25372 11558
rect 25320 11494 25372 11500
rect 25332 10470 25360 11494
rect 25780 11144 25832 11150
rect 25780 11086 25832 11092
rect 25688 11008 25740 11014
rect 25688 10950 25740 10956
rect 25320 10464 25372 10470
rect 25320 10406 25372 10412
rect 25332 10062 25360 10406
rect 25320 10056 25372 10062
rect 25320 9998 25372 10004
rect 25136 9444 25188 9450
rect 25136 9386 25188 9392
rect 25228 9376 25280 9382
rect 25228 9318 25280 9324
rect 25240 8634 25268 9318
rect 25228 8628 25280 8634
rect 25228 8570 25280 8576
rect 25332 7954 25360 9998
rect 25700 9994 25728 10950
rect 25792 10810 25820 11086
rect 25780 10804 25832 10810
rect 25780 10746 25832 10752
rect 25688 9988 25740 9994
rect 25688 9930 25740 9936
rect 25792 9654 25820 10746
rect 27172 9654 27200 11766
rect 28368 10810 28396 13126
rect 28460 12986 28488 13126
rect 28448 12980 28500 12986
rect 28448 12922 28500 12928
rect 28644 12238 28672 17478
rect 29012 16046 29040 17478
rect 29380 17202 29408 17682
rect 29472 17270 29500 17750
rect 29460 17264 29512 17270
rect 29460 17206 29512 17212
rect 29368 17196 29420 17202
rect 29368 17138 29420 17144
rect 29380 16794 29408 17138
rect 29368 16788 29420 16794
rect 29368 16730 29420 16736
rect 28816 16040 28868 16046
rect 28816 15982 28868 15988
rect 29000 16040 29052 16046
rect 29000 15982 29052 15988
rect 28828 15706 28856 15982
rect 28908 15904 28960 15910
rect 28908 15846 28960 15852
rect 28816 15700 28868 15706
rect 28816 15642 28868 15648
rect 28920 13530 28948 15846
rect 29380 15570 29408 16730
rect 29368 15564 29420 15570
rect 29368 15506 29420 15512
rect 29656 15502 29684 18566
rect 29736 18080 29788 18086
rect 29736 18022 29788 18028
rect 29644 15496 29696 15502
rect 29644 15438 29696 15444
rect 29748 14346 29776 18022
rect 29932 17678 29960 18634
rect 30024 18426 30052 18634
rect 30012 18420 30064 18426
rect 30012 18362 30064 18368
rect 30104 18352 30156 18358
rect 30104 18294 30156 18300
rect 30012 17876 30064 17882
rect 30012 17818 30064 17824
rect 29920 17672 29972 17678
rect 29920 17614 29972 17620
rect 30024 17610 30052 17818
rect 30012 17604 30064 17610
rect 30012 17546 30064 17552
rect 29736 14340 29788 14346
rect 29736 14282 29788 14288
rect 29000 14272 29052 14278
rect 29000 14214 29052 14220
rect 28908 13524 28960 13530
rect 28908 13466 28960 13472
rect 28816 12844 28868 12850
rect 28816 12786 28868 12792
rect 28828 12442 28856 12786
rect 29012 12782 29040 14214
rect 30024 14006 30052 17546
rect 30116 17542 30144 18294
rect 30668 18290 30696 19926
rect 32232 19446 32260 20198
rect 32220 19440 32272 19446
rect 32220 19382 32272 19388
rect 32128 19304 32180 19310
rect 32128 19246 32180 19252
rect 30748 18624 30800 18630
rect 30748 18566 30800 18572
rect 30656 18284 30708 18290
rect 30656 18226 30708 18232
rect 30760 18222 30788 18566
rect 30748 18216 30800 18222
rect 30748 18158 30800 18164
rect 32140 18154 32168 19246
rect 32324 18766 32352 20878
rect 32508 20346 32536 21100
rect 32600 20466 32628 21626
rect 33048 21616 33100 21622
rect 33048 21558 33100 21564
rect 33060 21078 33088 21558
rect 33692 21480 33744 21486
rect 33692 21422 33744 21428
rect 33704 21146 33732 21422
rect 33692 21140 33744 21146
rect 33692 21082 33744 21088
rect 33048 21072 33100 21078
rect 33048 21014 33100 21020
rect 33060 20534 33088 21014
rect 33704 21010 33732 21082
rect 33692 21004 33744 21010
rect 33692 20946 33744 20952
rect 33048 20528 33100 20534
rect 33048 20470 33100 20476
rect 32588 20460 32640 20466
rect 32588 20402 32640 20408
rect 32508 20318 32628 20346
rect 33888 20330 33916 25842
rect 34716 24818 34744 26454
rect 35360 26382 35388 26726
rect 35348 26376 35400 26382
rect 35348 26318 35400 26324
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 34704 24812 34756 24818
rect 34704 24754 34756 24760
rect 34716 23730 34744 24754
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 34704 23724 34756 23730
rect 34704 23666 34756 23672
rect 35348 23724 35400 23730
rect 35348 23666 35400 23672
rect 34716 23186 34744 23666
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 34704 23180 34756 23186
rect 34704 23122 34756 23128
rect 34716 22710 34744 23122
rect 34888 23044 34940 23050
rect 34888 22986 34940 22992
rect 34704 22704 34756 22710
rect 34704 22646 34756 22652
rect 34520 22636 34572 22642
rect 34520 22578 34572 22584
rect 34532 21146 34560 22578
rect 34900 22522 34928 22986
rect 34716 22494 34928 22522
rect 34520 21140 34572 21146
rect 34520 21082 34572 21088
rect 34060 20800 34112 20806
rect 34060 20742 34112 20748
rect 34072 20466 34100 20742
rect 34060 20460 34112 20466
rect 34060 20402 34112 20408
rect 32600 19990 32628 20318
rect 33876 20324 33928 20330
rect 33876 20266 33928 20272
rect 32588 19984 32640 19990
rect 32588 19926 32640 19932
rect 32404 19848 32456 19854
rect 32404 19790 32456 19796
rect 32416 19514 32444 19790
rect 32496 19712 32548 19718
rect 32496 19654 32548 19660
rect 32404 19508 32456 19514
rect 32404 19450 32456 19456
rect 32508 18766 32536 19654
rect 32600 19378 32628 19926
rect 34716 19922 34744 22494
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 34796 22024 34848 22030
rect 34796 21966 34848 21972
rect 34808 21350 34836 21966
rect 35360 21962 35388 23666
rect 35532 22024 35584 22030
rect 35532 21966 35584 21972
rect 35348 21956 35400 21962
rect 35348 21898 35400 21904
rect 35544 21554 35572 21966
rect 35532 21548 35584 21554
rect 35532 21490 35584 21496
rect 34796 21344 34848 21350
rect 34796 21286 34848 21292
rect 34808 20942 34836 21286
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 34796 20936 34848 20942
rect 34796 20878 34848 20884
rect 34888 20868 34940 20874
rect 34888 20810 34940 20816
rect 34900 20602 34928 20810
rect 35348 20800 35400 20806
rect 35348 20742 35400 20748
rect 34888 20596 34940 20602
rect 34888 20538 34940 20544
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 34704 19916 34756 19922
rect 34704 19858 34756 19864
rect 33600 19848 33652 19854
rect 33600 19790 33652 19796
rect 33612 19446 33640 19790
rect 34980 19712 35032 19718
rect 34980 19654 35032 19660
rect 33600 19440 33652 19446
rect 33600 19382 33652 19388
rect 32588 19372 32640 19378
rect 32588 19314 32640 19320
rect 33612 18970 33640 19382
rect 34992 19310 35020 19654
rect 35360 19378 35388 20742
rect 35348 19372 35400 19378
rect 35348 19314 35400 19320
rect 34980 19304 35032 19310
rect 34980 19246 35032 19252
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 33600 18964 33652 18970
rect 33600 18906 33652 18912
rect 32312 18760 32364 18766
rect 32312 18702 32364 18708
rect 32496 18760 32548 18766
rect 32496 18702 32548 18708
rect 32324 18358 32352 18702
rect 32312 18352 32364 18358
rect 32312 18294 32364 18300
rect 32128 18148 32180 18154
rect 32128 18090 32180 18096
rect 31024 18080 31076 18086
rect 31024 18022 31076 18028
rect 34796 18080 34848 18086
rect 34796 18022 34848 18028
rect 31036 17678 31064 18022
rect 34808 17678 34836 18022
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 31024 17672 31076 17678
rect 31024 17614 31076 17620
rect 34796 17672 34848 17678
rect 34980 17672 35032 17678
rect 34848 17620 34928 17626
rect 34796 17614 34928 17620
rect 34980 17614 35032 17620
rect 34808 17598 34928 17614
rect 30104 17536 30156 17542
rect 30104 17478 30156 17484
rect 32588 17536 32640 17542
rect 32588 17478 32640 17484
rect 34796 17536 34848 17542
rect 34796 17478 34848 17484
rect 30116 16590 30144 17478
rect 30748 16992 30800 16998
rect 30748 16934 30800 16940
rect 30760 16590 30788 16934
rect 32600 16590 32628 17478
rect 34612 16992 34664 16998
rect 34612 16934 34664 16940
rect 32772 16720 32824 16726
rect 32772 16662 32824 16668
rect 33324 16720 33376 16726
rect 33324 16662 33376 16668
rect 30104 16584 30156 16590
rect 30104 16526 30156 16532
rect 30748 16584 30800 16590
rect 30748 16526 30800 16532
rect 31024 16584 31076 16590
rect 31024 16526 31076 16532
rect 32588 16584 32640 16590
rect 32640 16544 32720 16572
rect 32588 16526 32640 16532
rect 30760 16114 30788 16526
rect 31036 16454 31064 16526
rect 31116 16516 31168 16522
rect 31116 16458 31168 16464
rect 31024 16448 31076 16454
rect 31024 16390 31076 16396
rect 31036 16182 31064 16390
rect 31024 16176 31076 16182
rect 31024 16118 31076 16124
rect 31128 16114 31156 16458
rect 32312 16448 32364 16454
rect 32312 16390 32364 16396
rect 32588 16448 32640 16454
rect 32588 16390 32640 16396
rect 32324 16182 32352 16390
rect 32312 16176 32364 16182
rect 32312 16118 32364 16124
rect 32600 16114 32628 16390
rect 30748 16108 30800 16114
rect 30748 16050 30800 16056
rect 31116 16108 31168 16114
rect 31116 16050 31168 16056
rect 32588 16108 32640 16114
rect 32588 16050 32640 16056
rect 32600 15978 32628 16050
rect 32692 16046 32720 16544
rect 32784 16522 32812 16662
rect 32864 16584 32916 16590
rect 32864 16526 32916 16532
rect 32956 16584 33008 16590
rect 32956 16526 33008 16532
rect 32772 16516 32824 16522
rect 32772 16458 32824 16464
rect 32680 16040 32732 16046
rect 32680 15982 32732 15988
rect 32588 15972 32640 15978
rect 32588 15914 32640 15920
rect 32036 15904 32088 15910
rect 32036 15846 32088 15852
rect 30932 15360 30984 15366
rect 30932 15302 30984 15308
rect 30944 15094 30972 15302
rect 30932 15088 30984 15094
rect 30932 15030 30984 15036
rect 30196 14816 30248 14822
rect 30196 14758 30248 14764
rect 31668 14816 31720 14822
rect 31668 14758 31720 14764
rect 30012 14000 30064 14006
rect 30012 13942 30064 13948
rect 30104 13932 30156 13938
rect 30104 13874 30156 13880
rect 30116 13326 30144 13874
rect 30208 13870 30236 14758
rect 30380 14340 30432 14346
rect 30380 14282 30432 14288
rect 30288 14272 30340 14278
rect 30288 14214 30340 14220
rect 30300 13938 30328 14214
rect 30288 13932 30340 13938
rect 30288 13874 30340 13880
rect 30196 13864 30248 13870
rect 30196 13806 30248 13812
rect 30300 13394 30328 13874
rect 30288 13388 30340 13394
rect 30288 13330 30340 13336
rect 29276 13320 29328 13326
rect 29276 13262 29328 13268
rect 30104 13320 30156 13326
rect 30104 13262 30156 13268
rect 29288 12986 29316 13262
rect 30288 13252 30340 13258
rect 30288 13194 30340 13200
rect 30300 12986 30328 13194
rect 29276 12980 29328 12986
rect 29276 12922 29328 12928
rect 30288 12980 30340 12986
rect 30288 12922 30340 12928
rect 29092 12844 29144 12850
rect 29092 12786 29144 12792
rect 29000 12776 29052 12782
rect 29000 12718 29052 12724
rect 28816 12436 28868 12442
rect 28816 12378 28868 12384
rect 28632 12232 28684 12238
rect 28632 12174 28684 12180
rect 29104 11898 29132 12786
rect 30392 12714 30420 14282
rect 31680 13938 31708 14758
rect 31852 14544 31904 14550
rect 31852 14486 31904 14492
rect 31760 14408 31812 14414
rect 31760 14350 31812 14356
rect 31668 13932 31720 13938
rect 31668 13874 31720 13880
rect 31772 13870 31800 14350
rect 31864 14074 31892 14486
rect 32048 14414 32076 15846
rect 32600 15706 32628 15914
rect 32588 15700 32640 15706
rect 32588 15642 32640 15648
rect 32876 15502 32904 16526
rect 32968 16182 32996 16526
rect 32956 16176 33008 16182
rect 32956 16118 33008 16124
rect 32968 15570 32996 16118
rect 32956 15564 33008 15570
rect 32956 15506 33008 15512
rect 33336 15502 33364 16662
rect 34624 16522 34652 16934
rect 34808 16658 34836 17478
rect 34900 17202 34928 17598
rect 34992 17270 35020 17614
rect 34980 17264 35032 17270
rect 34980 17206 35032 17212
rect 34888 17196 34940 17202
rect 34888 17138 34940 17144
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 34796 16652 34848 16658
rect 34796 16594 34848 16600
rect 34612 16516 34664 16522
rect 34612 16458 34664 16464
rect 35348 16516 35400 16522
rect 35348 16458 35400 16464
rect 34704 16448 34756 16454
rect 34704 16390 34756 16396
rect 34796 16448 34848 16454
rect 34796 16390 34848 16396
rect 34716 16114 34744 16390
rect 33692 16108 33744 16114
rect 33692 16050 33744 16056
rect 34704 16108 34756 16114
rect 34704 16050 34756 16056
rect 33704 15706 33732 16050
rect 34612 15904 34664 15910
rect 34612 15846 34664 15852
rect 33692 15700 33744 15706
rect 33692 15642 33744 15648
rect 32864 15496 32916 15502
rect 32864 15438 32916 15444
rect 33324 15496 33376 15502
rect 33324 15438 33376 15444
rect 34520 14612 34572 14618
rect 34440 14572 34520 14600
rect 32036 14408 32088 14414
rect 32036 14350 32088 14356
rect 32220 14408 32272 14414
rect 32220 14350 32272 14356
rect 33600 14408 33652 14414
rect 33600 14350 33652 14356
rect 33784 14408 33836 14414
rect 33784 14350 33836 14356
rect 32232 14074 32260 14350
rect 33416 14272 33468 14278
rect 33416 14214 33468 14220
rect 31852 14068 31904 14074
rect 31852 14010 31904 14016
rect 32220 14068 32272 14074
rect 32220 14010 32272 14016
rect 33232 13932 33284 13938
rect 33232 13874 33284 13880
rect 31760 13864 31812 13870
rect 31760 13806 31812 13812
rect 33048 13796 33100 13802
rect 33048 13738 33100 13744
rect 30748 13728 30800 13734
rect 30748 13670 30800 13676
rect 31024 13728 31076 13734
rect 31024 13670 31076 13676
rect 32864 13728 32916 13734
rect 32864 13670 32916 13676
rect 30760 12850 30788 13670
rect 31036 13326 31064 13670
rect 31024 13320 31076 13326
rect 31024 13262 31076 13268
rect 32220 13320 32272 13326
rect 32220 13262 32272 13268
rect 30748 12844 30800 12850
rect 30748 12786 30800 12792
rect 31036 12782 31064 13262
rect 32232 12986 32260 13262
rect 32312 13184 32364 13190
rect 32312 13126 32364 13132
rect 32220 12980 32272 12986
rect 32220 12922 32272 12928
rect 31208 12844 31260 12850
rect 31484 12844 31536 12850
rect 31260 12804 31484 12832
rect 31208 12786 31260 12792
rect 31484 12786 31536 12792
rect 31024 12776 31076 12782
rect 31024 12718 31076 12724
rect 30380 12708 30432 12714
rect 30380 12650 30432 12656
rect 30840 12708 30892 12714
rect 30840 12650 30892 12656
rect 30472 12640 30524 12646
rect 30472 12582 30524 12588
rect 30484 12238 30512 12582
rect 30472 12232 30524 12238
rect 30472 12174 30524 12180
rect 29092 11892 29144 11898
rect 29092 11834 29144 11840
rect 30472 11552 30524 11558
rect 30472 11494 30524 11500
rect 28356 10804 28408 10810
rect 28356 10746 28408 10752
rect 30484 10742 30512 11494
rect 30288 10736 30340 10742
rect 30288 10678 30340 10684
rect 30472 10736 30524 10742
rect 30472 10678 30524 10684
rect 29920 10668 29972 10674
rect 29920 10610 29972 10616
rect 28908 10600 28960 10606
rect 28908 10542 28960 10548
rect 27344 10056 27396 10062
rect 27344 9998 27396 10004
rect 25780 9648 25832 9654
rect 25780 9590 25832 9596
rect 27160 9648 27212 9654
rect 27160 9590 27212 9596
rect 25504 9580 25556 9586
rect 25504 9522 25556 9528
rect 25516 8974 25544 9522
rect 26240 9512 26292 9518
rect 26240 9454 26292 9460
rect 25504 8968 25556 8974
rect 25504 8910 25556 8916
rect 25320 7948 25372 7954
rect 25320 7890 25372 7896
rect 25516 7410 25544 8910
rect 26252 8906 26280 9454
rect 26240 8900 26292 8906
rect 26240 8842 26292 8848
rect 27160 8832 27212 8838
rect 27160 8774 27212 8780
rect 27172 8566 27200 8774
rect 27160 8560 27212 8566
rect 27160 8502 27212 8508
rect 27356 8498 27384 9998
rect 27620 9988 27672 9994
rect 27620 9930 27672 9936
rect 27632 9450 27660 9930
rect 28920 9722 28948 10542
rect 29552 9920 29604 9926
rect 29552 9862 29604 9868
rect 28908 9716 28960 9722
rect 28908 9658 28960 9664
rect 29184 9580 29236 9586
rect 29184 9522 29236 9528
rect 27620 9444 27672 9450
rect 27620 9386 27672 9392
rect 29196 9178 29224 9522
rect 29184 9172 29236 9178
rect 29184 9114 29236 9120
rect 29564 8974 29592 9862
rect 29932 9722 29960 10610
rect 29920 9716 29972 9722
rect 29920 9658 29972 9664
rect 28632 8968 28684 8974
rect 28632 8910 28684 8916
rect 29552 8968 29604 8974
rect 29552 8910 29604 8916
rect 28644 8634 28672 8910
rect 29184 8832 29236 8838
rect 29184 8774 29236 8780
rect 28632 8628 28684 8634
rect 28632 8570 28684 8576
rect 29196 8498 29224 8774
rect 27344 8492 27396 8498
rect 27344 8434 27396 8440
rect 29184 8492 29236 8498
rect 29184 8434 29236 8440
rect 30300 8430 30328 10678
rect 30852 10674 30880 12650
rect 32324 12238 32352 13126
rect 32876 12238 32904 13670
rect 33060 13462 33088 13738
rect 33048 13456 33100 13462
rect 33048 13398 33100 13404
rect 32312 12232 32364 12238
rect 32312 12174 32364 12180
rect 32864 12232 32916 12238
rect 32864 12174 32916 12180
rect 31944 12096 31996 12102
rect 31944 12038 31996 12044
rect 31956 11762 31984 12038
rect 33060 11762 33088 13398
rect 33244 12986 33272 13874
rect 33428 13394 33456 14214
rect 33612 14006 33640 14350
rect 33600 14000 33652 14006
rect 33600 13942 33652 13948
rect 33416 13388 33468 13394
rect 33416 13330 33468 13336
rect 33232 12980 33284 12986
rect 33232 12922 33284 12928
rect 33612 12306 33640 13942
rect 33796 12986 33824 14350
rect 34440 13938 34468 14572
rect 34520 14554 34572 14560
rect 34624 14414 34652 15846
rect 34716 15570 34744 16050
rect 34808 15638 34836 16390
rect 35360 16046 35388 16458
rect 35348 16040 35400 16046
rect 35348 15982 35400 15988
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 34796 15632 34848 15638
rect 34796 15574 34848 15580
rect 35532 15632 35584 15638
rect 35532 15574 35584 15580
rect 34704 15564 34756 15570
rect 34704 15506 34756 15512
rect 34716 15026 34744 15506
rect 35348 15360 35400 15366
rect 35348 15302 35400 15308
rect 34704 15020 34756 15026
rect 34704 14962 34756 14968
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 34612 14408 34664 14414
rect 34612 14350 34664 14356
rect 35360 14346 35388 15302
rect 35544 15026 35572 15574
rect 35532 15020 35584 15026
rect 35532 14962 35584 14968
rect 35532 14612 35584 14618
rect 35532 14554 35584 14560
rect 35544 14346 35572 14554
rect 34520 14340 34572 14346
rect 34520 14282 34572 14288
rect 35348 14340 35400 14346
rect 35348 14282 35400 14288
rect 35532 14340 35584 14346
rect 35532 14282 35584 14288
rect 34428 13932 34480 13938
rect 34428 13874 34480 13880
rect 34336 13728 34388 13734
rect 34336 13670 34388 13676
rect 34348 13326 34376 13670
rect 34532 13326 34560 14282
rect 34704 14272 34756 14278
rect 34704 14214 34756 14220
rect 34980 14272 35032 14278
rect 34980 14214 35032 14220
rect 34612 13796 34664 13802
rect 34612 13738 34664 13744
rect 34336 13320 34388 13326
rect 34336 13262 34388 13268
rect 34520 13320 34572 13326
rect 34520 13262 34572 13268
rect 33784 12980 33836 12986
rect 33784 12922 33836 12928
rect 34532 12306 34560 13262
rect 33416 12300 33468 12306
rect 33416 12242 33468 12248
rect 33600 12300 33652 12306
rect 33600 12242 33652 12248
rect 34520 12300 34572 12306
rect 34520 12242 34572 12248
rect 31944 11756 31996 11762
rect 31944 11698 31996 11704
rect 33048 11756 33100 11762
rect 33048 11698 33100 11704
rect 30840 10668 30892 10674
rect 30840 10610 30892 10616
rect 32588 10668 32640 10674
rect 32588 10610 32640 10616
rect 30564 10464 30616 10470
rect 30564 10406 30616 10412
rect 30380 9920 30432 9926
rect 30380 9862 30432 9868
rect 30392 9586 30420 9862
rect 30576 9722 30604 10406
rect 30852 10062 30880 10610
rect 31116 10464 31168 10470
rect 31116 10406 31168 10412
rect 32312 10464 32364 10470
rect 32312 10406 32364 10412
rect 30840 10056 30892 10062
rect 30840 9998 30892 10004
rect 30564 9716 30616 9722
rect 30564 9658 30616 9664
rect 30852 9654 30880 9998
rect 31128 9994 31156 10406
rect 31484 10056 31536 10062
rect 31484 9998 31536 10004
rect 31116 9988 31168 9994
rect 31116 9930 31168 9936
rect 30840 9648 30892 9654
rect 30840 9590 30892 9596
rect 30380 9580 30432 9586
rect 30380 9522 30432 9528
rect 30564 9512 30616 9518
rect 30564 9454 30616 9460
rect 30576 8634 30604 9454
rect 30564 8628 30616 8634
rect 30564 8570 30616 8576
rect 30852 8566 30880 9590
rect 31496 9042 31524 9998
rect 32324 9586 32352 10406
rect 32600 10266 32628 10610
rect 33060 10606 33088 11698
rect 33232 11552 33284 11558
rect 33232 11494 33284 11500
rect 33048 10600 33100 10606
rect 33048 10542 33100 10548
rect 33048 10464 33100 10470
rect 33048 10406 33100 10412
rect 32588 10260 32640 10266
rect 32588 10202 32640 10208
rect 33060 10130 33088 10406
rect 33048 10124 33100 10130
rect 33048 10066 33100 10072
rect 33244 10062 33272 11494
rect 33428 11014 33456 12242
rect 33508 12096 33560 12102
rect 33508 12038 33560 12044
rect 33520 11150 33548 12038
rect 33612 11830 33640 12242
rect 33600 11824 33652 11830
rect 33600 11766 33652 11772
rect 34428 11824 34480 11830
rect 34428 11766 34480 11772
rect 33692 11756 33744 11762
rect 33692 11698 33744 11704
rect 33704 11218 33732 11698
rect 34336 11552 34388 11558
rect 34336 11494 34388 11500
rect 33692 11212 33744 11218
rect 33692 11154 33744 11160
rect 33508 11144 33560 11150
rect 33508 11086 33560 11092
rect 33324 11008 33376 11014
rect 33324 10950 33376 10956
rect 33416 11008 33468 11014
rect 33416 10950 33468 10956
rect 33336 10810 33364 10950
rect 33324 10804 33376 10810
rect 33324 10746 33376 10752
rect 33324 10668 33376 10674
rect 33324 10610 33376 10616
rect 33232 10056 33284 10062
rect 33232 9998 33284 10004
rect 33336 9654 33364 10610
rect 33428 10130 33456 10950
rect 33416 10124 33468 10130
rect 33416 10066 33468 10072
rect 33324 9648 33376 9654
rect 33324 9590 33376 9596
rect 32312 9580 32364 9586
rect 32312 9522 32364 9528
rect 33428 9518 33456 10066
rect 34348 9586 34376 11494
rect 34440 11150 34468 11766
rect 34624 11762 34652 13738
rect 34716 12986 34744 14214
rect 34796 13932 34848 13938
rect 34796 13874 34848 13880
rect 34808 13530 34836 13874
rect 34992 13870 35020 14214
rect 34980 13864 35032 13870
rect 34980 13806 35032 13812
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 34796 13524 34848 13530
rect 34796 13466 34848 13472
rect 35360 13258 35388 14282
rect 35348 13252 35400 13258
rect 35348 13194 35400 13200
rect 35532 13252 35584 13258
rect 35532 13194 35584 13200
rect 35256 13184 35308 13190
rect 35256 13126 35308 13132
rect 34704 12980 34756 12986
rect 34704 12922 34756 12928
rect 34716 12442 34744 12922
rect 34796 12844 34848 12850
rect 34796 12786 34848 12792
rect 34704 12436 34756 12442
rect 34704 12378 34756 12384
rect 34808 12306 34836 12786
rect 35268 12782 35296 13126
rect 35544 12782 35572 13194
rect 35256 12776 35308 12782
rect 35256 12718 35308 12724
rect 35532 12776 35584 12782
rect 35532 12718 35584 12724
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 35636 12434 35664 27814
rect 36004 22094 36032 37182
rect 36084 36100 36136 36106
rect 36084 36042 36136 36048
rect 36096 35494 36124 36042
rect 36084 35488 36136 35494
rect 36084 35430 36136 35436
rect 36268 34400 36320 34406
rect 36268 34342 36320 34348
rect 36280 34066 36308 34342
rect 36268 34060 36320 34066
rect 36268 34002 36320 34008
rect 36372 32842 36400 37674
rect 36464 37262 36492 37742
rect 36452 37256 36504 37262
rect 36452 37198 36504 37204
rect 36464 36854 36492 37198
rect 36544 37188 36596 37194
rect 36544 37130 36596 37136
rect 36556 36922 36584 37130
rect 36924 37126 36952 37810
rect 37568 37330 37596 37810
rect 38108 37800 38160 37806
rect 38108 37742 38160 37748
rect 37556 37324 37608 37330
rect 37556 37266 37608 37272
rect 36636 37120 36688 37126
rect 36636 37062 36688 37068
rect 36912 37120 36964 37126
rect 36912 37062 36964 37068
rect 36544 36916 36596 36922
rect 36544 36858 36596 36864
rect 36452 36848 36504 36854
rect 36452 36790 36504 36796
rect 36556 36174 36584 36858
rect 36648 36174 36676 37062
rect 37568 36922 37596 37266
rect 37832 37120 37884 37126
rect 37832 37062 37884 37068
rect 37556 36916 37608 36922
rect 37556 36858 37608 36864
rect 36820 36848 36872 36854
rect 36820 36790 36872 36796
rect 36832 36174 36860 36790
rect 36544 36168 36596 36174
rect 36544 36110 36596 36116
rect 36636 36168 36688 36174
rect 36636 36110 36688 36116
rect 36820 36168 36872 36174
rect 36820 36110 36872 36116
rect 37556 35012 37608 35018
rect 37556 34954 37608 34960
rect 36820 34944 36872 34950
rect 36820 34886 36872 34892
rect 37280 34944 37332 34950
rect 37280 34886 37332 34892
rect 36832 34678 36860 34886
rect 36820 34672 36872 34678
rect 36820 34614 36872 34620
rect 36832 33998 36860 34614
rect 37292 34082 37320 34886
rect 37568 34202 37596 34954
rect 37556 34196 37608 34202
rect 37556 34138 37608 34144
rect 37200 34066 37320 34082
rect 37188 34060 37320 34066
rect 37240 34054 37320 34060
rect 37188 34002 37240 34008
rect 36820 33992 36872 33998
rect 36820 33934 36872 33940
rect 37844 32978 37872 37062
rect 38016 35216 38068 35222
rect 38016 35158 38068 35164
rect 38028 34746 38056 35158
rect 38120 35154 38148 37742
rect 38672 36802 38700 37810
rect 38752 37664 38804 37670
rect 38752 37606 38804 37612
rect 38764 37398 38792 37606
rect 38752 37392 38804 37398
rect 38752 37334 38804 37340
rect 38764 36922 38792 37334
rect 38752 36916 38804 36922
rect 38752 36858 38804 36864
rect 38856 36854 38884 37946
rect 38948 37738 38976 38286
rect 39120 38004 39172 38010
rect 39120 37946 39172 37952
rect 39132 37874 39160 37946
rect 39120 37868 39172 37874
rect 39120 37810 39172 37816
rect 39132 37754 39160 37810
rect 38936 37732 38988 37738
rect 39132 37726 39252 37754
rect 38936 37674 38988 37680
rect 38844 36848 38896 36854
rect 38292 36780 38344 36786
rect 38672 36774 38792 36802
rect 38844 36790 38896 36796
rect 38292 36722 38344 36728
rect 38304 35630 38332 36722
rect 38476 36236 38528 36242
rect 38476 36178 38528 36184
rect 38292 35624 38344 35630
rect 38292 35566 38344 35572
rect 38108 35148 38160 35154
rect 38108 35090 38160 35096
rect 38120 34950 38148 35090
rect 38108 34944 38160 34950
rect 38108 34886 38160 34892
rect 38016 34740 38068 34746
rect 38016 34682 38068 34688
rect 38028 33998 38056 34682
rect 38304 34202 38332 35566
rect 38488 35494 38516 36178
rect 38764 36174 38792 36774
rect 38856 36650 38884 36790
rect 38844 36644 38896 36650
rect 38844 36586 38896 36592
rect 38844 36372 38896 36378
rect 38844 36314 38896 36320
rect 38752 36168 38804 36174
rect 38856 36122 38884 36314
rect 38804 36116 38884 36122
rect 38752 36110 38884 36116
rect 38764 36094 38884 36110
rect 38856 35630 38884 36094
rect 38948 35630 38976 37674
rect 39028 37664 39080 37670
rect 39028 37606 39080 37612
rect 39120 37664 39172 37670
rect 39120 37606 39172 37612
rect 39040 36242 39068 37606
rect 39132 37194 39160 37606
rect 39224 37262 39252 37726
rect 39304 37460 39356 37466
rect 39304 37402 39356 37408
rect 39212 37256 39264 37262
rect 39212 37198 39264 37204
rect 39120 37188 39172 37194
rect 39120 37130 39172 37136
rect 39120 36848 39172 36854
rect 39120 36790 39172 36796
rect 39028 36236 39080 36242
rect 39028 36178 39080 36184
rect 39132 36174 39160 36790
rect 39224 36786 39252 37198
rect 39212 36780 39264 36786
rect 39212 36722 39264 36728
rect 39224 36582 39252 36722
rect 39212 36576 39264 36582
rect 39212 36518 39264 36524
rect 39120 36168 39172 36174
rect 39120 36110 39172 36116
rect 38844 35624 38896 35630
rect 38844 35566 38896 35572
rect 38936 35624 38988 35630
rect 38936 35566 38988 35572
rect 38476 35488 38528 35494
rect 38476 35430 38528 35436
rect 38488 34678 38516 35430
rect 38856 35086 38884 35566
rect 38948 35154 38976 35566
rect 38936 35148 38988 35154
rect 38936 35090 38988 35096
rect 38752 35080 38804 35086
rect 38752 35022 38804 35028
rect 38844 35080 38896 35086
rect 38844 35022 38896 35028
rect 38476 34672 38528 34678
rect 38476 34614 38528 34620
rect 38384 34604 38436 34610
rect 38384 34546 38436 34552
rect 38292 34196 38344 34202
rect 38292 34138 38344 34144
rect 38016 33992 38068 33998
rect 38016 33934 38068 33940
rect 38396 33844 38424 34546
rect 38764 34542 38792 35022
rect 38844 34604 38896 34610
rect 38844 34546 38896 34552
rect 38752 34536 38804 34542
rect 38752 34478 38804 34484
rect 38660 34400 38712 34406
rect 38660 34342 38712 34348
rect 38672 33998 38700 34342
rect 38660 33992 38712 33998
rect 38660 33934 38712 33940
rect 38764 33930 38792 34478
rect 38856 34134 38884 34546
rect 38844 34128 38896 34134
rect 38844 34070 38896 34076
rect 38948 34066 38976 35090
rect 39212 34740 39264 34746
rect 39212 34682 39264 34688
rect 38936 34060 38988 34066
rect 38936 34002 38988 34008
rect 38752 33924 38804 33930
rect 38752 33866 38804 33872
rect 38476 33856 38528 33862
rect 38396 33816 38476 33844
rect 38476 33798 38528 33804
rect 38384 33448 38436 33454
rect 38384 33390 38436 33396
rect 38292 33312 38344 33318
rect 38292 33254 38344 33260
rect 37832 32972 37884 32978
rect 37832 32914 37884 32920
rect 37004 32904 37056 32910
rect 37004 32846 37056 32852
rect 38200 32904 38252 32910
rect 38200 32846 38252 32852
rect 36360 32836 36412 32842
rect 36360 32778 36412 32784
rect 36452 32836 36504 32842
rect 36452 32778 36504 32784
rect 36728 32836 36780 32842
rect 36728 32778 36780 32784
rect 36372 32366 36400 32778
rect 36464 32570 36492 32778
rect 36636 32768 36688 32774
rect 36636 32710 36688 32716
rect 36648 32570 36676 32710
rect 36452 32564 36504 32570
rect 36452 32506 36504 32512
rect 36636 32564 36688 32570
rect 36636 32506 36688 32512
rect 36740 32434 36768 32778
rect 36728 32428 36780 32434
rect 36728 32370 36780 32376
rect 36360 32360 36412 32366
rect 36360 32302 36412 32308
rect 37016 32230 37044 32846
rect 37924 32836 37976 32842
rect 37924 32778 37976 32784
rect 37004 32224 37056 32230
rect 37004 32166 37056 32172
rect 37016 31822 37044 32166
rect 37936 31890 37964 32778
rect 37924 31884 37976 31890
rect 37924 31826 37976 31832
rect 37004 31816 37056 31822
rect 37004 31758 37056 31764
rect 37280 31816 37332 31822
rect 37280 31758 37332 31764
rect 37016 30734 37044 31758
rect 37292 31414 37320 31758
rect 37280 31408 37332 31414
rect 37280 31350 37332 31356
rect 37936 31346 37964 31826
rect 37924 31340 37976 31346
rect 38212 31328 38240 32846
rect 38304 31482 38332 33254
rect 38396 33114 38424 33390
rect 38488 33386 38516 33798
rect 39028 33584 39080 33590
rect 39028 33526 39080 33532
rect 38936 33516 38988 33522
rect 38936 33458 38988 33464
rect 38476 33380 38528 33386
rect 38476 33322 38528 33328
rect 38384 33108 38436 33114
rect 38384 33050 38436 33056
rect 38488 31482 38516 33322
rect 38660 32904 38712 32910
rect 38660 32846 38712 32852
rect 38672 32570 38700 32846
rect 38660 32564 38712 32570
rect 38660 32506 38712 32512
rect 38672 31890 38700 32506
rect 38948 32366 38976 33458
rect 38936 32360 38988 32366
rect 38936 32302 38988 32308
rect 38660 31884 38712 31890
rect 38660 31826 38712 31832
rect 39040 31482 39068 33526
rect 39120 32768 39172 32774
rect 39120 32710 39172 32716
rect 39132 32434 39160 32710
rect 39120 32428 39172 32434
rect 39120 32370 39172 32376
rect 39224 32230 39252 34682
rect 39316 33318 39344 37402
rect 39396 36848 39448 36854
rect 39396 36790 39448 36796
rect 39408 36378 39436 36790
rect 39396 36372 39448 36378
rect 39396 36314 39448 36320
rect 39394 35456 39450 35465
rect 39394 35391 39450 35400
rect 39304 33312 39356 33318
rect 39304 33254 39356 33260
rect 39212 32224 39264 32230
rect 39212 32166 39264 32172
rect 38292 31476 38344 31482
rect 38292 31418 38344 31424
rect 38476 31476 38528 31482
rect 38476 31418 38528 31424
rect 39028 31476 39080 31482
rect 39028 31418 39080 31424
rect 38292 31340 38344 31346
rect 38212 31300 38292 31328
rect 37924 31282 37976 31288
rect 38292 31282 38344 31288
rect 37936 30802 37964 31282
rect 37924 30796 37976 30802
rect 37924 30738 37976 30744
rect 38304 30734 38332 31282
rect 38568 30932 38620 30938
rect 38568 30874 38620 30880
rect 39120 30932 39172 30938
rect 39120 30874 39172 30880
rect 37004 30728 37056 30734
rect 37004 30670 37056 30676
rect 38292 30728 38344 30734
rect 38580 30716 38608 30874
rect 38344 30688 38608 30716
rect 38292 30670 38344 30676
rect 36452 30592 36504 30598
rect 36452 30534 36504 30540
rect 37924 30592 37976 30598
rect 37924 30534 37976 30540
rect 36464 30258 36492 30534
rect 36452 30252 36504 30258
rect 36452 30194 36504 30200
rect 37832 30252 37884 30258
rect 37832 30194 37884 30200
rect 37740 30048 37792 30054
rect 37740 29990 37792 29996
rect 37752 29850 37780 29990
rect 37740 29844 37792 29850
rect 37740 29786 37792 29792
rect 37556 29504 37608 29510
rect 37556 29446 37608 29452
rect 37568 29170 37596 29446
rect 37844 29306 37872 30194
rect 37936 29578 37964 30534
rect 38580 30122 38608 30688
rect 38568 30116 38620 30122
rect 38568 30058 38620 30064
rect 39132 29782 39160 30874
rect 39120 29776 39172 29782
rect 39120 29718 39172 29724
rect 39132 29646 39160 29718
rect 39120 29640 39172 29646
rect 39120 29582 39172 29588
rect 37924 29572 37976 29578
rect 37924 29514 37976 29520
rect 37832 29300 37884 29306
rect 37832 29242 37884 29248
rect 37556 29164 37608 29170
rect 37556 29106 37608 29112
rect 36360 24812 36412 24818
rect 36360 24754 36412 24760
rect 39304 24812 39356 24818
rect 39304 24754 39356 24760
rect 36372 24410 36400 24754
rect 36360 24404 36412 24410
rect 36360 24346 36412 24352
rect 37556 24336 37608 24342
rect 37554 24304 37556 24313
rect 37608 24304 37610 24313
rect 37554 24239 37610 24248
rect 38660 24200 38712 24206
rect 38660 24142 38712 24148
rect 39120 24200 39172 24206
rect 39120 24142 39172 24148
rect 38016 23724 38068 23730
rect 38016 23666 38068 23672
rect 37096 23044 37148 23050
rect 37096 22986 37148 22992
rect 35912 22066 36032 22094
rect 37108 22094 37136 22986
rect 37108 22066 37228 22094
rect 35716 21956 35768 21962
rect 35716 21898 35768 21904
rect 35728 21554 35756 21898
rect 35716 21548 35768 21554
rect 35716 21490 35768 21496
rect 35912 20398 35940 22066
rect 36360 21888 36412 21894
rect 36360 21830 36412 21836
rect 36372 21554 36400 21830
rect 36360 21548 36412 21554
rect 36360 21490 36412 21496
rect 36176 21344 36228 21350
rect 36176 21286 36228 21292
rect 36188 20466 36216 21286
rect 36372 21010 36400 21490
rect 37200 21146 37228 22066
rect 37280 21480 37332 21486
rect 37280 21422 37332 21428
rect 37188 21140 37240 21146
rect 37188 21082 37240 21088
rect 36360 21004 36412 21010
rect 36360 20946 36412 20952
rect 37188 21004 37240 21010
rect 37188 20946 37240 20952
rect 36268 20936 36320 20942
rect 36268 20878 36320 20884
rect 36912 20936 36964 20942
rect 36912 20878 36964 20884
rect 36280 20534 36308 20878
rect 36820 20868 36872 20874
rect 36820 20810 36872 20816
rect 36268 20528 36320 20534
rect 36268 20470 36320 20476
rect 36176 20460 36228 20466
rect 36176 20402 36228 20408
rect 35900 20392 35952 20398
rect 35900 20334 35952 20340
rect 35912 19786 35940 20334
rect 36188 20330 36216 20402
rect 36176 20324 36228 20330
rect 36176 20266 36228 20272
rect 36832 19854 36860 20810
rect 36924 20466 36952 20878
rect 37200 20534 37228 20946
rect 37188 20528 37240 20534
rect 37188 20470 37240 20476
rect 36912 20460 36964 20466
rect 36912 20402 36964 20408
rect 37096 20460 37148 20466
rect 37096 20402 37148 20408
rect 37108 19922 37136 20402
rect 37096 19916 37148 19922
rect 37096 19858 37148 19864
rect 36820 19848 36872 19854
rect 36820 19790 36872 19796
rect 37108 19786 37136 19858
rect 37200 19854 37228 20470
rect 37292 20262 37320 21422
rect 38028 21146 38056 23666
rect 38672 23322 38700 24142
rect 39028 23520 39080 23526
rect 39028 23462 39080 23468
rect 38660 23316 38712 23322
rect 38660 23258 38712 23264
rect 38936 23112 38988 23118
rect 38936 23054 38988 23060
rect 38844 22636 38896 22642
rect 38844 22578 38896 22584
rect 38856 21690 38884 22578
rect 38948 22098 38976 23054
rect 38936 22092 38988 22098
rect 38936 22034 38988 22040
rect 38844 21684 38896 21690
rect 38844 21626 38896 21632
rect 38948 21570 38976 22034
rect 39040 22030 39068 23462
rect 39028 22024 39080 22030
rect 39028 21966 39080 21972
rect 38764 21542 38976 21570
rect 38476 21412 38528 21418
rect 38476 21354 38528 21360
rect 38016 21140 38068 21146
rect 38016 21082 38068 21088
rect 37924 20936 37976 20942
rect 37924 20878 37976 20884
rect 37832 20868 37884 20874
rect 37832 20810 37884 20816
rect 37844 20466 37872 20810
rect 37832 20460 37884 20466
rect 37832 20402 37884 20408
rect 37556 20392 37608 20398
rect 37556 20334 37608 20340
rect 37280 20256 37332 20262
rect 37280 20198 37332 20204
rect 37292 19990 37320 20198
rect 37280 19984 37332 19990
rect 37280 19926 37332 19932
rect 37188 19848 37240 19854
rect 37188 19790 37240 19796
rect 35900 19780 35952 19786
rect 35900 19722 35952 19728
rect 37096 19780 37148 19786
rect 37096 19722 37148 19728
rect 36636 19712 36688 19718
rect 36636 19654 36688 19660
rect 36360 18284 36412 18290
rect 36360 18226 36412 18232
rect 36372 17746 36400 18226
rect 36360 17740 36412 17746
rect 36360 17682 36412 17688
rect 36648 17678 36676 19654
rect 37200 19514 37228 19790
rect 37188 19508 37240 19514
rect 37188 19450 37240 19456
rect 37568 18290 37596 20334
rect 37936 19854 37964 20878
rect 38488 19854 38516 21354
rect 38764 21010 38792 21542
rect 38752 21004 38804 21010
rect 38752 20946 38804 20952
rect 37924 19848 37976 19854
rect 37924 19790 37976 19796
rect 38476 19848 38528 19854
rect 38476 19790 38528 19796
rect 38016 19712 38068 19718
rect 38016 19654 38068 19660
rect 38028 18358 38056 19654
rect 38488 19378 38516 19790
rect 38476 19372 38528 19378
rect 38476 19314 38528 19320
rect 38016 18352 38068 18358
rect 38016 18294 38068 18300
rect 37556 18284 37608 18290
rect 37556 18226 37608 18232
rect 38764 17678 38792 20946
rect 39132 20058 39160 24142
rect 39316 22098 39344 24754
rect 39408 23254 39436 35391
rect 39672 33108 39724 33114
rect 39672 33050 39724 33056
rect 39488 33040 39540 33046
rect 39488 32982 39540 32988
rect 39500 32570 39528 32982
rect 39488 32564 39540 32570
rect 39488 32506 39540 32512
rect 39488 32360 39540 32366
rect 39488 32302 39540 32308
rect 39500 31482 39528 32302
rect 39684 32230 39712 33050
rect 39672 32224 39724 32230
rect 39672 32166 39724 32172
rect 39488 31476 39540 31482
rect 39488 31418 39540 31424
rect 39500 30002 39528 31418
rect 39684 31414 39712 32166
rect 39672 31408 39724 31414
rect 39672 31350 39724 31356
rect 39580 31340 39632 31346
rect 39580 31282 39632 31288
rect 39592 30938 39620 31282
rect 39580 30932 39632 30938
rect 39580 30874 39632 30880
rect 39672 30252 39724 30258
rect 39672 30194 39724 30200
rect 39580 30048 39632 30054
rect 39500 29996 39580 30002
rect 39500 29990 39632 29996
rect 39500 29974 39620 29990
rect 39500 29578 39528 29974
rect 39684 29850 39712 30194
rect 39672 29844 39724 29850
rect 39672 29786 39724 29792
rect 39488 29572 39540 29578
rect 39488 29514 39540 29520
rect 39396 23248 39448 23254
rect 39396 23190 39448 23196
rect 39580 22976 39632 22982
rect 39580 22918 39632 22924
rect 39304 22092 39356 22098
rect 39304 22034 39356 22040
rect 39304 21480 39356 21486
rect 39304 21422 39356 21428
rect 39316 21146 39344 21422
rect 39304 21140 39356 21146
rect 39304 21082 39356 21088
rect 39592 20505 39620 22918
rect 39672 22024 39724 22030
rect 39672 21966 39724 21972
rect 39684 21554 39712 21966
rect 39672 21548 39724 21554
rect 39672 21490 39724 21496
rect 39578 20496 39634 20505
rect 39578 20431 39634 20440
rect 39120 20052 39172 20058
rect 39120 19994 39172 20000
rect 38936 18760 38988 18766
rect 38936 18702 38988 18708
rect 39028 18760 39080 18766
rect 39028 18702 39080 18708
rect 39580 18760 39632 18766
rect 39580 18702 39632 18708
rect 38948 18426 38976 18702
rect 38936 18420 38988 18426
rect 38936 18362 38988 18368
rect 39040 17746 39068 18702
rect 39396 18624 39448 18630
rect 39396 18566 39448 18572
rect 39408 18290 39436 18566
rect 39592 18426 39620 18702
rect 39580 18420 39632 18426
rect 39580 18362 39632 18368
rect 39396 18284 39448 18290
rect 39396 18226 39448 18232
rect 39028 17740 39080 17746
rect 39028 17682 39080 17688
rect 39776 17678 39804 39034
rect 40236 39030 40264 39238
rect 40224 39024 40276 39030
rect 40224 38966 40276 38972
rect 40040 37868 40092 37874
rect 40040 37810 40092 37816
rect 40052 37466 40080 37810
rect 40040 37460 40092 37466
rect 40040 37402 40092 37408
rect 39948 36304 40000 36310
rect 39948 36246 40000 36252
rect 39960 35766 39988 36246
rect 39948 35760 40000 35766
rect 39948 35702 40000 35708
rect 40132 35216 40184 35222
rect 40132 35158 40184 35164
rect 39856 34060 39908 34066
rect 39856 34002 39908 34008
rect 39868 32434 39896 34002
rect 40144 33998 40172 35158
rect 40224 34944 40276 34950
rect 40224 34886 40276 34892
rect 40236 34678 40264 34886
rect 40224 34672 40276 34678
rect 40224 34614 40276 34620
rect 40132 33992 40184 33998
rect 40132 33934 40184 33940
rect 39948 33312 40000 33318
rect 39948 33254 40000 33260
rect 39856 32428 39908 32434
rect 39856 32370 39908 32376
rect 39960 31346 39988 33254
rect 40316 32904 40368 32910
rect 40316 32846 40368 32852
rect 40224 32428 40276 32434
rect 40224 32370 40276 32376
rect 40236 31482 40264 32370
rect 40224 31476 40276 31482
rect 40224 31418 40276 31424
rect 40328 31346 40356 32846
rect 39948 31340 40000 31346
rect 39948 31282 40000 31288
rect 40316 31340 40368 31346
rect 40316 31282 40368 31288
rect 40040 25288 40092 25294
rect 40040 25230 40092 25236
rect 40052 24818 40080 25230
rect 40224 25220 40276 25226
rect 40224 25162 40276 25168
rect 40236 24886 40264 25162
rect 40224 24880 40276 24886
rect 40224 24822 40276 24828
rect 40040 24812 40092 24818
rect 40040 24754 40092 24760
rect 40040 24608 40092 24614
rect 40040 24550 40092 24556
rect 40052 24274 40080 24550
rect 40420 24274 40448 43302
rect 40590 43200 40646 43302
rect 41878 43200 41934 44000
rect 42522 43200 42578 44000
rect 43166 43200 43222 44000
rect 43810 43200 43866 44000
rect 41326 42936 41382 42945
rect 41326 42871 41382 42880
rect 41144 41064 41196 41070
rect 41144 41006 41196 41012
rect 40500 40452 40552 40458
rect 40500 40394 40552 40400
rect 40512 39642 40540 40394
rect 41156 39642 41184 41006
rect 41340 40186 41368 42871
rect 41892 40594 41920 43200
rect 42536 41206 42564 43200
rect 42524 41200 42576 41206
rect 42524 41142 42576 41148
rect 41880 40588 41932 40594
rect 41880 40530 41932 40536
rect 41328 40180 41380 40186
rect 41328 40122 41380 40128
rect 41972 39976 42024 39982
rect 41972 39918 42024 39924
rect 41420 39840 41472 39846
rect 41420 39782 41472 39788
rect 40500 39636 40552 39642
rect 40500 39578 40552 39584
rect 41144 39636 41196 39642
rect 41144 39578 41196 39584
rect 41432 39438 41460 39782
rect 41984 39642 42012 39918
rect 41972 39636 42024 39642
rect 41972 39578 42024 39584
rect 41878 39536 41934 39545
rect 41878 39471 41934 39480
rect 41236 39432 41288 39438
rect 41236 39374 41288 39380
rect 41420 39432 41472 39438
rect 41420 39374 41472 39380
rect 41248 39098 41276 39374
rect 41236 39092 41288 39098
rect 41236 39034 41288 39040
rect 40684 35080 40736 35086
rect 40684 35022 40736 35028
rect 40696 34542 40724 35022
rect 40684 34536 40736 34542
rect 40684 34478 40736 34484
rect 41248 28082 41276 39034
rect 41328 38412 41380 38418
rect 41328 38354 41380 38360
rect 41340 38185 41368 38354
rect 41326 38176 41382 38185
rect 41326 38111 41382 38120
rect 41328 36236 41380 36242
rect 41328 36178 41380 36184
rect 41340 36145 41368 36178
rect 41326 36136 41382 36145
rect 41326 36071 41382 36080
rect 41328 33448 41380 33454
rect 41326 33416 41328 33425
rect 41380 33416 41382 33425
rect 41326 33351 41382 33360
rect 41326 32056 41382 32065
rect 41326 31991 41382 32000
rect 41340 31890 41368 31991
rect 41328 31884 41380 31890
rect 41328 31826 41380 31832
rect 41432 31346 41460 39374
rect 41892 39030 41920 39471
rect 42248 39364 42300 39370
rect 42248 39306 42300 39312
rect 41880 39024 41932 39030
rect 41880 38966 41932 38972
rect 42156 38344 42208 38350
rect 42156 38286 42208 38292
rect 41696 38276 41748 38282
rect 41696 38218 41748 38224
rect 41708 38010 41736 38218
rect 41696 38004 41748 38010
rect 41696 37946 41748 37952
rect 42168 37466 42196 38286
rect 42156 37460 42208 37466
rect 42156 37402 42208 37408
rect 41604 36780 41656 36786
rect 41604 36722 41656 36728
rect 41616 33998 41644 36722
rect 41972 36576 42024 36582
rect 41972 36518 42024 36524
rect 41984 36242 42012 36518
rect 41972 36236 42024 36242
rect 41972 36178 42024 36184
rect 42156 36168 42208 36174
rect 42156 36110 42208 36116
rect 42168 35698 42196 36110
rect 42156 35692 42208 35698
rect 42156 35634 42208 35640
rect 41972 35080 42024 35086
rect 41972 35022 42024 35028
rect 41878 34776 41934 34785
rect 41878 34711 41934 34720
rect 41892 34678 41920 34711
rect 41880 34672 41932 34678
rect 41880 34614 41932 34620
rect 41604 33992 41656 33998
rect 41604 33934 41656 33940
rect 41512 32836 41564 32842
rect 41512 32778 41564 32784
rect 41524 31482 41552 32778
rect 41512 31476 41564 31482
rect 41512 31418 41564 31424
rect 41420 31340 41472 31346
rect 41472 31300 41552 31328
rect 41420 31282 41472 31288
rect 41326 28656 41382 28665
rect 41326 28591 41328 28600
rect 41380 28591 41382 28600
rect 41328 28562 41380 28568
rect 41420 28484 41472 28490
rect 41420 28426 41472 28432
rect 41432 28218 41460 28426
rect 41420 28212 41472 28218
rect 41420 28154 41472 28160
rect 41236 28076 41288 28082
rect 41236 28018 41288 28024
rect 41524 27470 41552 31300
rect 41512 27464 41564 27470
rect 41512 27406 41564 27412
rect 41328 26920 41380 26926
rect 41328 26862 41380 26868
rect 41340 25945 41368 26862
rect 41326 25936 41382 25945
rect 41326 25871 41382 25880
rect 41512 25288 41564 25294
rect 41234 25256 41290 25265
rect 41512 25230 41564 25236
rect 41234 25191 41290 25200
rect 40500 25152 40552 25158
rect 40500 25094 40552 25100
rect 40040 24268 40092 24274
rect 40040 24210 40092 24216
rect 40408 24268 40460 24274
rect 40408 24210 40460 24216
rect 40512 23186 40540 25094
rect 41248 24750 41276 25191
rect 41236 24744 41288 24750
rect 41236 24686 41288 24692
rect 41326 23896 41382 23905
rect 41326 23831 41382 23840
rect 41340 23662 41368 23831
rect 41328 23656 41380 23662
rect 41328 23598 41380 23604
rect 40500 23180 40552 23186
rect 40500 23122 40552 23128
rect 39948 23112 40000 23118
rect 39948 23054 40000 23060
rect 40316 23112 40368 23118
rect 40316 23054 40368 23060
rect 39960 22642 39988 23054
rect 40328 22778 40356 23054
rect 40316 22772 40368 22778
rect 40316 22714 40368 22720
rect 39948 22636 40000 22642
rect 39948 22578 40000 22584
rect 40684 22432 40736 22438
rect 40684 22374 40736 22380
rect 40696 22098 40724 22374
rect 40684 22092 40736 22098
rect 40684 22034 40736 22040
rect 40960 21480 41012 21486
rect 40960 21422 41012 21428
rect 40972 21146 41000 21422
rect 40960 21140 41012 21146
rect 40960 21082 41012 21088
rect 41524 20942 41552 25230
rect 40316 20936 40368 20942
rect 40316 20878 40368 20884
rect 40868 20936 40920 20942
rect 40868 20878 40920 20884
rect 41512 20936 41564 20942
rect 41512 20878 41564 20884
rect 40328 20602 40356 20878
rect 40316 20596 40368 20602
rect 40316 20538 40368 20544
rect 40224 20256 40276 20262
rect 40224 20198 40276 20204
rect 40236 19446 40264 20198
rect 40880 20058 40908 20878
rect 40868 20052 40920 20058
rect 40868 19994 40920 20000
rect 40316 19848 40368 19854
rect 40316 19790 40368 19796
rect 40224 19440 40276 19446
rect 40224 19382 40276 19388
rect 40040 19372 40092 19378
rect 40040 19314 40092 19320
rect 40052 17882 40080 19314
rect 40328 19242 40356 19790
rect 40408 19712 40460 19718
rect 40408 19654 40460 19660
rect 40316 19236 40368 19242
rect 40316 19178 40368 19184
rect 40420 18834 40448 19654
rect 41236 19304 41288 19310
rect 41236 19246 41288 19252
rect 41248 19145 41276 19246
rect 41234 19136 41290 19145
rect 41234 19071 41290 19080
rect 40408 18828 40460 18834
rect 40408 18770 40460 18776
rect 41326 18456 41382 18465
rect 41326 18391 41382 18400
rect 41340 18222 41368 18391
rect 41328 18216 41380 18222
rect 41328 18158 41380 18164
rect 40040 17876 40092 17882
rect 40040 17818 40092 17824
rect 36636 17672 36688 17678
rect 36636 17614 36688 17620
rect 38476 17672 38528 17678
rect 38476 17614 38528 17620
rect 38752 17672 38804 17678
rect 38752 17614 38804 17620
rect 39764 17672 39816 17678
rect 39764 17614 39816 17620
rect 41144 17672 41196 17678
rect 41144 17614 41196 17620
rect 37924 17536 37976 17542
rect 37924 17478 37976 17484
rect 37936 17202 37964 17478
rect 37924 17196 37976 17202
rect 37924 17138 37976 17144
rect 37648 16992 37700 16998
rect 37648 16934 37700 16940
rect 37660 16590 37688 16934
rect 37648 16584 37700 16590
rect 37648 16526 37700 16532
rect 37280 16448 37332 16454
rect 37280 16390 37332 16396
rect 37292 16114 37320 16390
rect 37280 16108 37332 16114
rect 37280 16050 37332 16056
rect 37464 16040 37516 16046
rect 37464 15982 37516 15988
rect 36084 15904 36136 15910
rect 36084 15846 36136 15852
rect 35900 15496 35952 15502
rect 35900 15438 35952 15444
rect 35808 14816 35860 14822
rect 35808 14758 35860 14764
rect 35716 14408 35768 14414
rect 35716 14350 35768 14356
rect 35728 13938 35756 14350
rect 35820 13938 35848 14758
rect 35912 14618 35940 15438
rect 35900 14612 35952 14618
rect 35900 14554 35952 14560
rect 36096 14414 36124 15846
rect 37476 15706 37504 15982
rect 37464 15700 37516 15706
rect 37464 15642 37516 15648
rect 36544 15496 36596 15502
rect 36544 15438 36596 15444
rect 36268 14612 36320 14618
rect 36268 14554 36320 14560
rect 36084 14408 36136 14414
rect 36084 14350 36136 14356
rect 35992 14068 36044 14074
rect 35992 14010 36044 14016
rect 35716 13932 35768 13938
rect 35716 13874 35768 13880
rect 35808 13932 35860 13938
rect 35808 13874 35860 13880
rect 35728 13462 35756 13874
rect 35716 13456 35768 13462
rect 35716 13398 35768 13404
rect 35716 13320 35768 13326
rect 35716 13262 35768 13268
rect 35728 12850 35756 13262
rect 35716 12844 35768 12850
rect 35716 12786 35768 12792
rect 35544 12406 35664 12434
rect 34796 12300 34848 12306
rect 34796 12242 34848 12248
rect 35164 12096 35216 12102
rect 34992 12044 35164 12050
rect 34992 12038 35216 12044
rect 34992 12022 35204 12038
rect 34992 11830 35020 12022
rect 34980 11824 35032 11830
rect 34980 11766 35032 11772
rect 34612 11756 34664 11762
rect 34612 11698 34664 11704
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 34428 11144 34480 11150
rect 34428 11086 34480 11092
rect 35440 11144 35492 11150
rect 35440 11086 35492 11092
rect 35452 10742 35480 11086
rect 35440 10736 35492 10742
rect 35440 10678 35492 10684
rect 35348 10668 35400 10674
rect 35348 10610 35400 10616
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 35360 10266 35388 10610
rect 35348 10260 35400 10266
rect 35348 10202 35400 10208
rect 35452 10062 35480 10678
rect 35440 10056 35492 10062
rect 35440 9998 35492 10004
rect 34704 9920 34756 9926
rect 34704 9862 34756 9868
rect 34716 9654 34744 9862
rect 34704 9648 34756 9654
rect 34704 9590 34756 9596
rect 34336 9580 34388 9586
rect 34336 9522 34388 9528
rect 33416 9512 33468 9518
rect 33416 9454 33468 9460
rect 32128 9376 32180 9382
rect 32128 9318 32180 9324
rect 31484 9036 31536 9042
rect 31484 8978 31536 8984
rect 32140 8974 32168 9318
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 32128 8968 32180 8974
rect 32128 8910 32180 8916
rect 31300 8832 31352 8838
rect 31300 8774 31352 8780
rect 30840 8560 30892 8566
rect 30840 8502 30892 8508
rect 30288 8424 30340 8430
rect 30288 8366 30340 8372
rect 31312 8362 31340 8774
rect 31300 8356 31352 8362
rect 31300 8298 31352 8304
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 25596 7812 25648 7818
rect 25596 7754 25648 7760
rect 25608 7546 25636 7754
rect 25596 7540 25648 7546
rect 25596 7482 25648 7488
rect 25504 7404 25556 7410
rect 25504 7346 25556 7352
rect 24584 7268 24636 7274
rect 24584 7210 24636 7216
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 20720 6656 20772 6662
rect 20720 6598 20772 6604
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 18604 4208 18656 4214
rect 18604 4150 18656 4156
rect 18144 3936 18196 3942
rect 18144 3878 18196 3884
rect 16856 3732 16908 3738
rect 16684 3692 16856 3720
rect 16684 3602 16712 3692
rect 16856 3674 16908 3680
rect 16672 3596 16724 3602
rect 16672 3538 16724 3544
rect 16856 3596 16908 3602
rect 16856 3538 16908 3544
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 14292 3058 14320 3470
rect 16764 3460 16816 3466
rect 16764 3402 16816 3408
rect 16776 3194 16804 3402
rect 16764 3188 16816 3194
rect 16764 3130 16816 3136
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 15200 2984 15252 2990
rect 15200 2926 15252 2932
rect 15476 2984 15528 2990
rect 15476 2926 15528 2932
rect 15212 2650 15240 2926
rect 15200 2644 15252 2650
rect 15200 2586 15252 2592
rect 13728 2508 13780 2514
rect 13728 2450 13780 2456
rect 11624 1686 11744 1714
rect 11624 800 11652 1686
rect 15488 800 15516 2926
rect 16868 2774 16896 3538
rect 16948 3392 17000 3398
rect 16948 3334 17000 3340
rect 16960 3194 16988 3334
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 18156 3058 18184 3878
rect 18616 3534 18644 4150
rect 22468 4072 22520 4078
rect 22468 4014 22520 4020
rect 22836 4072 22888 4078
rect 22836 4014 22888 4020
rect 23204 4072 23256 4078
rect 23204 4014 23256 4020
rect 19524 3936 19576 3942
rect 19524 3878 19576 3884
rect 21824 3936 21876 3942
rect 21824 3878 21876 3884
rect 19536 3602 19564 3878
rect 19524 3596 19576 3602
rect 19524 3538 19576 3544
rect 19984 3596 20036 3602
rect 19984 3538 20036 3544
rect 18604 3528 18656 3534
rect 18604 3470 18656 3476
rect 18328 3392 18380 3398
rect 18328 3334 18380 3340
rect 18340 3126 18368 3334
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 18328 3120 18380 3126
rect 18328 3062 18380 3068
rect 18144 3052 18196 3058
rect 18144 2994 18196 3000
rect 18696 2984 18748 2990
rect 18696 2926 18748 2932
rect 16776 2746 16896 2774
rect 16776 800 16804 2746
rect 18708 800 18736 2926
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 19996 800 20024 3538
rect 20536 3460 20588 3466
rect 20536 3402 20588 3408
rect 20548 3194 20576 3402
rect 20536 3188 20588 3194
rect 20536 3130 20588 3136
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 20640 2446 20668 2994
rect 21836 2514 21864 3878
rect 22480 3738 22508 4014
rect 22468 3732 22520 3738
rect 22468 3674 22520 3680
rect 22848 3194 22876 4014
rect 22836 3188 22888 3194
rect 22836 3130 22888 3136
rect 22008 2848 22060 2854
rect 22008 2790 22060 2796
rect 22020 2514 22048 2790
rect 21824 2508 21876 2514
rect 21824 2450 21876 2456
rect 22008 2508 22060 2514
rect 22008 2450 22060 2456
rect 22560 2508 22612 2514
rect 22560 2450 22612 2456
rect 20628 2440 20680 2446
rect 20628 2382 20680 2388
rect 22572 800 22600 2450
rect 23216 800 23244 4014
rect 34704 3936 34756 3942
rect 34704 3878 34756 3884
rect 34716 3602 34744 3878
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 34704 3596 34756 3602
rect 34888 3596 34940 3602
rect 34704 3538 34756 3544
rect 34808 3556 34888 3584
rect 23480 3528 23532 3534
rect 23480 3470 23532 3476
rect 27620 3528 27672 3534
rect 27620 3470 27672 3476
rect 27804 3528 27856 3534
rect 27804 3470 27856 3476
rect 23492 3058 23520 3470
rect 23664 3392 23716 3398
rect 23664 3334 23716 3340
rect 23676 3126 23704 3334
rect 23664 3120 23716 3126
rect 23664 3062 23716 3068
rect 23480 3052 23532 3058
rect 23480 2994 23532 3000
rect 23848 2984 23900 2990
rect 23848 2926 23900 2932
rect 23860 800 23888 2926
rect 27632 2446 27660 3470
rect 27816 3058 27844 3470
rect 27804 3052 27856 3058
rect 27804 2994 27856 3000
rect 27988 2984 28040 2990
rect 27988 2926 28040 2932
rect 28356 2984 28408 2990
rect 28356 2926 28408 2932
rect 28000 2650 28028 2926
rect 27988 2644 28040 2650
rect 27988 2586 28040 2592
rect 27620 2440 27672 2446
rect 27620 2382 27672 2388
rect 28368 800 28396 2926
rect 34808 800 34836 3556
rect 34888 3538 34940 3544
rect 35544 3466 35572 12406
rect 35624 12164 35676 12170
rect 35624 12106 35676 12112
rect 35636 11626 35664 12106
rect 35624 11620 35676 11626
rect 35624 11562 35676 11568
rect 35728 11150 35756 12786
rect 35820 12170 35848 13874
rect 36004 12986 36032 14010
rect 35992 12980 36044 12986
rect 35992 12922 36044 12928
rect 36096 12238 36124 14350
rect 36176 13864 36228 13870
rect 36176 13806 36228 13812
rect 36188 13326 36216 13806
rect 36176 13320 36228 13326
rect 36176 13262 36228 13268
rect 36188 13190 36216 13262
rect 36280 13258 36308 14554
rect 36556 13530 36584 15438
rect 38488 14890 38516 17614
rect 38764 17270 38792 17614
rect 39776 17338 39804 17614
rect 39764 17332 39816 17338
rect 39764 17274 39816 17280
rect 38752 17264 38804 17270
rect 38752 17206 38804 17212
rect 40960 16108 41012 16114
rect 40960 16050 41012 16056
rect 38936 16040 38988 16046
rect 38936 15982 38988 15988
rect 38476 14884 38528 14890
rect 38476 14826 38528 14832
rect 37188 14408 37240 14414
rect 37188 14350 37240 14356
rect 36636 14272 36688 14278
rect 36636 14214 36688 14220
rect 36544 13524 36596 13530
rect 36544 13466 36596 13472
rect 36268 13252 36320 13258
rect 36268 13194 36320 13200
rect 36176 13184 36228 13190
rect 36176 13126 36228 13132
rect 36084 12232 36136 12238
rect 36084 12174 36136 12180
rect 35808 12164 35860 12170
rect 35808 12106 35860 12112
rect 35992 12096 36044 12102
rect 35992 12038 36044 12044
rect 36004 11694 36032 12038
rect 36096 11830 36124 12174
rect 36188 11898 36216 13126
rect 36280 12850 36308 13194
rect 36648 12850 36676 14214
rect 36820 13796 36872 13802
rect 36820 13738 36872 13744
rect 36832 13530 36860 13738
rect 36820 13524 36872 13530
rect 36820 13466 36872 13472
rect 37200 12850 37228 14350
rect 37372 13932 37424 13938
rect 37372 13874 37424 13880
rect 37384 13326 37412 13874
rect 37372 13320 37424 13326
rect 37372 13262 37424 13268
rect 37464 13184 37516 13190
rect 37464 13126 37516 13132
rect 37476 12918 37504 13126
rect 37464 12912 37516 12918
rect 37464 12854 37516 12860
rect 36268 12844 36320 12850
rect 36268 12786 36320 12792
rect 36636 12844 36688 12850
rect 36636 12786 36688 12792
rect 37188 12844 37240 12850
rect 37188 12786 37240 12792
rect 36280 12170 36308 12786
rect 36360 12708 36412 12714
rect 36360 12650 36412 12656
rect 36372 12434 36400 12650
rect 36372 12406 36492 12434
rect 36268 12164 36320 12170
rect 36268 12106 36320 12112
rect 36176 11892 36228 11898
rect 36176 11834 36228 11840
rect 36084 11824 36136 11830
rect 36084 11766 36136 11772
rect 36280 11762 36308 12106
rect 36360 12096 36412 12102
rect 36360 12038 36412 12044
rect 36268 11756 36320 11762
rect 36268 11698 36320 11704
rect 35992 11688 36044 11694
rect 35992 11630 36044 11636
rect 36268 11620 36320 11626
rect 36268 11562 36320 11568
rect 35992 11552 36044 11558
rect 35992 11494 36044 11500
rect 35900 11280 35952 11286
rect 35900 11222 35952 11228
rect 35716 11144 35768 11150
rect 35716 11086 35768 11092
rect 35624 11008 35676 11014
rect 35624 10950 35676 10956
rect 35636 10810 35664 10950
rect 35624 10804 35676 10810
rect 35624 10746 35676 10752
rect 35912 10674 35940 11222
rect 36004 11150 36032 11494
rect 36176 11212 36228 11218
rect 36176 11154 36228 11160
rect 35992 11144 36044 11150
rect 35992 11086 36044 11092
rect 35900 10668 35952 10674
rect 35900 10610 35952 10616
rect 35716 10464 35768 10470
rect 35716 10406 35768 10412
rect 35728 10062 35756 10406
rect 36188 10198 36216 11154
rect 36280 10606 36308 11562
rect 36372 11286 36400 12038
rect 36464 11286 36492 12406
rect 37004 12232 37056 12238
rect 37004 12174 37056 12180
rect 37016 11898 37044 12174
rect 37004 11892 37056 11898
rect 37004 11834 37056 11840
rect 37004 11756 37056 11762
rect 37004 11698 37056 11704
rect 36820 11688 36872 11694
rect 36820 11630 36872 11636
rect 36360 11280 36412 11286
rect 36360 11222 36412 11228
rect 36452 11280 36504 11286
rect 36452 11222 36504 11228
rect 36464 11150 36492 11222
rect 36832 11150 36860 11630
rect 37016 11150 37044 11698
rect 36452 11144 36504 11150
rect 36452 11086 36504 11092
rect 36820 11144 36872 11150
rect 36820 11086 36872 11092
rect 37004 11144 37056 11150
rect 37004 11086 37056 11092
rect 36268 10600 36320 10606
rect 36268 10542 36320 10548
rect 36176 10192 36228 10198
rect 36176 10134 36228 10140
rect 36832 10130 36860 11086
rect 37200 10674 37228 12786
rect 37556 11008 37608 11014
rect 37556 10950 37608 10956
rect 37188 10668 37240 10674
rect 37188 10610 37240 10616
rect 36820 10124 36872 10130
rect 36820 10066 36872 10072
rect 37568 10062 37596 10950
rect 35716 10056 35768 10062
rect 35716 9998 35768 10004
rect 37556 10056 37608 10062
rect 37556 9998 37608 10004
rect 38476 5704 38528 5710
rect 38476 5646 38528 5652
rect 38488 5234 38516 5646
rect 38660 5568 38712 5574
rect 38660 5510 38712 5516
rect 38672 5302 38700 5510
rect 38660 5296 38712 5302
rect 38660 5238 38712 5244
rect 38476 5228 38528 5234
rect 38476 5170 38528 5176
rect 36728 4616 36780 4622
rect 36728 4558 36780 4564
rect 37556 4616 37608 4622
rect 37556 4558 37608 4564
rect 35624 3936 35676 3942
rect 35624 3878 35676 3884
rect 35532 3460 35584 3466
rect 35532 3402 35584 3408
rect 35636 3126 35664 3878
rect 36740 3602 36768 4558
rect 37464 3936 37516 3942
rect 37464 3878 37516 3884
rect 36728 3596 36780 3602
rect 36728 3538 36780 3544
rect 37372 3596 37424 3602
rect 37372 3538 37424 3544
rect 37188 3460 37240 3466
rect 37188 3402 37240 3408
rect 36360 3392 36412 3398
rect 36360 3334 36412 3340
rect 35624 3120 35676 3126
rect 35624 3062 35676 3068
rect 35808 2984 35860 2990
rect 35808 2926 35860 2932
rect 36084 2984 36136 2990
rect 36084 2926 36136 2932
rect 35440 2916 35492 2922
rect 35440 2858 35492 2864
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 35452 800 35480 2858
rect 35820 2650 35848 2926
rect 35808 2644 35860 2650
rect 35808 2586 35860 2592
rect 35900 2440 35952 2446
rect 35900 2382 35952 2388
rect 35912 2106 35940 2382
rect 35900 2100 35952 2106
rect 35900 2042 35952 2048
rect 36096 800 36124 2926
rect 36372 2446 36400 3334
rect 37200 2650 37228 3402
rect 37188 2644 37240 2650
rect 37188 2586 37240 2592
rect 36360 2440 36412 2446
rect 36360 2382 36412 2388
rect 37384 800 37412 3538
rect 37476 2514 37504 3878
rect 37568 3058 37596 4558
rect 37832 4140 37884 4146
rect 37832 4082 37884 4088
rect 37648 3936 37700 3942
rect 37648 3878 37700 3884
rect 37556 3052 37608 3058
rect 37556 2994 37608 3000
rect 37660 2514 37688 3878
rect 37464 2508 37516 2514
rect 37464 2450 37516 2456
rect 37648 2508 37700 2514
rect 37648 2450 37700 2456
rect 37844 2378 37872 4082
rect 38660 3936 38712 3942
rect 38660 3878 38712 3884
rect 38672 3126 38700 3878
rect 38660 3120 38712 3126
rect 38660 3062 38712 3068
rect 38948 2922 38976 15982
rect 40316 15904 40368 15910
rect 40316 15846 40368 15852
rect 40500 15904 40552 15910
rect 40500 15846 40552 15852
rect 40328 15570 40356 15846
rect 40512 15570 40540 15846
rect 40316 15564 40368 15570
rect 40316 15506 40368 15512
rect 40500 15564 40552 15570
rect 40500 15506 40552 15512
rect 40776 12640 40828 12646
rect 40776 12582 40828 12588
rect 40788 12306 40816 12582
rect 40972 12434 41000 16050
rect 40972 12406 41092 12434
rect 40776 12300 40828 12306
rect 40776 12242 40828 12248
rect 40316 11552 40368 11558
rect 40316 11494 40368 11500
rect 40328 11218 40356 11494
rect 40316 11212 40368 11218
rect 40316 11154 40368 11160
rect 40316 10464 40368 10470
rect 40316 10406 40368 10412
rect 40328 10130 40356 10406
rect 40316 10124 40368 10130
rect 40316 10066 40368 10072
rect 40500 7744 40552 7750
rect 40500 7686 40552 7692
rect 40512 6730 40540 7686
rect 40960 7200 41012 7206
rect 40960 7142 41012 7148
rect 40972 6866 41000 7142
rect 40960 6860 41012 6866
rect 40960 6802 41012 6808
rect 40500 6724 40552 6730
rect 40500 6666 40552 6672
rect 40316 6112 40368 6118
rect 40316 6054 40368 6060
rect 39856 5704 39908 5710
rect 39856 5646 39908 5652
rect 39028 4616 39080 4622
rect 39028 4558 39080 4564
rect 39120 4616 39172 4622
rect 39120 4558 39172 4564
rect 39040 4146 39068 4558
rect 39028 4140 39080 4146
rect 39028 4082 39080 4088
rect 39132 4078 39160 4558
rect 39764 4480 39816 4486
rect 39764 4422 39816 4428
rect 39776 4214 39804 4422
rect 39764 4208 39816 4214
rect 39764 4150 39816 4156
rect 39120 4072 39172 4078
rect 39120 4014 39172 4020
rect 39764 3460 39816 3466
rect 39764 3402 39816 3408
rect 39304 2984 39356 2990
rect 39304 2926 39356 2932
rect 38936 2916 38988 2922
rect 38936 2858 38988 2864
rect 37832 2372 37884 2378
rect 37832 2314 37884 2320
rect 39316 800 39344 2926
rect 6564 734 6776 762
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 23846 0 23902 800
rect 25134 0 25190 800
rect 25778 0 25834 800
rect 26422 0 26478 800
rect 27066 0 27122 800
rect 28354 0 28410 800
rect 28998 0 29054 800
rect 29642 0 29698 800
rect 30930 0 30986 800
rect 31574 0 31630 800
rect 32218 0 32274 800
rect 32862 0 32918 800
rect 34150 0 34206 800
rect 34794 0 34850 800
rect 35438 0 35494 800
rect 36082 0 36138 800
rect 37370 0 37426 800
rect 38014 0 38070 800
rect 38658 0 38714 800
rect 39302 0 39358 800
rect 39776 785 39804 3402
rect 39868 3058 39896 5646
rect 40040 5024 40092 5030
rect 40040 4966 40092 4972
rect 40052 3126 40080 4966
rect 40328 4690 40356 6054
rect 41064 5234 41092 12406
rect 41156 9586 41184 17614
rect 41420 16516 41472 16522
rect 41420 16458 41472 16464
rect 41432 16250 41460 16458
rect 41420 16244 41472 16250
rect 41420 16186 41472 16192
rect 41524 15638 41552 20878
rect 41512 15632 41564 15638
rect 41512 15574 41564 15580
rect 41326 15056 41382 15065
rect 41326 14991 41382 15000
rect 41340 14958 41368 14991
rect 41328 14952 41380 14958
rect 41328 14894 41380 14900
rect 41420 14952 41472 14958
rect 41420 14894 41472 14900
rect 41432 14618 41460 14894
rect 41420 14612 41472 14618
rect 41420 14554 41472 14560
rect 41236 14408 41288 14414
rect 41236 14350 41288 14356
rect 41144 9580 41196 9586
rect 41144 9522 41196 9528
rect 41248 5710 41276 14350
rect 41328 13388 41380 13394
rect 41328 13330 41380 13336
rect 41340 13025 41368 13330
rect 41512 13252 41564 13258
rect 41512 13194 41564 13200
rect 41326 13016 41382 13025
rect 41524 12986 41552 13194
rect 41326 12951 41382 12960
rect 41512 12980 41564 12986
rect 41512 12922 41564 12928
rect 41418 12880 41474 12889
rect 41418 12815 41420 12824
rect 41472 12815 41474 12824
rect 41420 12786 41472 12792
rect 41432 11762 41460 12786
rect 41512 12164 41564 12170
rect 41512 12106 41564 12112
rect 41524 11898 41552 12106
rect 41512 11892 41564 11898
rect 41512 11834 41564 11840
rect 41420 11756 41472 11762
rect 41420 11698 41472 11704
rect 41420 11076 41472 11082
rect 41420 11018 41472 11024
rect 41432 10810 41460 11018
rect 41420 10804 41472 10810
rect 41420 10746 41472 10752
rect 41420 9988 41472 9994
rect 41420 9930 41472 9936
rect 41432 9654 41460 9930
rect 41420 9648 41472 9654
rect 41420 9590 41472 9596
rect 41616 7886 41644 33934
rect 41696 33856 41748 33862
rect 41696 33798 41748 33804
rect 41708 33590 41736 33798
rect 41696 33584 41748 33590
rect 41696 33526 41748 33532
rect 41984 33522 42012 35022
rect 41972 33516 42024 33522
rect 41972 33458 42024 33464
rect 42156 32836 42208 32842
rect 42156 32778 42208 32784
rect 42168 32745 42196 32778
rect 42154 32736 42210 32745
rect 42154 32671 42210 32680
rect 42156 31816 42208 31822
rect 42156 31758 42208 31764
rect 41972 31748 42024 31754
rect 41972 31690 42024 31696
rect 41984 30938 42012 31690
rect 41972 30932 42024 30938
rect 41972 30874 42024 30880
rect 41880 30728 41932 30734
rect 41880 30670 41932 30676
rect 41788 28960 41840 28966
rect 41788 28902 41840 28908
rect 41800 28626 41828 28902
rect 41788 28620 41840 28626
rect 41788 28562 41840 28568
rect 41696 27328 41748 27334
rect 41696 27270 41748 27276
rect 41708 27062 41736 27270
rect 41696 27056 41748 27062
rect 41696 26998 41748 27004
rect 41892 27010 41920 30670
rect 42168 30258 42196 31758
rect 42156 30252 42208 30258
rect 42156 30194 42208 30200
rect 42064 29572 42116 29578
rect 42064 29514 42116 29520
rect 41972 29504 42024 29510
rect 41972 29446 42024 29452
rect 41984 27130 42012 29446
rect 42076 29345 42104 29514
rect 42062 29336 42118 29345
rect 42062 29271 42118 29280
rect 41972 27124 42024 27130
rect 41972 27066 42024 27072
rect 41892 26982 42012 27010
rect 41880 26920 41932 26926
rect 41880 26862 41932 26868
rect 41892 26586 41920 26862
rect 41880 26580 41932 26586
rect 41880 26522 41932 26528
rect 41880 25696 41932 25702
rect 41880 25638 41932 25644
rect 41788 25288 41840 25294
rect 41788 25230 41840 25236
rect 41696 23656 41748 23662
rect 41696 23598 41748 23604
rect 41708 21146 41736 23598
rect 41696 21140 41748 21146
rect 41696 21082 41748 21088
rect 41696 20256 41748 20262
rect 41696 20198 41748 20204
rect 41708 19922 41736 20198
rect 41696 19916 41748 19922
rect 41696 19858 41748 19864
rect 41696 18216 41748 18222
rect 41696 18158 41748 18164
rect 41708 17882 41736 18158
rect 41696 17876 41748 17882
rect 41696 17818 41748 17824
rect 41696 16652 41748 16658
rect 41696 16594 41748 16600
rect 41708 16425 41736 16594
rect 41694 16416 41750 16425
rect 41694 16351 41750 16360
rect 41800 13818 41828 25230
rect 41892 23730 41920 25638
rect 41880 23724 41932 23730
rect 41880 23666 41932 23672
rect 41878 23216 41934 23225
rect 41878 23151 41934 23160
rect 41892 21622 41920 23151
rect 41984 22642 42012 26982
rect 41972 22636 42024 22642
rect 41972 22578 42024 22584
rect 42154 22536 42210 22545
rect 42154 22471 42210 22480
rect 42168 22098 42196 22471
rect 42156 22092 42208 22098
rect 42156 22034 42208 22040
rect 41880 21616 41932 21622
rect 41880 21558 41932 21564
rect 42154 19816 42210 19825
rect 42154 19751 42156 19760
rect 42208 19751 42210 19760
rect 42156 19722 42208 19728
rect 42064 18692 42116 18698
rect 42064 18634 42116 18640
rect 41880 18216 41932 18222
rect 41880 18158 41932 18164
rect 41892 17882 41920 18158
rect 41880 17876 41932 17882
rect 41880 17818 41932 17824
rect 41880 16040 41932 16046
rect 41880 15982 41932 15988
rect 41892 14498 41920 15982
rect 41972 14952 42024 14958
rect 41972 14894 42024 14900
rect 41984 14618 42012 14894
rect 41972 14612 42024 14618
rect 41972 14554 42024 14560
rect 41892 14470 42012 14498
rect 41708 13790 41828 13818
rect 41708 12850 41736 13790
rect 41788 13728 41840 13734
rect 41788 13670 41840 13676
rect 41800 13394 41828 13670
rect 41788 13388 41840 13394
rect 41788 13330 41840 13336
rect 41696 12844 41748 12850
rect 41696 12786 41748 12792
rect 41604 7880 41656 7886
rect 41604 7822 41656 7828
rect 41880 7404 41932 7410
rect 41880 7346 41932 7352
rect 41892 6905 41920 7346
rect 41878 6896 41934 6905
rect 41878 6831 41934 6840
rect 41788 6112 41840 6118
rect 41788 6054 41840 6060
rect 41696 5772 41748 5778
rect 41696 5714 41748 5720
rect 41236 5704 41288 5710
rect 41236 5646 41288 5652
rect 41052 5228 41104 5234
rect 41052 5170 41104 5176
rect 41420 5228 41472 5234
rect 41420 5170 41472 5176
rect 40316 4684 40368 4690
rect 40316 4626 40368 4632
rect 41326 4176 41382 4185
rect 41326 4111 41382 4120
rect 41340 4078 41368 4111
rect 41328 4072 41380 4078
rect 41328 4014 41380 4020
rect 41236 3392 41288 3398
rect 41236 3334 41288 3340
rect 40040 3120 40092 3126
rect 40040 3062 40092 3068
rect 39856 3052 39908 3058
rect 39856 2994 39908 3000
rect 40592 2984 40644 2990
rect 40592 2926 40644 2932
rect 39948 2372 40000 2378
rect 39948 2314 40000 2320
rect 39960 2145 39988 2314
rect 39946 2136 40002 2145
rect 39946 2071 40002 2080
rect 40604 800 40632 2926
rect 41248 800 41276 3334
rect 41432 2582 41460 5170
rect 41512 5024 41564 5030
rect 41512 4966 41564 4972
rect 41524 4690 41552 4966
rect 41512 4684 41564 4690
rect 41512 4626 41564 4632
rect 41420 2576 41472 2582
rect 41420 2518 41472 2524
rect 41328 2508 41380 2514
rect 41328 2450 41380 2456
rect 39762 776 39818 785
rect 39762 711 39818 720
rect 40590 0 40646 800
rect 41234 0 41290 800
rect 41340 105 41368 2450
rect 41708 2378 41736 5714
rect 41800 3602 41828 6054
rect 41984 5710 42012 14470
rect 41972 5704 42024 5710
rect 41972 5646 42024 5652
rect 42076 5658 42104 18634
rect 42156 16992 42208 16998
rect 42156 16934 42208 16940
rect 42168 16658 42196 16934
rect 42156 16652 42208 16658
rect 42156 16594 42208 16600
rect 42154 15736 42210 15745
rect 42154 15671 42210 15680
rect 42168 15570 42196 15671
rect 42156 15564 42208 15570
rect 42156 15506 42208 15512
rect 42154 12336 42210 12345
rect 42154 12271 42156 12280
rect 42208 12271 42210 12280
rect 42156 12242 42208 12248
rect 42156 11076 42208 11082
rect 42156 11018 42208 11024
rect 42168 10985 42196 11018
rect 42154 10976 42210 10985
rect 42154 10911 42210 10920
rect 42260 10674 42288 39306
rect 42340 37868 42392 37874
rect 42340 37810 42392 37816
rect 42352 16114 42380 37810
rect 42340 16108 42392 16114
rect 42340 16050 42392 16056
rect 42248 10668 42300 10674
rect 42248 10610 42300 10616
rect 42154 10296 42210 10305
rect 42154 10231 42210 10240
rect 42168 10130 42196 10231
rect 42156 10124 42208 10130
rect 42156 10066 42208 10072
rect 42156 6724 42208 6730
rect 42156 6666 42208 6672
rect 42168 6225 42196 6666
rect 42154 6216 42210 6225
rect 42154 6151 42210 6160
rect 42076 5630 42196 5658
rect 41972 5568 42024 5574
rect 41972 5510 42024 5516
rect 42064 5568 42116 5574
rect 42064 5510 42116 5516
rect 41880 4684 41932 4690
rect 41880 4626 41932 4632
rect 41788 3596 41840 3602
rect 41788 3538 41840 3544
rect 41696 2372 41748 2378
rect 41696 2314 41748 2320
rect 41892 800 41920 4626
rect 41984 3466 42012 5510
rect 41972 3460 42024 3466
rect 41972 3402 42024 3408
rect 42076 2514 42104 5510
rect 42168 3398 42196 5630
rect 43168 5160 43220 5166
rect 43168 5102 43220 5108
rect 42156 3392 42208 3398
rect 42156 3334 42208 3340
rect 42064 2508 42116 2514
rect 42064 2450 42116 2456
rect 43180 800 43208 5102
rect 41326 96 41382 105
rect 41326 31 41382 40
rect 41878 0 41934 800
rect 43166 0 43222 800
rect 43810 0 43866 800
<< via2 >>
rect 1858 40840 1914 40896
rect 2870 42880 2926 42936
rect 2962 41520 3018 41576
rect 1858 21800 1914 21856
rect 1858 19760 1914 19816
rect 1858 16360 1914 16416
rect 1398 8916 1400 8936
rect 1400 8916 1452 8936
rect 1452 8916 1454 8936
rect 1398 8880 1454 8916
rect 1858 5480 1914 5536
rect 1398 3476 1400 3496
rect 1400 3476 1452 3496
rect 1452 3476 1454 3496
rect 1398 3440 1454 3476
rect 2778 38120 2834 38176
rect 3514 40160 3570 40216
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 3606 36760 3662 36816
rect 2870 36080 2926 36136
rect 2778 28620 2834 28656
rect 2778 28600 2780 28620
rect 2780 28600 2832 28620
rect 2832 28600 2834 28620
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 2778 21120 2834 21176
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 2778 17720 2834 17776
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 2778 15000 2834 15056
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 2870 13640 2926 13696
rect 2778 12300 2834 12336
rect 2778 12280 2780 12300
rect 2780 12280 2832 12300
rect 2832 12280 2834 12300
rect 2778 10240 2834 10296
rect 2778 8200 2834 8256
rect 2778 4800 2834 4856
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4066 6860 4122 6896
rect 4066 6840 4068 6860
rect 4068 6840 4120 6860
rect 4120 6840 4122 6860
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 3146 4140 3202 4176
rect 3146 4120 3148 4140
rect 3148 4120 3200 4140
rect 3200 4120 3202 4140
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 2778 1400 2834 1456
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 3422 2080 3478 2136
rect 5630 24268 5686 24304
rect 5630 24248 5632 24268
rect 5632 24248 5684 24268
rect 5684 24248 5686 24268
rect 8206 39480 8262 39536
rect 9586 38956 9642 38992
rect 9586 38936 9588 38956
rect 9588 38936 9640 38956
rect 9640 38936 9642 38956
rect 12346 38836 12348 38856
rect 12348 38836 12400 38856
rect 12400 38836 12402 38856
rect 12346 38800 12402 38836
rect 11702 12824 11758 12880
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 14462 36372 14518 36408
rect 14462 36352 14464 36372
rect 14464 36352 14516 36372
rect 14516 36352 14518 36372
rect 18234 36352 18290 36408
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 13266 17620 13268 17640
rect 13268 17620 13320 17640
rect 13320 17620 13322 17640
rect 13266 17584 13322 17620
rect 14830 20848 14886 20904
rect 15290 17604 15346 17640
rect 15290 17584 15292 17604
rect 15292 17584 15344 17604
rect 15344 17584 15346 17604
rect 16578 20884 16580 20904
rect 16580 20884 16632 20904
rect 16632 20884 16634 20904
rect 16578 20848 16634 20884
rect 14278 15580 14280 15600
rect 14280 15580 14332 15600
rect 14332 15580 14334 15600
rect 14278 15544 14334 15580
rect 15842 17584 15898 17640
rect 16118 15564 16174 15600
rect 16118 15544 16120 15564
rect 16120 15544 16172 15564
rect 16172 15544 16174 15564
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 17590 20868 17646 20904
rect 17590 20848 17592 20868
rect 17592 20848 17644 20868
rect 17644 20848 17646 20868
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 32862 39480 32918 39536
rect 29274 38936 29330 38992
rect 39302 41520 39358 41576
rect 39302 40160 39358 40216
rect 26606 38800 26662 38856
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 29182 28600 29238 28656
rect 29090 28328 29146 28384
rect 27802 22092 27858 22128
rect 27802 22072 27804 22092
rect 27804 22072 27856 22092
rect 27856 22072 27858 22092
rect 28906 22108 28954 22128
rect 28954 22108 28962 22128
rect 28906 22072 28962 22108
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 39394 35400 39450 35456
rect 37554 24284 37556 24304
rect 37556 24284 37608 24304
rect 37608 24284 37610 24304
rect 37554 24248 37610 24284
rect 39578 20440 39634 20496
rect 41326 42880 41382 42936
rect 41878 39480 41934 39536
rect 41326 38120 41382 38176
rect 41326 36080 41382 36136
rect 41326 33396 41328 33416
rect 41328 33396 41380 33416
rect 41380 33396 41382 33416
rect 41326 33360 41382 33396
rect 41326 32000 41382 32056
rect 41878 34720 41934 34776
rect 41326 28620 41382 28656
rect 41326 28600 41328 28620
rect 41328 28600 41380 28620
rect 41380 28600 41382 28620
rect 41326 25880 41382 25936
rect 41234 25200 41290 25256
rect 41326 23840 41382 23896
rect 41234 19080 41290 19136
rect 41326 18400 41382 18456
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 41326 15000 41382 15056
rect 41326 12960 41382 13016
rect 41418 12844 41474 12880
rect 41418 12824 41420 12844
rect 41420 12824 41472 12844
rect 41472 12824 41474 12844
rect 42154 32680 42210 32736
rect 42062 29280 42118 29336
rect 41694 16360 41750 16416
rect 41878 23160 41934 23216
rect 42154 22480 42210 22536
rect 42154 19780 42210 19816
rect 42154 19760 42156 19780
rect 42156 19760 42208 19780
rect 42208 19760 42210 19780
rect 41878 6840 41934 6896
rect 41326 4120 41382 4176
rect 39946 2080 40002 2136
rect 39762 720 39818 776
rect 42154 15680 42210 15736
rect 42154 12300 42210 12336
rect 42154 12280 42156 12300
rect 42156 12280 42208 12300
rect 42208 12280 42210 12300
rect 42154 10920 42210 10976
rect 42154 10240 42210 10296
rect 42154 6160 42210 6216
rect 41326 40 41382 96
<< metal3 >>
rect 0 43528 800 43648
rect 0 42938 800 42968
rect 2865 42938 2931 42941
rect 0 42936 2931 42938
rect 0 42880 2870 42936
rect 2926 42880 2931 42936
rect 0 42878 2931 42880
rect 0 42848 800 42878
rect 2865 42875 2931 42878
rect 41321 42938 41387 42941
rect 43200 42938 44000 42968
rect 41321 42936 44000 42938
rect 41321 42880 41326 42936
rect 41382 42880 44000 42936
rect 41321 42878 44000 42880
rect 41321 42875 41387 42878
rect 43200 42848 44000 42878
rect 43200 42168 44000 42288
rect 0 41578 800 41608
rect 2957 41578 3023 41581
rect 0 41576 3023 41578
rect 0 41520 2962 41576
rect 3018 41520 3023 41576
rect 0 41518 3023 41520
rect 0 41488 800 41518
rect 2957 41515 3023 41518
rect 39297 41578 39363 41581
rect 43200 41578 44000 41608
rect 39297 41576 44000 41578
rect 39297 41520 39302 41576
rect 39358 41520 44000 41576
rect 39297 41518 44000 41520
rect 39297 41515 39363 41518
rect 43200 41488 44000 41518
rect 19568 41376 19888 41377
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 41311 19888 41312
rect 0 40898 800 40928
rect 1853 40898 1919 40901
rect 0 40896 1919 40898
rect 0 40840 1858 40896
rect 1914 40840 1919 40896
rect 0 40838 1919 40840
rect 0 40808 800 40838
rect 1853 40835 1919 40838
rect 4208 40832 4528 40833
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 40767 4528 40768
rect 34928 40832 35248 40833
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 40767 35248 40768
rect 19568 40288 19888 40289
rect 0 40218 800 40248
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 40223 19888 40224
rect 3509 40218 3575 40221
rect 0 40216 3575 40218
rect 0 40160 3514 40216
rect 3570 40160 3575 40216
rect 0 40158 3575 40160
rect 0 40128 800 40158
rect 3509 40155 3575 40158
rect 39297 40218 39363 40221
rect 43200 40218 44000 40248
rect 39297 40216 44000 40218
rect 39297 40160 39302 40216
rect 39358 40160 44000 40216
rect 39297 40158 44000 40160
rect 39297 40155 39363 40158
rect 43200 40128 44000 40158
rect 4208 39744 4528 39745
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 39679 4528 39680
rect 34928 39744 35248 39745
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 39679 35248 39680
rect 0 39448 800 39568
rect 8201 39538 8267 39541
rect 32857 39538 32923 39541
rect 8201 39536 32923 39538
rect 8201 39480 8206 39536
rect 8262 39480 32862 39536
rect 32918 39480 32923 39536
rect 8201 39478 32923 39480
rect 8201 39475 8267 39478
rect 32857 39475 32923 39478
rect 41873 39538 41939 39541
rect 43200 39538 44000 39568
rect 41873 39536 44000 39538
rect 41873 39480 41878 39536
rect 41934 39480 44000 39536
rect 41873 39478 44000 39480
rect 41873 39475 41939 39478
rect 43200 39448 44000 39478
rect 19568 39200 19888 39201
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 39135 19888 39136
rect 9581 38994 9647 38997
rect 29269 38994 29335 38997
rect 9581 38992 29335 38994
rect 9581 38936 9586 38992
rect 9642 38936 29274 38992
rect 29330 38936 29335 38992
rect 9581 38934 29335 38936
rect 9581 38931 9647 38934
rect 29269 38931 29335 38934
rect 12341 38858 12407 38861
rect 26601 38858 26667 38861
rect 12341 38856 26667 38858
rect 12341 38800 12346 38856
rect 12402 38800 26606 38856
rect 26662 38800 26667 38856
rect 12341 38798 26667 38800
rect 12341 38795 12407 38798
rect 26601 38795 26667 38798
rect 43200 38768 44000 38888
rect 4208 38656 4528 38657
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 38591 4528 38592
rect 34928 38656 35248 38657
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 38591 35248 38592
rect 0 38178 800 38208
rect 2773 38178 2839 38181
rect 0 38176 2839 38178
rect 0 38120 2778 38176
rect 2834 38120 2839 38176
rect 0 38118 2839 38120
rect 0 38088 800 38118
rect 2773 38115 2839 38118
rect 41321 38178 41387 38181
rect 43200 38178 44000 38208
rect 41321 38176 44000 38178
rect 41321 38120 41326 38176
rect 41382 38120 44000 38176
rect 41321 38118 44000 38120
rect 41321 38115 41387 38118
rect 19568 38112 19888 38113
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 43200 38088 44000 38118
rect 19568 38047 19888 38048
rect 4208 37568 4528 37569
rect 0 37408 800 37528
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 0 36818 800 36848
rect 3601 36818 3667 36821
rect 0 36816 3667 36818
rect 0 36760 3606 36816
rect 3662 36760 3667 36816
rect 0 36758 3667 36760
rect 0 36728 800 36758
rect 3601 36755 3667 36758
rect 43200 36728 44000 36848
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 14457 36410 14523 36413
rect 18229 36410 18295 36413
rect 14457 36408 18295 36410
rect 14457 36352 14462 36408
rect 14518 36352 18234 36408
rect 18290 36352 18295 36408
rect 14457 36350 18295 36352
rect 14457 36347 14523 36350
rect 18229 36347 18295 36350
rect 0 36138 800 36168
rect 2865 36138 2931 36141
rect 0 36136 2931 36138
rect 0 36080 2870 36136
rect 2926 36080 2931 36136
rect 0 36078 2931 36080
rect 0 36048 800 36078
rect 2865 36075 2931 36078
rect 41321 36138 41387 36141
rect 43200 36138 44000 36168
rect 41321 36136 44000 36138
rect 41321 36080 41326 36136
rect 41382 36080 44000 36136
rect 41321 36078 44000 36080
rect 41321 36075 41387 36078
rect 43200 36048 44000 36078
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 39389 35458 39455 35461
rect 43200 35458 44000 35488
rect 39389 35456 44000 35458
rect 39389 35400 39394 35456
rect 39450 35400 44000 35456
rect 39389 35398 44000 35400
rect 39389 35395 39455 35398
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 43200 35368 44000 35398
rect 34928 35327 35248 35328
rect 19568 34848 19888 34849
rect 0 34688 800 34808
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 41873 34778 41939 34781
rect 43200 34778 44000 34808
rect 41873 34776 44000 34778
rect 41873 34720 41878 34776
rect 41934 34720 44000 34776
rect 41873 34718 44000 34720
rect 41873 34715 41939 34718
rect 43200 34688 44000 34718
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 0 34008 800 34128
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 0 33328 800 33448
rect 41321 33418 41387 33421
rect 43200 33418 44000 33448
rect 41321 33416 44000 33418
rect 41321 33360 41326 33416
rect 41382 33360 44000 33416
rect 41321 33358 44000 33360
rect 41321 33355 41387 33358
rect 43200 33328 44000 33358
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 0 32648 800 32768
rect 42149 32738 42215 32741
rect 43200 32738 44000 32768
rect 42149 32736 44000 32738
rect 42149 32680 42154 32736
rect 42210 32680 44000 32736
rect 42149 32678 44000 32680
rect 42149 32675 42215 32678
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 43200 32648 44000 32678
rect 19568 32607 19888 32608
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 41321 32058 41387 32061
rect 43200 32058 44000 32088
rect 41321 32056 44000 32058
rect 41321 32000 41326 32056
rect 41382 32000 44000 32056
rect 41321 31998 44000 32000
rect 41321 31995 41387 31998
rect 43200 31968 44000 31998
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 0 31288 800 31408
rect 43200 31288 44000 31408
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 0 30608 800 30728
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 0 29928 800 30048
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 43200 29928 44000 30048
rect 34928 29887 35248 29888
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 42057 29338 42123 29341
rect 43200 29338 44000 29368
rect 42057 29336 44000 29338
rect 42057 29280 42062 29336
rect 42118 29280 44000 29336
rect 42057 29278 44000 29280
rect 42057 29275 42123 29278
rect 43200 29248 44000 29278
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 0 28658 800 28688
rect 2773 28658 2839 28661
rect 29177 28658 29243 28661
rect 0 28656 2839 28658
rect 0 28600 2778 28656
rect 2834 28600 2839 28656
rect 0 28598 2839 28600
rect 0 28568 800 28598
rect 2773 28595 2839 28598
rect 29134 28656 29243 28658
rect 29134 28600 29182 28656
rect 29238 28600 29243 28656
rect 29134 28595 29243 28600
rect 41321 28658 41387 28661
rect 43200 28658 44000 28688
rect 41321 28656 44000 28658
rect 41321 28600 41326 28656
rect 41382 28600 44000 28656
rect 41321 28598 44000 28600
rect 41321 28595 41387 28598
rect 29134 28389 29194 28595
rect 43200 28568 44000 28598
rect 29085 28384 29194 28389
rect 29085 28328 29090 28384
rect 29146 28328 29194 28384
rect 29085 28326 29194 28328
rect 29085 28323 29151 28326
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 0 27888 800 28008
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 0 27208 800 27328
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 43200 27208 44000 27328
rect 19568 27167 19888 27168
rect 4208 26688 4528 26689
rect 0 26528 800 26648
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 43200 26528 44000 26648
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 41321 25938 41387 25941
rect 43200 25938 44000 25968
rect 41321 25936 44000 25938
rect 41321 25880 41326 25936
rect 41382 25880 44000 25936
rect 41321 25878 44000 25880
rect 41321 25875 41387 25878
rect 43200 25848 44000 25878
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 0 25168 800 25288
rect 41229 25258 41295 25261
rect 43200 25258 44000 25288
rect 41229 25256 44000 25258
rect 41229 25200 41234 25256
rect 41290 25200 44000 25256
rect 41229 25198 44000 25200
rect 41229 25195 41295 25198
rect 43200 25168 44000 25198
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 0 24488 800 24608
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 5625 24306 5691 24309
rect 37549 24306 37615 24309
rect 5625 24304 37615 24306
rect 5625 24248 5630 24304
rect 5686 24248 37554 24304
rect 37610 24248 37615 24304
rect 5625 24246 37615 24248
rect 5625 24243 5691 24246
rect 37549 24243 37615 24246
rect 19568 23968 19888 23969
rect 0 23808 800 23928
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 41321 23898 41387 23901
rect 43200 23898 44000 23928
rect 41321 23896 44000 23898
rect 41321 23840 41326 23896
rect 41382 23840 44000 23896
rect 41321 23838 44000 23840
rect 41321 23835 41387 23838
rect 43200 23808 44000 23838
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 0 23128 800 23248
rect 41873 23218 41939 23221
rect 43200 23218 44000 23248
rect 41873 23216 44000 23218
rect 41873 23160 41878 23216
rect 41934 23160 44000 23216
rect 41873 23158 44000 23160
rect 41873 23155 41939 23158
rect 43200 23128 44000 23158
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 42149 22538 42215 22541
rect 43200 22538 44000 22568
rect 42149 22536 44000 22538
rect 42149 22480 42154 22536
rect 42210 22480 44000 22536
rect 42149 22478 44000 22480
rect 42149 22475 42215 22478
rect 43200 22448 44000 22478
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 27797 22130 27863 22133
rect 28901 22130 28967 22133
rect 27797 22128 28967 22130
rect 27797 22072 27802 22128
rect 27858 22072 28906 22128
rect 28962 22072 28967 22128
rect 27797 22070 28967 22072
rect 27797 22067 27863 22070
rect 28901 22067 28967 22070
rect 0 21858 800 21888
rect 1853 21858 1919 21861
rect 0 21856 1919 21858
rect 0 21800 1858 21856
rect 1914 21800 1919 21856
rect 0 21798 1919 21800
rect 0 21768 800 21798
rect 1853 21795 1919 21798
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 43200 21768 44000 21888
rect 19568 21727 19888 21728
rect 4208 21248 4528 21249
rect 0 21178 800 21208
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 2773 21178 2839 21181
rect 0 21176 2839 21178
rect 0 21120 2778 21176
rect 2834 21120 2839 21176
rect 0 21118 2839 21120
rect 0 21088 800 21118
rect 2773 21115 2839 21118
rect 14825 20906 14891 20909
rect 16573 20906 16639 20909
rect 17585 20906 17651 20909
rect 14825 20904 17651 20906
rect 14825 20848 14830 20904
rect 14886 20848 16578 20904
rect 16634 20848 17590 20904
rect 17646 20848 17651 20904
rect 14825 20846 17651 20848
rect 14825 20843 14891 20846
rect 16573 20843 16639 20846
rect 17585 20843 17651 20846
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 0 20408 800 20528
rect 39573 20498 39639 20501
rect 43200 20498 44000 20528
rect 39573 20496 44000 20498
rect 39573 20440 39578 20496
rect 39634 20440 44000 20496
rect 39573 20438 44000 20440
rect 39573 20435 39639 20438
rect 43200 20408 44000 20438
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 0 19818 800 19848
rect 1853 19818 1919 19821
rect 0 19816 1919 19818
rect 0 19760 1858 19816
rect 1914 19760 1919 19816
rect 0 19758 1919 19760
rect 0 19728 800 19758
rect 1853 19755 1919 19758
rect 42149 19818 42215 19821
rect 43200 19818 44000 19848
rect 42149 19816 44000 19818
rect 42149 19760 42154 19816
rect 42210 19760 44000 19816
rect 42149 19758 44000 19760
rect 42149 19755 42215 19758
rect 43200 19728 44000 19758
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 41229 19138 41295 19141
rect 43200 19138 44000 19168
rect 41229 19136 44000 19138
rect 41229 19080 41234 19136
rect 41290 19080 44000 19136
rect 41229 19078 44000 19080
rect 41229 19075 41295 19078
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 43200 19048 44000 19078
rect 34928 19007 35248 19008
rect 19568 18528 19888 18529
rect 0 18368 800 18488
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 41321 18458 41387 18461
rect 43200 18458 44000 18488
rect 41321 18456 44000 18458
rect 41321 18400 41326 18456
rect 41382 18400 44000 18456
rect 41321 18398 44000 18400
rect 41321 18395 41387 18398
rect 43200 18368 44000 18398
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 0 17778 800 17808
rect 2773 17778 2839 17781
rect 0 17776 2839 17778
rect 0 17720 2778 17776
rect 2834 17720 2839 17776
rect 0 17718 2839 17720
rect 0 17688 800 17718
rect 2773 17715 2839 17718
rect 13261 17642 13327 17645
rect 15285 17642 15351 17645
rect 15837 17642 15903 17645
rect 13261 17640 15903 17642
rect 13261 17584 13266 17640
rect 13322 17584 15290 17640
rect 15346 17584 15842 17640
rect 15898 17584 15903 17640
rect 13261 17582 15903 17584
rect 13261 17579 13327 17582
rect 15285 17579 15351 17582
rect 15837 17579 15903 17582
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 0 17008 800 17128
rect 43200 17008 44000 17128
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 0 16418 800 16448
rect 1853 16418 1919 16421
rect 0 16416 1919 16418
rect 0 16360 1858 16416
rect 1914 16360 1919 16416
rect 0 16358 1919 16360
rect 0 16328 800 16358
rect 1853 16355 1919 16358
rect 41689 16418 41755 16421
rect 43200 16418 44000 16448
rect 41689 16416 44000 16418
rect 41689 16360 41694 16416
rect 41750 16360 44000 16416
rect 41689 16358 44000 16360
rect 41689 16355 41755 16358
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 43200 16328 44000 16358
rect 19568 16287 19888 16288
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 42149 15738 42215 15741
rect 43200 15738 44000 15768
rect 42149 15736 44000 15738
rect 42149 15680 42154 15736
rect 42210 15680 44000 15736
rect 42149 15678 44000 15680
rect 42149 15675 42215 15678
rect 43200 15648 44000 15678
rect 14273 15602 14339 15605
rect 16113 15602 16179 15605
rect 14273 15600 16179 15602
rect 14273 15544 14278 15600
rect 14334 15544 16118 15600
rect 16174 15544 16179 15600
rect 14273 15542 16179 15544
rect 14273 15539 14339 15542
rect 16113 15539 16179 15542
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 0 15058 800 15088
rect 2773 15058 2839 15061
rect 0 15056 2839 15058
rect 0 15000 2778 15056
rect 2834 15000 2839 15056
rect 0 14998 2839 15000
rect 0 14968 800 14998
rect 2773 14995 2839 14998
rect 41321 15058 41387 15061
rect 43200 15058 44000 15088
rect 41321 15056 44000 15058
rect 41321 15000 41326 15056
rect 41382 15000 44000 15056
rect 41321 14998 44000 15000
rect 41321 14995 41387 14998
rect 43200 14968 44000 14998
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 0 14288 800 14408
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 0 13698 800 13728
rect 2865 13698 2931 13701
rect 0 13696 2931 13698
rect 0 13640 2870 13696
rect 2926 13640 2931 13696
rect 0 13638 2931 13640
rect 0 13608 800 13638
rect 2865 13635 2931 13638
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 43200 13608 44000 13728
rect 34928 13567 35248 13568
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 41321 13018 41387 13021
rect 43200 13018 44000 13048
rect 41321 13016 44000 13018
rect 41321 12960 41326 13016
rect 41382 12960 44000 13016
rect 41321 12958 44000 12960
rect 41321 12955 41387 12958
rect 43200 12928 44000 12958
rect 11697 12882 11763 12885
rect 41413 12882 41479 12885
rect 11697 12880 41479 12882
rect 11697 12824 11702 12880
rect 11758 12824 41418 12880
rect 41474 12824 41479 12880
rect 11697 12822 41479 12824
rect 11697 12819 11763 12822
rect 41413 12819 41479 12822
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 0 12338 800 12368
rect 2773 12338 2839 12341
rect 0 12336 2839 12338
rect 0 12280 2778 12336
rect 2834 12280 2839 12336
rect 0 12278 2839 12280
rect 0 12248 800 12278
rect 2773 12275 2839 12278
rect 42149 12338 42215 12341
rect 43200 12338 44000 12368
rect 42149 12336 44000 12338
rect 42149 12280 42154 12336
rect 42210 12280 44000 12336
rect 42149 12278 44000 12280
rect 42149 12275 42215 12278
rect 43200 12248 44000 12278
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 0 11568 800 11688
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 0 10888 800 11008
rect 42149 10978 42215 10981
rect 43200 10978 44000 11008
rect 42149 10976 44000 10978
rect 42149 10920 42154 10976
rect 42210 10920 44000 10976
rect 42149 10918 44000 10920
rect 42149 10915 42215 10918
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 43200 10888 44000 10918
rect 19568 10847 19888 10848
rect 4208 10368 4528 10369
rect 0 10298 800 10328
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 2773 10298 2839 10301
rect 0 10296 2839 10298
rect 0 10240 2778 10296
rect 2834 10240 2839 10296
rect 0 10238 2839 10240
rect 0 10208 800 10238
rect 2773 10235 2839 10238
rect 42149 10298 42215 10301
rect 43200 10298 44000 10328
rect 42149 10296 44000 10298
rect 42149 10240 42154 10296
rect 42210 10240 44000 10296
rect 42149 10238 44000 10240
rect 42149 10235 42215 10238
rect 43200 10208 44000 10238
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 43200 9528 44000 9648
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 0 8938 800 8968
rect 1393 8938 1459 8941
rect 0 8936 1459 8938
rect 0 8880 1398 8936
rect 1454 8880 1459 8936
rect 0 8878 1459 8880
rect 0 8848 800 8878
rect 1393 8875 1459 8878
rect 43200 8848 44000 8968
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 0 8258 800 8288
rect 2773 8258 2839 8261
rect 0 8256 2839 8258
rect 0 8200 2778 8256
rect 2834 8200 2839 8256
rect 0 8198 2839 8200
rect 0 8168 800 8198
rect 2773 8195 2839 8198
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 19568 7648 19888 7649
rect 0 7488 800 7608
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 43200 7488 44000 7608
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 0 6898 800 6928
rect 4061 6898 4127 6901
rect 0 6896 4127 6898
rect 0 6840 4066 6896
rect 4122 6840 4127 6896
rect 0 6838 4127 6840
rect 0 6808 800 6838
rect 4061 6835 4127 6838
rect 41873 6898 41939 6901
rect 43200 6898 44000 6928
rect 41873 6896 44000 6898
rect 41873 6840 41878 6896
rect 41934 6840 44000 6896
rect 41873 6838 44000 6840
rect 41873 6835 41939 6838
rect 43200 6808 44000 6838
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 42149 6218 42215 6221
rect 43200 6218 44000 6248
rect 42149 6216 44000 6218
rect 42149 6160 42154 6216
rect 42210 6160 44000 6216
rect 42149 6158 44000 6160
rect 42149 6155 42215 6158
rect 43200 6128 44000 6158
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 0 5538 800 5568
rect 1853 5538 1919 5541
rect 0 5536 1919 5538
rect 0 5480 1858 5536
rect 1914 5480 1919 5536
rect 0 5478 1919 5480
rect 0 5448 800 5478
rect 1853 5475 1919 5478
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 43200 5448 44000 5568
rect 19568 5407 19888 5408
rect 4208 4928 4528 4929
rect 0 4858 800 4888
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 2773 4858 2839 4861
rect 0 4856 2839 4858
rect 0 4800 2778 4856
rect 2834 4800 2839 4856
rect 0 4798 2839 4800
rect 0 4768 800 4798
rect 2773 4795 2839 4798
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 0 4178 800 4208
rect 3141 4178 3207 4181
rect 0 4176 3207 4178
rect 0 4120 3146 4176
rect 3202 4120 3207 4176
rect 0 4118 3207 4120
rect 0 4088 800 4118
rect 3141 4115 3207 4118
rect 41321 4178 41387 4181
rect 43200 4178 44000 4208
rect 41321 4176 44000 4178
rect 41321 4120 41326 4176
rect 41382 4120 44000 4176
rect 41321 4118 44000 4120
rect 41321 4115 41387 4118
rect 43200 4088 44000 4118
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 0 3498 800 3528
rect 1393 3498 1459 3501
rect 0 3496 1459 3498
rect 0 3440 1398 3496
rect 1454 3440 1459 3496
rect 0 3438 1459 3440
rect 0 3408 800 3438
rect 1393 3435 1459 3438
rect 43200 3408 44000 3528
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 43200 2728 44000 2848
rect 34928 2687 35248 2688
rect 19568 2208 19888 2209
rect 0 2138 800 2168
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 3417 2138 3483 2141
rect 0 2136 3483 2138
rect 0 2080 3422 2136
rect 3478 2080 3483 2136
rect 0 2078 3483 2080
rect 0 2048 800 2078
rect 3417 2075 3483 2078
rect 39941 2138 40007 2141
rect 43200 2138 44000 2168
rect 39941 2136 44000 2138
rect 39941 2080 39946 2136
rect 40002 2080 44000 2136
rect 39941 2078 44000 2080
rect 39941 2075 40007 2078
rect 43200 2048 44000 2078
rect 0 1458 800 1488
rect 2773 1458 2839 1461
rect 0 1456 2839 1458
rect 0 1400 2778 1456
rect 2834 1400 2839 1456
rect 0 1398 2839 1400
rect 0 1368 800 1398
rect 2773 1395 2839 1398
rect 0 688 800 808
rect 39757 778 39823 781
rect 43200 778 44000 808
rect 39757 776 44000 778
rect 39757 720 39762 776
rect 39818 720 44000 776
rect 39757 718 44000 720
rect 39757 715 39823 718
rect 43200 688 44000 718
rect 41321 98 41387 101
rect 43200 98 44000 128
rect 41321 96 44000 98
rect 41321 40 41326 96
rect 41382 40 44000 96
rect 41321 38 44000 40
rect 41321 35 41387 38
rect 43200 8 44000 38
<< via3 >>
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 40832 4528 41392
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 41376 19888 41392
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 40832 35248 41392
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__decap_6  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2208 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2944 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50
timestamp 1644511149
transform 1 0 5704 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78
timestamp 1644511149
transform 1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1644511149
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_116 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11776 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_128
timestamp 1644511149
transform 1 0 12880 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_149 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_155
timestamp 1644511149
transform 1 0 15364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1644511149
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_181
timestamp 1644511149
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1644511149
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_209
timestamp 1644511149
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1644511149
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_246
timestamp 1644511149
transform 1 0 23736 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_265
timestamp 1644511149
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1644511149
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_289
timestamp 1644511149
transform 1 0 27692 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_293
timestamp 1644511149
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1644511149
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_309
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_321
timestamp 1644511149
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1644511149
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_349
timestamp 1644511149
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1644511149
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_373
timestamp 1644511149
transform 1 0 35420 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_379
timestamp 1644511149
transform 1 0 35972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_386
timestamp 1644511149
transform 1 0 36616 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_416
timestamp 1644511149
transform 1 0 39376 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_421
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_444
timestamp 1644511149
transform 1 0 41952 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_449
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_24
timestamp 1644511149
transform 1 0 3312 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_49
timestamp 1644511149
transform 1 0 5612 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1644511149
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_60
timestamp 1644511149
transform 1 0 6624 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_87
timestamp 1644511149
transform 1 0 9108 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_95
timestamp 1644511149
transform 1 0 9844 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_100
timestamp 1644511149
transform 1 0 10304 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_104
timestamp 1644511149
transform 1 0 10672 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1644511149
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_134
timestamp 1644511149
transform 1 0 13432 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_142
timestamp 1644511149
transform 1 0 14168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1644511149
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_172
timestamp 1644511149
transform 1 0 16928 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_184
timestamp 1644511149
transform 1 0 18032 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_206
timestamp 1644511149
transform 1 0 20056 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_213
timestamp 1644511149
transform 1 0 20700 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_221
timestamp 1644511149
transform 1 0 21436 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_229
timestamp 1644511149
transform 1 0 22172 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_233
timestamp 1644511149
transform 1 0 22540 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_237
timestamp 1644511149
transform 1 0 22908 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_264
timestamp 1644511149
transform 1 0 25392 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1644511149
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_289
timestamp 1644511149
transform 1 0 27692 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_311
timestamp 1644511149
transform 1 0 29716 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_323
timestamp 1644511149
transform 1 0 30820 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1644511149
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_349
timestamp 1644511149
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_361
timestamp 1644511149
transform 1 0 34316 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_388
timestamp 1644511149
transform 1 0 36800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_393
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_417
timestamp 1644511149
transform 1 0 39468 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_442
timestamp 1644511149
transform 1 0 41768 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_449
timestamp 1644511149
transform 1 0 42412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1644511149
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_29
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_35
timestamp 1644511149
transform 1 0 4324 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_60
timestamp 1644511149
transform 1 0 6624 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_66
timestamp 1644511149
transform 1 0 7176 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_70
timestamp 1644511149
transform 1 0 7544 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_74
timestamp 1644511149
transform 1 0 7912 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_78
timestamp 1644511149
transform 1 0 8280 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_107
timestamp 1644511149
transform 1 0 10948 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_132
timestamp 1644511149
transform 1 0 13248 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_152
timestamp 1644511149
transform 1 0 15088 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_159
timestamp 1644511149
transform 1 0 15732 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_184
timestamp 1644511149
transform 1 0 18032 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_191
timestamp 1644511149
transform 1 0 18676 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1644511149
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_221
timestamp 1644511149
transform 1 0 21436 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_229
timestamp 1644511149
transform 1 0 22172 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_233
timestamp 1644511149
transform 1 0 22540 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_240
timestamp 1644511149
transform 1 0 23184 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_247
timestamp 1644511149
transform 1 0 23828 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1644511149
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_265
timestamp 1644511149
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_277
timestamp 1644511149
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_289
timestamp 1644511149
transform 1 0 27692 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_293
timestamp 1644511149
transform 1 0 28060 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_305
timestamp 1644511149
transform 1 0 29164 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_321
timestamp 1644511149
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_333
timestamp 1644511149
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_345
timestamp 1644511149
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1644511149
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1644511149
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_386
timestamp 1644511149
transform 1 0 36616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_411
timestamp 1644511149
transform 1 0 38916 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1644511149
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_421
timestamp 1644511149
transform 1 0 39836 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_425
timestamp 1644511149
transform 1 0 40204 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_447
timestamp 1644511149
transform 1 0 42228 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_12
timestamp 1644511149
transform 1 0 2208 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_20
timestamp 1644511149
transform 1 0 2944 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_43
timestamp 1644511149
transform 1 0 5060 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_50
timestamp 1644511149
transform 1 0 5704 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_60
timestamp 1644511149
transform 1 0 6624 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_72
timestamp 1644511149
transform 1 0 7728 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_84
timestamp 1644511149
transform 1 0 8832 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_91
timestamp 1644511149
transform 1 0 9476 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_98
timestamp 1644511149
transform 1 0 10120 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_104
timestamp 1644511149
transform 1 0 10672 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 1644511149
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_116
timestamp 1644511149
transform 1 0 11776 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_128
timestamp 1644511149
transform 1 0 12880 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_140
timestamp 1644511149
transform 1 0 13984 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_152
timestamp 1644511149
transform 1 0 15088 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1644511149
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_181
timestamp 1644511149
transform 1 0 17756 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_188
timestamp 1644511149
transform 1 0 18400 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_200
timestamp 1644511149
transform 1 0 19504 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_204
timestamp 1644511149
transform 1 0 19872 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_216
timestamp 1644511149
transform 1 0 20976 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_229
timestamp 1644511149
transform 1 0 22172 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_233
timestamp 1644511149
transform 1 0 22540 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_255
timestamp 1644511149
transform 1 0 24564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_267
timestamp 1644511149
transform 1 0 25668 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1644511149
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_305
timestamp 1644511149
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_317
timestamp 1644511149
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1644511149
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1644511149
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_349
timestamp 1644511149
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_361
timestamp 1644511149
transform 1 0 34316 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_366
timestamp 1644511149
transform 1 0 34776 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_374
timestamp 1644511149
transform 1 0 35512 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_378
timestamp 1644511149
transform 1 0 35880 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_384
timestamp 1644511149
transform 1 0 36432 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_388
timestamp 1644511149
transform 1 0 36800 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_402
timestamp 1644511149
transform 1 0 38088 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_406
timestamp 1644511149
transform 1 0 38456 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_410
timestamp 1644511149
transform 1 0 38824 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_439
timestamp 1644511149
transform 1 0 41492 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1644511149
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_449
timestamp 1644511149
transform 1 0 42412 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_6
timestamp 1644511149
transform 1 0 1656 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_13
timestamp 1644511149
transform 1 0 2300 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_20
timestamp 1644511149
transform 1 0 2944 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_32
timestamp 1644511149
transform 1 0 4048 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_39
timestamp 1644511149
transform 1 0 4692 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_46
timestamp 1644511149
transform 1 0 5336 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_58
timestamp 1644511149
transform 1 0 6440 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_70
timestamp 1644511149
transform 1 0 7544 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1644511149
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_97
timestamp 1644511149
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_109
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_121
timestamp 1644511149
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1644511149
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1644511149
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1644511149
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_209
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_221
timestamp 1644511149
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_233
timestamp 1644511149
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1644511149
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1644511149
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_277
timestamp 1644511149
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_289
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1644511149
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1644511149
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_345
timestamp 1644511149
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1644511149
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_388
timestamp 1644511149
transform 1 0 36800 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_396
timestamp 1644511149
transform 1 0 37536 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_402
timestamp 1644511149
transform 1 0 38088 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_409
timestamp 1644511149
transform 1 0 38732 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_416
timestamp 1644511149
transform 1 0 39376 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_421
timestamp 1644511149
transform 1 0 39836 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_425
timestamp 1644511149
transform 1 0 40204 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_447
timestamp 1644511149
transform 1 0 42228 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_30
timestamp 1644511149
transform 1 0 3864 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_37
timestamp 1644511149
transform 1 0 4508 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_49
timestamp 1644511149
transform 1 0 5612 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_193
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_205
timestamp 1644511149
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1644511149
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_249
timestamp 1644511149
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_261
timestamp 1644511149
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1644511149
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_373
timestamp 1644511149
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1644511149
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_405
timestamp 1644511149
transform 1 0 38364 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_427
timestamp 1644511149
transform 1 0 40388 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_434
timestamp 1644511149
transform 1 0 41032 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1644511149
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1644511149
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_449
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1644511149
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_32
timestamp 1644511149
transform 1 0 4048 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_39
timestamp 1644511149
transform 1 0 4692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_51
timestamp 1644511149
transform 1 0 5796 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_63
timestamp 1644511149
transform 1 0 6900 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_75
timestamp 1644511149
transform 1 0 8004 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_397
timestamp 1644511149
transform 1 0 37628 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_402
timestamp 1644511149
transform 1 0 38088 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_406
timestamp 1644511149
transform 1 0 38456 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_410
timestamp 1644511149
transform 1 0 38824 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_418
timestamp 1644511149
transform 1 0 39560 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_424
timestamp 1644511149
transform 1 0 40112 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_433
timestamp 1644511149
transform 1 0 40940 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_440
timestamp 1644511149
transform 1 0 41584 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_447
timestamp 1644511149
transform 1 0 42228 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_6
timestamp 1644511149
transform 1 0 1656 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_13
timestamp 1644511149
transform 1 0 2300 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_20
timestamp 1644511149
transform 1 0 2944 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_28
timestamp 1644511149
transform 1 0 3680 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 1644511149
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_417
timestamp 1644511149
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_429
timestamp 1644511149
transform 1 0 40572 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_436
timestamp 1644511149
transform 1 0 41216 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_443
timestamp 1644511149
transform 1 0 41860 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1644511149
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_449
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_35
timestamp 1644511149
transform 1 0 4324 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_47
timestamp 1644511149
transform 1 0 5428 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_59
timestamp 1644511149
transform 1 0 6532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_71
timestamp 1644511149
transform 1 0 7636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_205
timestamp 1644511149
transform 1 0 19964 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_211
timestamp 1644511149
transform 1 0 20516 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_223
timestamp 1644511149
transform 1 0 21620 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_235
timestamp 1644511149
transform 1 0 22724 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_247
timestamp 1644511149
transform 1 0 23828 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_389
timestamp 1644511149
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_401
timestamp 1644511149
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1644511149
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1644511149
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_421
timestamp 1644511149
transform 1 0 39836 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_425
timestamp 1644511149
transform 1 0 40204 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_447
timestamp 1644511149
transform 1 0 42228 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1644511149
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_173
timestamp 1644511149
transform 1 0 17020 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_178
timestamp 1644511149
transform 1 0 17480 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_193
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_215
timestamp 1644511149
transform 1 0 20884 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_254
timestamp 1644511149
transform 1 0 24472 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_266
timestamp 1644511149
transform 1 0 25576 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp 1644511149
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_317
timestamp 1644511149
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1644511149
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_361
timestamp 1644511149
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1644511149
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_417
timestamp 1644511149
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_429
timestamp 1644511149
transform 1 0 40572 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_436
timestamp 1644511149
transform 1 0 41216 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_444
timestamp 1644511149
transform 1 0 41952 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_449
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1644511149
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_187
timestamp 1644511149
transform 1 0 18308 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_213
timestamp 1644511149
transform 1 0 20700 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_233
timestamp 1644511149
transform 1 0 22540 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_240
timestamp 1644511149
transform 1 0 23184 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_247
timestamp 1644511149
transform 1 0 23828 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_261
timestamp 1644511149
transform 1 0 25116 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_280
timestamp 1644511149
transform 1 0 26864 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_292
timestamp 1644511149
transform 1 0 27968 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_304
timestamp 1644511149
transform 1 0 29072 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_345
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1644511149
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_401
timestamp 1644511149
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1644511149
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1644511149
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_433
timestamp 1644511149
transform 1 0 40940 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_442
timestamp 1644511149
transform 1 0 41768 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_450
timestamp 1644511149
transform 1 0 42504 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_28
timestamp 1644511149
transform 1 0 3680 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_40
timestamp 1644511149
transform 1 0 4784 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1644511149
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_145
timestamp 1644511149
transform 1 0 14444 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_164
timestamp 1644511149
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_179
timestamp 1644511149
transform 1 0 17572 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_185
timestamp 1644511149
transform 1 0 18124 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_192
timestamp 1644511149
transform 1 0 18768 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_207
timestamp 1644511149
transform 1 0 20148 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_230
timestamp 1644511149
transform 1 0 22264 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_254
timestamp 1644511149
transform 1 0 24472 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_266
timestamp 1644511149
transform 1 0 25576 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp 1644511149
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_300
timestamp 1644511149
transform 1 0 28704 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_320
timestamp 1644511149
transform 1 0 30544 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_330
timestamp 1644511149
transform 1 0 31464 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_373
timestamp 1644511149
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1644511149
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1644511149
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_417
timestamp 1644511149
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_429
timestamp 1644511149
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1644511149
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1644511149
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_449
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1644511149
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_159
timestamp 1644511149
transform 1 0 15732 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_168
timestamp 1644511149
transform 1 0 16560 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_180
timestamp 1644511149
transform 1 0 17664 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_186
timestamp 1644511149
transform 1 0 18216 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1644511149
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_201
timestamp 1644511149
transform 1 0 19596 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_207
timestamp 1644511149
transform 1 0 20148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_224
timestamp 1644511149
transform 1 0 21712 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_233
timestamp 1644511149
transform 1 0 22540 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_242
timestamp 1644511149
transform 1 0 23368 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1644511149
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_271
timestamp 1644511149
transform 1 0 26036 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_277
timestamp 1644511149
transform 1 0 26588 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_284
timestamp 1644511149
transform 1 0 27232 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_304
timestamp 1644511149
transform 1 0 29072 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_317
timestamp 1644511149
transform 1 0 30268 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_329
timestamp 1644511149
transform 1 0 31372 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_346
timestamp 1644511149
transform 1 0 32936 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_358
timestamp 1644511149
transform 1 0 34040 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1644511149
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1644511149
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_433
timestamp 1644511149
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_445
timestamp 1644511149
transform 1 0 42044 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_7
timestamp 1644511149
transform 1 0 1748 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_14
timestamp 1644511149
transform 1 0 2392 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_21
timestamp 1644511149
transform 1 0 3036 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_33
timestamp 1644511149
transform 1 0 4140 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_45
timestamp 1644511149
transform 1 0 5244 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_53
timestamp 1644511149
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_191
timestamp 1644511149
transform 1 0 18676 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_203
timestamp 1644511149
transform 1 0 19780 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_215
timestamp 1644511149
transform 1 0 20884 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_230
timestamp 1644511149
transform 1 0 22264 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_257
timestamp 1644511149
transform 1 0 24748 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_267
timestamp 1644511149
transform 1 0 25668 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_276
timestamp 1644511149
transform 1 0 26496 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_284
timestamp 1644511149
transform 1 0 27232 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_290
timestamp 1644511149
transform 1 0 27784 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_307
timestamp 1644511149
transform 1 0 29348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_313
timestamp 1644511149
transform 1 0 29900 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_323
timestamp 1644511149
transform 1 0 30820 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_340
timestamp 1644511149
transform 1 0 32384 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_348
timestamp 1644511149
transform 1 0 33120 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_358
timestamp 1644511149
transform 1 0 34040 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_370
timestamp 1644511149
transform 1 0 35144 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_382
timestamp 1644511149
transform 1 0 36248 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_390
timestamp 1644511149
transform 1 0 36984 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_417
timestamp 1644511149
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_429
timestamp 1644511149
transform 1 0 40572 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_440
timestamp 1644511149
transform 1 0 41584 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_449
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_12
timestamp 1644511149
transform 1 0 2208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_19
timestamp 1644511149
transform 1 0 2852 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_161
timestamp 1644511149
transform 1 0 15916 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_170
timestamp 1644511149
transform 1 0 16744 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_192
timestamp 1644511149
transform 1 0 18768 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_205
timestamp 1644511149
transform 1 0 19964 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_217
timestamp 1644511149
transform 1 0 21068 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_223
timestamp 1644511149
transform 1 0 21620 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_227
timestamp 1644511149
transform 1 0 21988 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_234
timestamp 1644511149
transform 1 0 22632 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_241
timestamp 1644511149
transform 1 0 23276 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_249
timestamp 1644511149
transform 1 0 24012 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_261
timestamp 1644511149
transform 1 0 25116 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_281
timestamp 1644511149
transform 1 0 26956 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1644511149
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1644511149
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_313
timestamp 1644511149
transform 1 0 29900 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_330
timestamp 1644511149
transform 1 0 31464 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_351
timestamp 1644511149
transform 1 0 33396 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_372
timestamp 1644511149
transform 1 0 35328 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_380
timestamp 1644511149
transform 1 0 36064 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_392
timestamp 1644511149
transform 1 0 37168 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_404
timestamp 1644511149
transform 1 0 38272 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_416
timestamp 1644511149
transform 1 0 39376 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_421
timestamp 1644511149
transform 1 0 39836 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_425
timestamp 1644511149
transform 1 0 40204 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_447
timestamp 1644511149
transform 1 0 42228 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1644511149
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_145
timestamp 1644511149
transform 1 0 14444 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1644511149
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_179
timestamp 1644511149
transform 1 0 17572 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_190
timestamp 1644511149
transform 1 0 18584 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_200
timestamp 1644511149
transform 1 0 19504 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_220
timestamp 1644511149
transform 1 0 21344 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_233
timestamp 1644511149
transform 1 0 22540 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_241
timestamp 1644511149
transform 1 0 23276 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_248
timestamp 1644511149
transform 1 0 23920 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_268
timestamp 1644511149
transform 1 0 25760 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_325
timestamp 1644511149
transform 1 0 31004 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_332
timestamp 1644511149
transform 1 0 31648 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_350
timestamp 1644511149
transform 1 0 33304 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_362
timestamp 1644511149
transform 1 0 34408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_372
timestamp 1644511149
transform 1 0 35328 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_384
timestamp 1644511149
transform 1 0 36432 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_417
timestamp 1644511149
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_429
timestamp 1644511149
transform 1 0 40572 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_433
timestamp 1644511149
transform 1 0 40940 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_440
timestamp 1644511149
transform 1 0 41584 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_449
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_9
timestamp 1644511149
transform 1 0 1932 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_21
timestamp 1644511149
transform 1 0 3036 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_191
timestamp 1644511149
transform 1 0 18676 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_206
timestamp 1644511149
transform 1 0 20056 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_214
timestamp 1644511149
transform 1 0 20792 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_219
timestamp 1644511149
transform 1 0 21252 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_226
timestamp 1644511149
transform 1 0 21896 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_238
timestamp 1644511149
transform 1 0 23000 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1644511149
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_265
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_275
timestamp 1644511149
transform 1 0 26404 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_287
timestamp 1644511149
transform 1 0 27508 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_299
timestamp 1644511149
transform 1 0 28612 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_349
timestamp 1644511149
transform 1 0 33212 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_358
timestamp 1644511149
transform 1 0 34040 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_370
timestamp 1644511149
transform 1 0 35144 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_374
timestamp 1644511149
transform 1 0 35512 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_384
timestamp 1644511149
transform 1 0 36432 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_391
timestamp 1644511149
transform 1 0 37076 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_398
timestamp 1644511149
transform 1 0 37720 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_410
timestamp 1644511149
transform 1 0 38824 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_418
timestamp 1644511149
transform 1 0 39560 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_421
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_425
timestamp 1644511149
transform 1 0 40204 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_447
timestamp 1644511149
transform 1 0 42228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_9
timestamp 1644511149
transform 1 0 1932 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_13
timestamp 1644511149
transform 1 0 2300 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_25
timestamp 1644511149
transform 1 0 3404 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_37
timestamp 1644511149
transform 1 0 4508 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_49
timestamp 1644511149
transform 1 0 5612 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_87
timestamp 1644511149
transform 1 0 9108 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_91
timestamp 1644511149
transform 1 0 9476 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_103
timestamp 1644511149
transform 1 0 10580 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_145
timestamp 1644511149
transform 1 0 14444 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_151
timestamp 1644511149
transform 1 0 14996 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_163
timestamp 1644511149
transform 1 0 16100 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_175
timestamp 1644511149
transform 1 0 17204 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_179
timestamp 1644511149
transform 1 0 17572 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_190
timestamp 1644511149
transform 1 0 18584 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_194
timestamp 1644511149
transform 1 0 18952 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_200
timestamp 1644511149
transform 1 0 19504 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_220
timestamp 1644511149
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_231
timestamp 1644511149
transform 1 0 22356 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_248
timestamp 1644511149
transform 1 0 23920 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_268
timestamp 1644511149
transform 1 0 25760 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_297
timestamp 1644511149
transform 1 0 28428 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_309
timestamp 1644511149
transform 1 0 29532 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_317
timestamp 1644511149
transform 1 0 30268 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_322
timestamp 1644511149
transform 1 0 30728 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_334
timestamp 1644511149
transform 1 0 31832 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_357
timestamp 1644511149
transform 1 0 33948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_365
timestamp 1644511149
transform 1 0 34684 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_387
timestamp 1644511149
transform 1 0 36708 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_417
timestamp 1644511149
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_429
timestamp 1644511149
transform 1 0 40572 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_434
timestamp 1644511149
transform 1 0 41032 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1644511149
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1644511149
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_449
timestamp 1644511149
transform 1 0 42412 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_24
timestamp 1644511149
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_125
timestamp 1644511149
transform 1 0 12604 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_129
timestamp 1644511149
transform 1 0 12972 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_137
timestamp 1644511149
transform 1 0 13708 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_159
timestamp 1644511149
transform 1 0 15732 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_163
timestamp 1644511149
transform 1 0 16100 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_169
timestamp 1644511149
transform 1 0 16652 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_180
timestamp 1644511149
transform 1 0 17664 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_190
timestamp 1644511149
transform 1 0 18584 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_18_200
timestamp 1644511149
transform 1 0 19504 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_206
timestamp 1644511149
transform 1 0 20056 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_212
timestamp 1644511149
transform 1 0 20608 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_220
timestamp 1644511149
transform 1 0 21344 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_232
timestamp 1644511149
transform 1 0 22448 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_244
timestamp 1644511149
transform 1 0 23552 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_258
timestamp 1644511149
transform 1 0 24840 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_270
timestamp 1644511149
transform 1 0 25944 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_287
timestamp 1644511149
transform 1 0 27508 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_295
timestamp 1644511149
transform 1 0 28244 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_304
timestamp 1644511149
transform 1 0 29072 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_313
timestamp 1644511149
transform 1 0 29900 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_327
timestamp 1644511149
transform 1 0 31188 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_344
timestamp 1644511149
transform 1 0 32752 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_360
timestamp 1644511149
transform 1 0 34224 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_370
timestamp 1644511149
transform 1 0 35144 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_378
timestamp 1644511149
transform 1 0 35880 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_384
timestamp 1644511149
transform 1 0 36432 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_391
timestamp 1644511149
transform 1 0 37076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_403
timestamp 1644511149
transform 1 0 38180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_415
timestamp 1644511149
transform 1 0 39284 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1644511149
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_421
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_425
timestamp 1644511149
transform 1 0 40204 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_447
timestamp 1644511149
transform 1 0 42228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_9
timestamp 1644511149
transform 1 0 1932 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_21
timestamp 1644511149
transform 1 0 3036 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_33
timestamp 1644511149
transform 1 0 4140 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_45
timestamp 1644511149
transform 1 0 5244 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 1644511149
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_119
timestamp 1644511149
transform 1 0 12052 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_141
timestamp 1644511149
transform 1 0 14076 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_149
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_154
timestamp 1644511149
transform 1 0 15272 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1644511149
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_179
timestamp 1644511149
transform 1 0 17572 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_203
timestamp 1644511149
transform 1 0 19780 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_211
timestamp 1644511149
transform 1 0 20516 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_219
timestamp 1644511149
transform 1 0 21252 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1644511149
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_230
timestamp 1644511149
transform 1 0 22264 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_242
timestamp 1644511149
transform 1 0 23368 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_254
timestamp 1644511149
transform 1 0 24472 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_265
timestamp 1644511149
transform 1 0 25484 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_271
timestamp 1644511149
transform 1 0 26036 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_276
timestamp 1644511149
transform 1 0 26496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_297
timestamp 1644511149
transform 1 0 28428 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_307
timestamp 1644511149
transform 1 0 29348 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_315
timestamp 1644511149
transform 1 0 30084 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_323
timestamp 1644511149
transform 1 0 30820 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_331
timestamp 1644511149
transform 1 0 31556 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_340
timestamp 1644511149
transform 1 0 32384 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_352
timestamp 1644511149
transform 1 0 33488 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_362
timestamp 1644511149
transform 1 0 34408 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_366
timestamp 1644511149
transform 1 0 34776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_375
timestamp 1644511149
transform 1 0 35604 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_387
timestamp 1644511149
transform 1 0 36708 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_401
timestamp 1644511149
transform 1 0 37996 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_413
timestamp 1644511149
transform 1 0 39100 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_425
timestamp 1644511149
transform 1 0 40204 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_434
timestamp 1644511149
transform 1 0 41032 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1644511149
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1644511149
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_449
timestamp 1644511149
transform 1 0 42412 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_9
timestamp 1644511149
transform 1 0 1932 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_13
timestamp 1644511149
transform 1 0 2300 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_20
timestamp 1644511149
transform 1 0 2944 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_117
timestamp 1644511149
transform 1 0 11868 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_128
timestamp 1644511149
transform 1 0 12880 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_161
timestamp 1644511149
transform 1 0 15916 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_171
timestamp 1644511149
transform 1 0 16836 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_185
timestamp 1644511149
transform 1 0 18124 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_193
timestamp 1644511149
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_205
timestamp 1644511149
transform 1 0 19964 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_218
timestamp 1644511149
transform 1 0 21160 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_227
timestamp 1644511149
transform 1 0 21988 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_231
timestamp 1644511149
transform 1 0 22356 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_248
timestamp 1644511149
transform 1 0 23920 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_259
timestamp 1644511149
transform 1 0 24932 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_269
timestamp 1644511149
transform 1 0 25852 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_273
timestamp 1644511149
transform 1 0 26220 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_277
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_289
timestamp 1644511149
transform 1 0 27692 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_293
timestamp 1644511149
transform 1 0 28060 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1644511149
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_318
timestamp 1644511149
transform 1 0 30360 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_337
timestamp 1644511149
transform 1 0 32108 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_345
timestamp 1644511149
transform 1 0 32844 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_355
timestamp 1644511149
transform 1 0 33764 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1644511149
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_369
timestamp 1644511149
transform 1 0 35052 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_383
timestamp 1644511149
transform 1 0 36340 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_390
timestamp 1644511149
transform 1 0 36984 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_397
timestamp 1644511149
transform 1 0 37628 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_409
timestamp 1644511149
transform 1 0 38732 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_417
timestamp 1644511149
transform 1 0 39468 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_421
timestamp 1644511149
transform 1 0 39836 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_425
timestamp 1644511149
transform 1 0 40204 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_447
timestamp 1644511149
transform 1 0 42228 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_30
timestamp 1644511149
transform 1 0 3864 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_42
timestamp 1644511149
transform 1 0 4968 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1644511149
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_157
timestamp 1644511149
transform 1 0 15548 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_165
timestamp 1644511149
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_174
timestamp 1644511149
transform 1 0 17112 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_187
timestamp 1644511149
transform 1 0 18308 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_199
timestamp 1644511149
transform 1 0 19412 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_206
timestamp 1644511149
transform 1 0 20056 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_214
timestamp 1644511149
transform 1 0 20792 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1644511149
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_229
timestamp 1644511149
transform 1 0 22172 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_249
timestamp 1644511149
transform 1 0 24012 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_253
timestamp 1644511149
transform 1 0 24380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_258
timestamp 1644511149
transform 1 0 24840 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_265
timestamp 1644511149
transform 1 0 25484 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_271
timestamp 1644511149
transform 1 0 26036 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_275
timestamp 1644511149
transform 1 0 26404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1644511149
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_291
timestamp 1644511149
transform 1 0 27876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_303
timestamp 1644511149
transform 1 0 28980 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_318
timestamp 1644511149
transform 1 0 30360 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_332
timestamp 1644511149
transform 1 0 31648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_340
timestamp 1644511149
transform 1 0 32384 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_344
timestamp 1644511149
transform 1 0 32752 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_354
timestamp 1644511149
transform 1 0 33672 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_360
timestamp 1644511149
transform 1 0 34224 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_369
timestamp 1644511149
transform 1 0 35052 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_417
timestamp 1644511149
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_429
timestamp 1644511149
transform 1 0 40572 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_437
timestamp 1644511149
transform 1 0 41308 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_443
timestamp 1644511149
transform 1 0 41860 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1644511149
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_449
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_14
timestamp 1644511149
transform 1 0 2392 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1644511149
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_117
timestamp 1644511149
transform 1 0 11868 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_123
timestamp 1644511149
transform 1 0 12420 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_131
timestamp 1644511149
transform 1 0 13156 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_135
timestamp 1644511149
transform 1 0 13524 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_152
timestamp 1644511149
transform 1 0 15088 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_163
timestamp 1644511149
transform 1 0 16100 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_175
timestamp 1644511149
transform 1 0 17204 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1644511149
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1644511149
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_202
timestamp 1644511149
transform 1 0 19688 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_214
timestamp 1644511149
transform 1 0 20792 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_227
timestamp 1644511149
transform 1 0 21988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_239
timestamp 1644511149
transform 1 0 23092 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1644511149
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1644511149
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_257
timestamp 1644511149
transform 1 0 24748 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_274
timestamp 1644511149
transform 1 0 26312 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_294
timestamp 1644511149
transform 1 0 28152 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_306
timestamp 1644511149
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_325
timestamp 1644511149
transform 1 0 31004 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_333
timestamp 1644511149
transform 1 0 31740 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_348
timestamp 1644511149
transform 1 0 33120 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_352
timestamp 1644511149
transform 1 0 33488 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_356
timestamp 1644511149
transform 1 0 33856 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_370
timestamp 1644511149
transform 1 0 35144 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_381
timestamp 1644511149
transform 1 0 36156 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_388
timestamp 1644511149
transform 1 0 36800 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_400
timestamp 1644511149
transform 1 0 37904 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_412
timestamp 1644511149
transform 1 0 39008 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_421
timestamp 1644511149
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_433
timestamp 1644511149
transform 1 0 40940 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_440
timestamp 1644511149
transform 1 0 41584 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_447
timestamp 1644511149
transform 1 0 42228 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_28
timestamp 1644511149
transform 1 0 3680 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_40
timestamp 1644511149
transform 1 0 4784 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1644511149
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_139
timestamp 1644511149
transform 1 0 13892 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_143
timestamp 1644511149
transform 1 0 14260 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_150
timestamp 1644511149
transform 1 0 14904 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_162
timestamp 1644511149
transform 1 0 16008 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_23_185
timestamp 1644511149
transform 1 0 18124 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_191
timestamp 1644511149
transform 1 0 18676 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_198
timestamp 1644511149
transform 1 0 19320 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_208
timestamp 1644511149
transform 1 0 20240 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_218
timestamp 1644511149
transform 1 0 21160 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_238
timestamp 1644511149
transform 1 0 23000 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_242
timestamp 1644511149
transform 1 0 23368 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_247
timestamp 1644511149
transform 1 0 23828 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_255
timestamp 1644511149
transform 1 0 24564 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_262
timestamp 1644511149
transform 1 0 25208 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_274
timestamp 1644511149
transform 1 0 26312 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_305
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_313
timestamp 1644511149
transform 1 0 29900 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_318
timestamp 1644511149
transform 1 0 30360 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_327
timestamp 1644511149
transform 1 0 31188 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1644511149
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_369
timestamp 1644511149
transform 1 0 35052 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_377
timestamp 1644511149
transform 1 0 35788 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_389
timestamp 1644511149
transform 1 0 36892 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_417
timestamp 1644511149
transform 1 0 39468 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_444
timestamp 1644511149
transform 1 0 41952 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_449
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_10
timestamp 1644511149
transform 1 0 2024 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_22
timestamp 1644511149
transform 1 0 3128 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_129
timestamp 1644511149
transform 1 0 12972 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1644511149
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_148
timestamp 1644511149
transform 1 0 14720 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_159
timestamp 1644511149
transform 1 0 15732 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_168
timestamp 1644511149
transform 1 0 16560 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_176
timestamp 1644511149
transform 1 0 17296 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_180
timestamp 1644511149
transform 1 0 17664 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_190
timestamp 1644511149
transform 1 0 18584 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_205
timestamp 1644511149
transform 1 0 19964 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_211
timestamp 1644511149
transform 1 0 20516 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_216
timestamp 1644511149
transform 1 0 20976 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_226
timestamp 1644511149
transform 1 0 21896 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_238
timestamp 1644511149
transform 1 0 23000 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1644511149
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_257
timestamp 1644511149
transform 1 0 24748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_265
timestamp 1644511149
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_277
timestamp 1644511149
transform 1 0 26588 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_285
timestamp 1644511149
transform 1 0 27324 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_302
timestamp 1644511149
transform 1 0 28888 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_325
timestamp 1644511149
transform 1 0 31004 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_337
timestamp 1644511149
transform 1 0 32108 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_355
timestamp 1644511149
transform 1 0 33764 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1644511149
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_371
timestamp 1644511149
transform 1 0 35236 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_385
timestamp 1644511149
transform 1 0 36524 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_391
timestamp 1644511149
transform 1 0 37076 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_395
timestamp 1644511149
transform 1 0 37444 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_407
timestamp 1644511149
transform 1 0 38548 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1644511149
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_421
timestamp 1644511149
transform 1 0 39836 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_425
timestamp 1644511149
transform 1 0 40204 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_447
timestamp 1644511149
transform 1 0 42228 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_6
timestamp 1644511149
transform 1 0 1656 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_13
timestamp 1644511149
transform 1 0 2300 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_25
timestamp 1644511149
transform 1 0 3404 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_37
timestamp 1644511149
transform 1 0 4508 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_49
timestamp 1644511149
transform 1 0 5612 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_130
timestamp 1644511149
transform 1 0 13064 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_144
timestamp 1644511149
transform 1 0 14352 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_153
timestamp 1644511149
transform 1 0 15180 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_160
timestamp 1644511149
transform 1 0 15824 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_181
timestamp 1644511149
transform 1 0 17756 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_189
timestamp 1644511149
transform 1 0 18492 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_197
timestamp 1644511149
transform 1 0 19228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_214
timestamp 1644511149
transform 1 0 20792 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1644511149
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_243
timestamp 1644511149
transform 1 0 23460 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_251
timestamp 1644511149
transform 1 0 24196 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_258
timestamp 1644511149
transform 1 0 24840 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_268
timestamp 1644511149
transform 1 0 25760 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_272
timestamp 1644511149
transform 1 0 26128 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_276
timestamp 1644511149
transform 1 0 26496 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_297
timestamp 1644511149
transform 1 0 28428 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_305
timestamp 1644511149
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_317
timestamp 1644511149
transform 1 0 30268 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_327
timestamp 1644511149
transform 1 0 31188 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1644511149
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_345
timestamp 1644511149
transform 1 0 32844 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_356
timestamp 1644511149
transform 1 0 33856 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_367
timestamp 1644511149
transform 1 0 34868 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_378
timestamp 1644511149
transform 1 0 35880 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_390
timestamp 1644511149
transform 1 0 36984 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_414
timestamp 1644511149
transform 1 0 39192 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_422
timestamp 1644511149
transform 1 0 39928 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_426
timestamp 1644511149
transform 1 0 40296 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_433
timestamp 1644511149
transform 1 0 40940 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_440
timestamp 1644511149
transform 1 0 41584 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_449
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1644511149
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_121
timestamp 1644511149
transform 1 0 12236 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_125
timestamp 1644511149
transform 1 0 12604 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1644511149
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_146
timestamp 1644511149
transform 1 0 14536 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_157
timestamp 1644511149
transform 1 0 15548 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_167
timestamp 1644511149
transform 1 0 16468 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_176
timestamp 1644511149
transform 1 0 17296 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_184
timestamp 1644511149
transform 1 0 18032 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_200
timestamp 1644511149
transform 1 0 19504 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_210
timestamp 1644511149
transform 1 0 20424 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_221
timestamp 1644511149
transform 1 0 21436 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_230
timestamp 1644511149
transform 1 0 22264 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_242
timestamp 1644511149
transform 1 0 23368 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1644511149
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_260
timestamp 1644511149
transform 1 0 25024 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_271
timestamp 1644511149
transform 1 0 26036 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_280
timestamp 1644511149
transform 1 0 26864 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_288
timestamp 1644511149
transform 1 0 27600 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_296
timestamp 1644511149
transform 1 0 28336 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_321
timestamp 1644511149
transform 1 0 30636 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_328
timestamp 1644511149
transform 1 0 31280 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_336
timestamp 1644511149
transform 1 0 32016 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_347
timestamp 1644511149
transform 1 0 33028 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_359
timestamp 1644511149
transform 1 0 34132 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_371
timestamp 1644511149
transform 1 0 35236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_383
timestamp 1644511149
transform 1 0 36340 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_398
timestamp 1644511149
transform 1 0 37720 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_410
timestamp 1644511149
transform 1 0 38824 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_418
timestamp 1644511149
transform 1 0 39560 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_421
timestamp 1644511149
transform 1 0 39836 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_425
timestamp 1644511149
transform 1 0 40204 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_447
timestamp 1644511149
transform 1 0 42228 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_30
timestamp 1644511149
transform 1 0 3864 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_42
timestamp 1644511149
transform 1 0 4968 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1644511149
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_129
timestamp 1644511149
transform 1 0 12972 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_141
timestamp 1644511149
transform 1 0 14076 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_148
timestamp 1644511149
transform 1 0 14720 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_152
timestamp 1644511149
transform 1 0 15088 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_159
timestamp 1644511149
transform 1 0 15732 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1644511149
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_176
timestamp 1644511149
transform 1 0 17296 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_189
timestamp 1644511149
transform 1 0 18492 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_196
timestamp 1644511149
transform 1 0 19136 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_202
timestamp 1644511149
transform 1 0 19688 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_213
timestamp 1644511149
transform 1 0 20700 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_221
timestamp 1644511149
transform 1 0 21436 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_228
timestamp 1644511149
transform 1 0 22080 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_248
timestamp 1644511149
transform 1 0 23920 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_260
timestamp 1644511149
transform 1 0 25024 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_276
timestamp 1644511149
transform 1 0 26496 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_293
timestamp 1644511149
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_305
timestamp 1644511149
transform 1 0 29164 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_323
timestamp 1644511149
transform 1 0 30820 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1644511149
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_361
timestamp 1644511149
transform 1 0 34316 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_369
timestamp 1644511149
transform 1 0 35052 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_381
timestamp 1644511149
transform 1 0 36156 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_389
timestamp 1644511149
transform 1 0 36892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_402
timestamp 1644511149
transform 1 0 38088 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_414
timestamp 1644511149
transform 1 0 39192 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_426
timestamp 1644511149
transform 1 0 40296 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_438
timestamp 1644511149
transform 1 0 41400 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_443
timestamp 1644511149
transform 1 0 41860 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1644511149
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_449
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_9
timestamp 1644511149
transform 1 0 1932 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_13
timestamp 1644511149
transform 1 0 2300 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_17
timestamp 1644511149
transform 1 0 2668 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_21
timestamp 1644511149
transform 1 0 3036 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_105
timestamp 1644511149
transform 1 0 10764 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_115
timestamp 1644511149
transform 1 0 11684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_127
timestamp 1644511149
transform 1 0 12788 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_131
timestamp 1644511149
transform 1 0 13156 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_136
timestamp 1644511149
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_149
timestamp 1644511149
transform 1 0 14812 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_158
timestamp 1644511149
transform 1 0 15640 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_166
timestamp 1644511149
transform 1 0 16376 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_172
timestamp 1644511149
transform 1 0 16928 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_178
timestamp 1644511149
transform 1 0 17480 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_186
timestamp 1644511149
transform 1 0 18216 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1644511149
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_203
timestamp 1644511149
transform 1 0 19780 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_207
timestamp 1644511149
transform 1 0 20148 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_225
timestamp 1644511149
transform 1 0 21804 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_231
timestamp 1644511149
transform 1 0 22356 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_248
timestamp 1644511149
transform 1 0 23920 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_265
timestamp 1644511149
transform 1 0 25484 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_284
timestamp 1644511149
transform 1 0 27232 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_304
timestamp 1644511149
transform 1 0 29072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_317
timestamp 1644511149
transform 1 0 30268 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_324
timestamp 1644511149
transform 1 0 30912 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_344
timestamp 1644511149
transform 1 0 32752 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_356
timestamp 1644511149
transform 1 0 33856 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_369
timestamp 1644511149
transform 1 0 35052 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_381
timestamp 1644511149
transform 1 0 36156 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_399
timestamp 1644511149
transform 1 0 37812 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_405
timestamp 1644511149
transform 1 0 38364 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_416
timestamp 1644511149
transform 1 0 39376 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_421
timestamp 1644511149
transform 1 0 39836 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_429
timestamp 1644511149
transform 1 0 40572 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_433
timestamp 1644511149
transform 1 0 40940 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_440
timestamp 1644511149
transform 1 0 41584 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_447
timestamp 1644511149
transform 1 0 42228 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1644511149
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1644511149
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1644511149
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1644511149
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_129
timestamp 1644511149
transform 1 0 12972 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_135
timestamp 1644511149
transform 1 0 13524 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_146
timestamp 1644511149
transform 1 0 14536 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_156
timestamp 1644511149
transform 1 0 15456 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_164
timestamp 1644511149
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_174
timestamp 1644511149
transform 1 0 17112 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_181
timestamp 1644511149
transform 1 0 17756 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_189
timestamp 1644511149
transform 1 0 18492 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_200
timestamp 1644511149
transform 1 0 19504 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_204
timestamp 1644511149
transform 1 0 19872 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1644511149
transform 1 0 20240 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1644511149
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_231
timestamp 1644511149
transform 1 0 22356 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_243
timestamp 1644511149
transform 1 0 23460 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_255
timestamp 1644511149
transform 1 0 24564 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_267
timestamp 1644511149
transform 1 0 25668 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1644511149
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_293
timestamp 1644511149
transform 1 0 28060 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_297
timestamp 1644511149
transform 1 0 28428 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_301
timestamp 1644511149
transform 1 0 28796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_312
timestamp 1644511149
transform 1 0 29808 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_318
timestamp 1644511149
transform 1 0 30360 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_326
timestamp 1644511149
transform 1 0 31096 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_334
timestamp 1644511149
transform 1 0 31832 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_341
timestamp 1644511149
transform 1 0 32476 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_349
timestamp 1644511149
transform 1 0 33212 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_367
timestamp 1644511149
transform 1 0 34868 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_379
timestamp 1644511149
transform 1 0 35972 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1644511149
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_393
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_412
timestamp 1644511149
transform 1 0 39008 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_419
timestamp 1644511149
transform 1 0 39652 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_444
timestamp 1644511149
transform 1 0 41952 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_449
timestamp 1644511149
transform 1 0 42412 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1644511149
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1644511149
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_105
timestamp 1644511149
transform 1 0 10764 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_116
timestamp 1644511149
transform 1 0 11776 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_128
timestamp 1644511149
transform 1 0 12880 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_136
timestamp 1644511149
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_145
timestamp 1644511149
transform 1 0 14444 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_151
timestamp 1644511149
transform 1 0 14996 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_165
timestamp 1644511149
transform 1 0 16284 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_173
timestamp 1644511149
transform 1 0 17020 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_184
timestamp 1644511149
transform 1 0 18032 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_203
timestamp 1644511149
transform 1 0 19780 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_211
timestamp 1644511149
transform 1 0 20516 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_231
timestamp 1644511149
transform 1 0 22356 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_238
timestamp 1644511149
transform 1 0 23000 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1644511149
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_269
timestamp 1644511149
transform 1 0 25852 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_281
timestamp 1644511149
transform 1 0 26956 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_293
timestamp 1644511149
transform 1 0 28060 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_304
timestamp 1644511149
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_317
timestamp 1644511149
transform 1 0 30268 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_324
timestamp 1644511149
transform 1 0 30912 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_336
timestamp 1644511149
transform 1 0 32016 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_354
timestamp 1644511149
transform 1 0 33672 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_362
timestamp 1644511149
transform 1 0 34408 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_377
timestamp 1644511149
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_389
timestamp 1644511149
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_401
timestamp 1644511149
transform 1 0 37996 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_409
timestamp 1644511149
transform 1 0 38732 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_415
timestamp 1644511149
transform 1 0 39284 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1644511149
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_421
timestamp 1644511149
transform 1 0 39836 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_446
timestamp 1644511149
transform 1 0 42136 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_450
timestamp 1644511149
transform 1 0 42504 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_12
timestamp 1644511149
transform 1 0 2208 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_24
timestamp 1644511149
transform 1 0 3312 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_36
timestamp 1644511149
transform 1 0 4416 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_48
timestamp 1644511149
transform 1 0 5520 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_101
timestamp 1644511149
transform 1 0 10396 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp 1644511149
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_122
timestamp 1644511149
transform 1 0 12328 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_144
timestamp 1644511149
transform 1 0 14352 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1644511149
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_174
timestamp 1644511149
transform 1 0 17112 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_180
timestamp 1644511149
transform 1 0 17664 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_197
timestamp 1644511149
transform 1 0 19228 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_204
timestamp 1644511149
transform 1 0 19872 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_216
timestamp 1644511149
transform 1 0 20976 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_247
timestamp 1644511149
transform 1 0 23828 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_256
timestamp 1644511149
transform 1 0 24656 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_264
timestamp 1644511149
transform 1 0 25392 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_271
timestamp 1644511149
transform 1 0 26036 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1644511149
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_284
timestamp 1644511149
transform 1 0 27232 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_296
timestamp 1644511149
transform 1 0 28336 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_306
timestamp 1644511149
transform 1 0 29256 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_316
timestamp 1644511149
transform 1 0 30176 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_328
timestamp 1644511149
transform 1 0 31280 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_343
timestamp 1644511149
transform 1 0 32660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_355
timestamp 1644511149
transform 1 0 33764 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_363
timestamp 1644511149
transform 1 0 34500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_372
timestamp 1644511149
transform 1 0 35328 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_384
timestamp 1644511149
transform 1 0 36432 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_398
timestamp 1644511149
transform 1 0 37720 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_410
timestamp 1644511149
transform 1 0 38824 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_419
timestamp 1644511149
transform 1 0 39652 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_444
timestamp 1644511149
transform 1 0 41952 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_449
timestamp 1644511149
transform 1 0 42412 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_24
timestamp 1644511149
transform 1 0 3312 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_63
timestamp 1644511149
transform 1 0 6900 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_75
timestamp 1644511149
transform 1 0 8004 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_103
timestamp 1644511149
transform 1 0 10580 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_116
timestamp 1644511149
transform 1 0 11776 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_128
timestamp 1644511149
transform 1 0 12880 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_153
timestamp 1644511149
transform 1 0 15180 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_169
timestamp 1644511149
transform 1 0 16652 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_181
timestamp 1644511149
transform 1 0 17756 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_187
timestamp 1644511149
transform 1 0 18308 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1644511149
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_214
timestamp 1644511149
transform 1 0 20792 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_222
timestamp 1644511149
transform 1 0 21528 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_227
timestamp 1644511149
transform 1 0 21988 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_247
timestamp 1644511149
transform 1 0 23828 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1644511149
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_261
timestamp 1644511149
transform 1 0 25116 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_275
timestamp 1644511149
transform 1 0 26404 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_286
timestamp 1644511149
transform 1 0 27416 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_294
timestamp 1644511149
transform 1 0 28152 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_306
timestamp 1644511149
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_319
timestamp 1644511149
transform 1 0 30452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_331
timestamp 1644511149
transform 1 0 31556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_343
timestamp 1644511149
transform 1 0 32660 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_355
timestamp 1644511149
transform 1 0 33764 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1644511149
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_372
timestamp 1644511149
transform 1 0 35328 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_384
timestamp 1644511149
transform 1 0 36432 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_392
timestamp 1644511149
transform 1 0 37168 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_402
timestamp 1644511149
transform 1 0 38088 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_409
timestamp 1644511149
transform 1 0 38732 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_416
timestamp 1644511149
transform 1 0 39376 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_421
timestamp 1644511149
transform 1 0 39836 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_425
timestamp 1644511149
transform 1 0 40204 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_447
timestamp 1644511149
transform 1 0 42228 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_9
timestamp 1644511149
transform 1 0 1932 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_21
timestamp 1644511149
transform 1 0 3036 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_33
timestamp 1644511149
transform 1 0 4140 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_45
timestamp 1644511149
transform 1 0 5244 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_52
timestamp 1644511149
transform 1 0 5888 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_93
timestamp 1644511149
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1644511149
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1644511149
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_125
timestamp 1644511149
transform 1 0 12604 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_144
timestamp 1644511149
transform 1 0 14352 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_148
timestamp 1644511149
transform 1 0 14720 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_154
timestamp 1644511149
transform 1 0 15272 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_163
timestamp 1644511149
transform 1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1644511149
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_174
timestamp 1644511149
transform 1 0 17112 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_186
timestamp 1644511149
transform 1 0 18216 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_194
timestamp 1644511149
transform 1 0 18952 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_200
timestamp 1644511149
transform 1 0 19504 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1644511149
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1644511149
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_237
timestamp 1644511149
transform 1 0 22908 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_245
timestamp 1644511149
transform 1 0 23644 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_253
timestamp 1644511149
transform 1 0 24380 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_263
timestamp 1644511149
transform 1 0 25300 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_271
timestamp 1644511149
transform 1 0 26036 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_276
timestamp 1644511149
transform 1 0 26496 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_288
timestamp 1644511149
transform 1 0 27600 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_301
timestamp 1644511149
transform 1 0 28796 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_318
timestamp 1644511149
transform 1 0 30360 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_325
timestamp 1644511149
transform 1 0 31004 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_332
timestamp 1644511149
transform 1 0 31648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_343
timestamp 1644511149
transform 1 0 32660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_355
timestamp 1644511149
transform 1 0 33764 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_359
timestamp 1644511149
transform 1 0 34132 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_371
timestamp 1644511149
transform 1 0 35236 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_379
timestamp 1644511149
transform 1 0 35972 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_388
timestamp 1644511149
transform 1 0 36800 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_397
timestamp 1644511149
transform 1 0 37628 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_406
timestamp 1644511149
transform 1 0 38456 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_426
timestamp 1644511149
transform 1 0 40296 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_432
timestamp 1644511149
transform 1 0 40848 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_436
timestamp 1644511149
transform 1 0 41216 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_443
timestamp 1644511149
transform 1 0 41860 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1644511149
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_449
timestamp 1644511149
transform 1 0 42412 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_12
timestamp 1644511149
transform 1 0 2208 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_19
timestamp 1644511149
transform 1 0 2852 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_51
timestamp 1644511149
transform 1 0 5796 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_75
timestamp 1644511149
transform 1 0 8004 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_109
timestamp 1644511149
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_121
timestamp 1644511149
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_136
timestamp 1644511149
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_149
timestamp 1644511149
transform 1 0 14812 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_155
timestamp 1644511149
transform 1 0 15364 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_164
timestamp 1644511149
transform 1 0 16192 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_176
timestamp 1644511149
transform 1 0 17296 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_184
timestamp 1644511149
transform 1 0 18032 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_202
timestamp 1644511149
transform 1 0 19688 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_209
timestamp 1644511149
transform 1 0 20332 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_213
timestamp 1644511149
transform 1 0 20700 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_220
timestamp 1644511149
transform 1 0 21344 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_228
timestamp 1644511149
transform 1 0 22080 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_240
timestamp 1644511149
transform 1 0 23184 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_258
timestamp 1644511149
transform 1 0 24840 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_272
timestamp 1644511149
transform 1 0 26128 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_285
timestamp 1644511149
transform 1 0 27324 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_294
timestamp 1644511149
transform 1 0 28152 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_303
timestamp 1644511149
transform 1 0 28980 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1644511149
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_328
timestamp 1644511149
transform 1 0 31280 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_348
timestamp 1644511149
transform 1 0 33120 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_352
timestamp 1644511149
transform 1 0 33488 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_360
timestamp 1644511149
transform 1 0 34224 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_372
timestamp 1644511149
transform 1 0 35328 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_383
timestamp 1644511149
transform 1 0 36340 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_393
timestamp 1644511149
transform 1 0 37260 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_403
timestamp 1644511149
transform 1 0 38180 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_411
timestamp 1644511149
transform 1 0 38916 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_416
timestamp 1644511149
transform 1 0 39376 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_421
timestamp 1644511149
transform 1 0 39836 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_428
timestamp 1644511149
transform 1 0 40480 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_435
timestamp 1644511149
transform 1 0 41124 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_442
timestamp 1644511149
transform 1 0 41768 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_450
timestamp 1644511149
transform 1 0 42504 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_7
timestamp 1644511149
transform 1 0 1748 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_29
timestamp 1644511149
transform 1 0 3772 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_41
timestamp 1644511149
transform 1 0 4876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_53
timestamp 1644511149
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_93
timestamp 1644511149
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1644511149
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1644511149
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_137
timestamp 1644511149
transform 1 0 13708 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_145
timestamp 1644511149
transform 1 0 14444 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_150
timestamp 1644511149
transform 1 0 14904 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_164
timestamp 1644511149
transform 1 0 16192 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_185
timestamp 1644511149
transform 1 0 18124 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_193
timestamp 1644511149
transform 1 0 18860 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_210
timestamp 1644511149
transform 1 0 20424 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1644511149
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_229
timestamp 1644511149
transform 1 0 22172 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_239
timestamp 1644511149
transform 1 0 23092 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_247
timestamp 1644511149
transform 1 0 23828 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_256
timestamp 1644511149
transform 1 0 24656 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_266
timestamp 1644511149
transform 1 0 25576 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1644511149
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1644511149
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_290
timestamp 1644511149
transform 1 0 27784 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_301
timestamp 1644511149
transform 1 0 28796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_312
timestamp 1644511149
transform 1 0 29808 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_324
timestamp 1644511149
transform 1 0 30912 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_342
timestamp 1644511149
transform 1 0 32568 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_354
timestamp 1644511149
transform 1 0 33672 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_366
timestamp 1644511149
transform 1 0 34776 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_377
timestamp 1644511149
transform 1 0 35788 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_384
timestamp 1644511149
transform 1 0 36432 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_402
timestamp 1644511149
transform 1 0 38088 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_409
timestamp 1644511149
transform 1 0 38732 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_415
timestamp 1644511149
transform 1 0 39284 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_419
timestamp 1644511149
transform 1 0 39652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_444
timestamp 1644511149
transform 1 0 41952 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_449
timestamp 1644511149
transform 1 0 42412 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_24
timestamp 1644511149
transform 1 0 3312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_109
timestamp 1644511149
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_121
timestamp 1644511149
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1644511149
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1644511149
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_157
timestamp 1644511149
transform 1 0 15548 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_168
timestamp 1644511149
transform 1 0 16560 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_180
timestamp 1644511149
transform 1 0 17664 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_187
timestamp 1644511149
transform 1 0 18308 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1644511149
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_197
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_205
timestamp 1644511149
transform 1 0 19964 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_211
timestamp 1644511149
transform 1 0 20516 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_216
timestamp 1644511149
transform 1 0 20976 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_236
timestamp 1644511149
transform 1 0 22816 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_248
timestamp 1644511149
transform 1 0 23920 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_256
timestamp 1644511149
transform 1 0 24656 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_264
timestamp 1644511149
transform 1 0 25392 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_271
timestamp 1644511149
transform 1 0 26036 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_277
timestamp 1644511149
transform 1 0 26588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_283
timestamp 1644511149
transform 1 0 27140 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_291
timestamp 1644511149
transform 1 0 27876 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_303
timestamp 1644511149
transform 1 0 28980 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1644511149
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_314
timestamp 1644511149
transform 1 0 29992 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_321
timestamp 1644511149
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_333
timestamp 1644511149
transform 1 0 31740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_338
timestamp 1644511149
transform 1 0 32200 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_360
timestamp 1644511149
transform 1 0 34224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_375
timestamp 1644511149
transform 1 0 35604 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_384
timestamp 1644511149
transform 1 0 36432 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_396
timestamp 1644511149
transform 1 0 37536 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_408
timestamp 1644511149
transform 1 0 38640 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_416
timestamp 1644511149
transform 1 0 39376 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_421
timestamp 1644511149
transform 1 0 39836 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_425
timestamp 1644511149
transform 1 0 40204 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_447
timestamp 1644511149
transform 1 0 42228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_12
timestamp 1644511149
transform 1 0 2208 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_24
timestamp 1644511149
transform 1 0 3312 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_36
timestamp 1644511149
transform 1 0 4416 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_48
timestamp 1644511149
transform 1 0 5520 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_93
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1644511149
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_125
timestamp 1644511149
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_137
timestamp 1644511149
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_149
timestamp 1644511149
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1644511149
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1644511149
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_181
timestamp 1644511149
transform 1 0 17756 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_185
timestamp 1644511149
transform 1 0 18124 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_189
timestamp 1644511149
transform 1 0 18492 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_193
timestamp 1644511149
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_205
timestamp 1644511149
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1644511149
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1644511149
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_238
timestamp 1644511149
transform 1 0 23000 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_242
timestamp 1644511149
transform 1 0 23368 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_250
timestamp 1644511149
transform 1 0 24104 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_262
timestamp 1644511149
transform 1 0 25208 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_271
timestamp 1644511149
transform 1 0 26036 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1644511149
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_290
timestamp 1644511149
transform 1 0 27784 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_298
timestamp 1644511149
transform 1 0 28520 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_309
timestamp 1644511149
transform 1 0 29532 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_318
timestamp 1644511149
transform 1 0 30360 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_330
timestamp 1644511149
transform 1 0 31464 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_341
timestamp 1644511149
transform 1 0 32476 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_353
timestamp 1644511149
transform 1 0 33580 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_371
timestamp 1644511149
transform 1 0 35236 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_383
timestamp 1644511149
transform 1 0 36340 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1644511149
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_401
timestamp 1644511149
transform 1 0 37996 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_405
timestamp 1644511149
transform 1 0 38364 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_425
timestamp 1644511149
transform 1 0 40204 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_434
timestamp 1644511149
transform 1 0 41032 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1644511149
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1644511149
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_449
timestamp 1644511149
transform 1 0 42412 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_9
timestamp 1644511149
transform 1 0 1932 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_21
timestamp 1644511149
transform 1 0 3036 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_121
timestamp 1644511149
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1644511149
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1644511149
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_153
timestamp 1644511149
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_165
timestamp 1644511149
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_177
timestamp 1644511149
transform 1 0 17388 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_181
timestamp 1644511149
transform 1 0 17756 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_192
timestamp 1644511149
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_206
timestamp 1644511149
transform 1 0 20056 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_218
timestamp 1644511149
transform 1 0 21160 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_230
timestamp 1644511149
transform 1 0 22264 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_235
timestamp 1644511149
transform 1 0 22724 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_248
timestamp 1644511149
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_263
timestamp 1644511149
transform 1 0 25300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_295
timestamp 1644511149
transform 1 0 28244 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_303
timestamp 1644511149
transform 1 0 28980 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1644511149
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_316
timestamp 1644511149
transform 1 0 30176 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_322
timestamp 1644511149
transform 1 0 30728 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_339
timestamp 1644511149
transform 1 0 32292 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_351
timestamp 1644511149
transform 1 0 33396 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1644511149
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_384
timestamp 1644511149
transform 1 0 36432 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_404
timestamp 1644511149
transform 1 0 38272 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1644511149
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1644511149
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_421
timestamp 1644511149
transform 1 0 39836 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_425
timestamp 1644511149
transform 1 0 40204 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_447
timestamp 1644511149
transform 1 0 42228 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_15
timestamp 1644511149
transform 1 0 2484 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_23
timestamp 1644511149
transform 1 0 3220 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1644511149
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1644511149
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1644511149
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_125
timestamp 1644511149
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_137
timestamp 1644511149
transform 1 0 13708 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_143
timestamp 1644511149
transform 1 0 14260 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_160
timestamp 1644511149
transform 1 0 15824 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_172
timestamp 1644511149
transform 1 0 16928 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_176
timestamp 1644511149
transform 1 0 17296 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_193
timestamp 1644511149
transform 1 0 18860 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_204
timestamp 1644511149
transform 1 0 19872 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_212
timestamp 1644511149
transform 1 0 20608 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_220
timestamp 1644511149
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_234
timestamp 1644511149
transform 1 0 22632 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_238
timestamp 1644511149
transform 1 0 23000 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_255
timestamp 1644511149
transform 1 0 24564 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_267
timestamp 1644511149
transform 1 0 25668 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_276
timestamp 1644511149
transform 1 0 26496 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_290
timestamp 1644511149
transform 1 0 27784 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_302
timestamp 1644511149
transform 1 0 28888 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_314
timestamp 1644511149
transform 1 0 29992 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_325
timestamp 1644511149
transform 1 0 31004 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_333
timestamp 1644511149
transform 1 0 31740 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_343
timestamp 1644511149
transform 1 0 32660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_355
timestamp 1644511149
transform 1 0 33764 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_367
timestamp 1644511149
transform 1 0 34868 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_388
timestamp 1644511149
transform 1 0 36800 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_393
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_397
timestamp 1644511149
transform 1 0 37628 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_414
timestamp 1644511149
transform 1 0 39192 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_422
timestamp 1644511149
transform 1 0 39928 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_444
timestamp 1644511149
transform 1 0 41952 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_449
timestamp 1644511149
transform 1 0 42412 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_50
timestamp 1644511149
transform 1 0 5704 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_62
timestamp 1644511149
transform 1 0 6808 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_74
timestamp 1644511149
transform 1 0 7912 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1644511149
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_109
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_121
timestamp 1644511149
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_136
timestamp 1644511149
transform 1 0 13616 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_145
timestamp 1644511149
transform 1 0 14444 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_153
timestamp 1644511149
transform 1 0 15180 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_162
timestamp 1644511149
transform 1 0 16008 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_170
timestamp 1644511149
transform 1 0 16744 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_176
timestamp 1644511149
transform 1 0 17296 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1644511149
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1644511149
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_209
timestamp 1644511149
transform 1 0 20332 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_213
timestamp 1644511149
transform 1 0 20700 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_224
timestamp 1644511149
transform 1 0 21712 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_238
timestamp 1644511149
transform 1 0 23000 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_247
timestamp 1644511149
transform 1 0 23828 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1644511149
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_257
timestamp 1644511149
transform 1 0 24748 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_269
timestamp 1644511149
transform 1 0 25852 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_274
timestamp 1644511149
transform 1 0 26312 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_281
timestamp 1644511149
transform 1 0 26956 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_293
timestamp 1644511149
transform 1 0 28060 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_299
timestamp 1644511149
transform 1 0 28612 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_304
timestamp 1644511149
transform 1 0 29072 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_314
timestamp 1644511149
transform 1 0 29992 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_318
timestamp 1644511149
transform 1 0 30360 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_322
timestamp 1644511149
transform 1 0 30728 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_332
timestamp 1644511149
transform 1 0 31648 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_338
timestamp 1644511149
transform 1 0 32200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_346
timestamp 1644511149
transform 1 0 32936 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_353
timestamp 1644511149
transform 1 0 33580 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_360
timestamp 1644511149
transform 1 0 34224 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_377
timestamp 1644511149
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_389
timestamp 1644511149
transform 1 0 36892 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_399
timestamp 1644511149
transform 1 0 37812 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_411
timestamp 1644511149
transform 1 0 38916 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_416
timestamp 1644511149
transform 1 0 39376 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_421
timestamp 1644511149
transform 1 0 39836 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_444
timestamp 1644511149
transform 1 0 41952 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_450
timestamp 1644511149
transform 1 0 42504 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_93
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1644511149
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_125
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_144
timestamp 1644511149
transform 1 0 14352 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_151
timestamp 1644511149
transform 1 0 14996 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_163
timestamp 1644511149
transform 1 0 16100 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1644511149
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_179
timestamp 1644511149
transform 1 0 17572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_191
timestamp 1644511149
transform 1 0 18676 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_199
timestamp 1644511149
transform 1 0 19412 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_216
timestamp 1644511149
transform 1 0 20976 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_234
timestamp 1644511149
transform 1 0 22632 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_241
timestamp 1644511149
transform 1 0 23276 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_253
timestamp 1644511149
transform 1 0 24380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_270
timestamp 1644511149
transform 1 0 25944 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_278
timestamp 1644511149
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_288
timestamp 1644511149
transform 1 0 27600 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_296
timestamp 1644511149
transform 1 0 28336 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_302
timestamp 1644511149
transform 1 0 28888 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_306
timestamp 1644511149
transform 1 0 29256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_310
timestamp 1644511149
transform 1 0 29624 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_322
timestamp 1644511149
transform 1 0 30728 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_326
timestamp 1644511149
transform 1 0 31096 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_332
timestamp 1644511149
transform 1 0 31648 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_347
timestamp 1644511149
transform 1 0 33028 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_367
timestamp 1644511149
transform 1 0 34868 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_387
timestamp 1644511149
transform 1 0 36708 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1644511149
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_405
timestamp 1644511149
transform 1 0 38364 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_413
timestamp 1644511149
transform 1 0 39100 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_418
timestamp 1644511149
transform 1 0 39560 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_422
timestamp 1644511149
transform 1 0 39928 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_444
timestamp 1644511149
transform 1 0 41952 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_449
timestamp 1644511149
transform 1 0 42412 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1644511149
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_97
timestamp 1644511149
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_109
timestamp 1644511149
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_121
timestamp 1644511149
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1644511149
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1644511149
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_145
timestamp 1644511149
transform 1 0 14444 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_149
timestamp 1644511149
transform 1 0 14812 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_158
timestamp 1644511149
transform 1 0 15640 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_174
timestamp 1644511149
transform 1 0 17112 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_178
timestamp 1644511149
transform 1 0 17480 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1644511149
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1644511149
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_205
timestamp 1644511149
transform 1 0 19964 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_210
timestamp 1644511149
transform 1 0 20424 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_222
timestamp 1644511149
transform 1 0 21528 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_234
timestamp 1644511149
transform 1 0 22632 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_246
timestamp 1644511149
transform 1 0 23736 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_261
timestamp 1644511149
transform 1 0 25116 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_270
timestamp 1644511149
transform 1 0 25944 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_276
timestamp 1644511149
transform 1 0 26496 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_287
timestamp 1644511149
transform 1 0 27508 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_295
timestamp 1644511149
transform 1 0 28244 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_303
timestamp 1644511149
transform 1 0 28980 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1644511149
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_42_321
timestamp 1644511149
transform 1 0 30636 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_327
timestamp 1644511149
transform 1 0 31188 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_334
timestamp 1644511149
transform 1 0 31832 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_346
timestamp 1644511149
transform 1 0 32936 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_353
timestamp 1644511149
transform 1 0 33580 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_361
timestamp 1644511149
transform 1 0 34316 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_377
timestamp 1644511149
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_389
timestamp 1644511149
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_401
timestamp 1644511149
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1644511149
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1644511149
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_421
timestamp 1644511149
transform 1 0 39836 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_427
timestamp 1644511149
transform 1 0 40388 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_431
timestamp 1644511149
transform 1 0 40756 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_438
timestamp 1644511149
transform 1 0 41400 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_445
timestamp 1644511149
transform 1 0 42044 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_125
timestamp 1644511149
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_137
timestamp 1644511149
transform 1 0 13708 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_143
timestamp 1644511149
transform 1 0 14260 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_150
timestamp 1644511149
transform 1 0 14904 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_154
timestamp 1644511149
transform 1 0 15272 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1644511149
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1644511149
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_175
timestamp 1644511149
transform 1 0 17204 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_192
timestamp 1644511149
transform 1 0 18768 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_204
timestamp 1644511149
transform 1 0 19872 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_212
timestamp 1644511149
transform 1 0 20608 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_219
timestamp 1644511149
transform 1 0 21252 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1644511149
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_237
timestamp 1644511149
transform 1 0 22908 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_241
timestamp 1644511149
transform 1 0 23276 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_261
timestamp 1644511149
transform 1 0 25116 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_271
timestamp 1644511149
transform 1 0 26036 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1644511149
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_286
timestamp 1644511149
transform 1 0 27416 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_304
timestamp 1644511149
transform 1 0 29072 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_326
timestamp 1644511149
transform 1 0 31096 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_334
timestamp 1644511149
transform 1 0 31832 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_342
timestamp 1644511149
transform 1 0 32568 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_354
timestamp 1644511149
transform 1 0 33672 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_359
timestamp 1644511149
transform 1 0 34132 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_371
timestamp 1644511149
transform 1 0 35236 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_383
timestamp 1644511149
transform 1 0 36340 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1644511149
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_405
timestamp 1644511149
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_417
timestamp 1644511149
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_429
timestamp 1644511149
transform 1 0 40572 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_437
timestamp 1644511149
transform 1 0 41308 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_443
timestamp 1644511149
transform 1 0 41860 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1644511149
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_449
timestamp 1644511149
transform 1 0 42412 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_117
timestamp 1644511149
transform 1 0 11868 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_136
timestamp 1644511149
transform 1 0 13616 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_149
timestamp 1644511149
transform 1 0 14812 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_159
timestamp 1644511149
transform 1 0 15732 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_169
timestamp 1644511149
transform 1 0 16652 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_176
timestamp 1644511149
transform 1 0 17296 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_188
timestamp 1644511149
transform 1 0 18400 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_206
timestamp 1644511149
transform 1 0 20056 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_210
timestamp 1644511149
transform 1 0 20424 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_214
timestamp 1644511149
transform 1 0 20792 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_226
timestamp 1644511149
transform 1 0 21896 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_232
timestamp 1644511149
transform 1 0 22448 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_243
timestamp 1644511149
transform 1 0 23460 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1644511149
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_256
timestamp 1644511149
transform 1 0 24656 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_267
timestamp 1644511149
transform 1 0 25668 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_287
timestamp 1644511149
transform 1 0 27508 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_295
timestamp 1644511149
transform 1 0 28244 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_304
timestamp 1644511149
transform 1 0 29072 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_316
timestamp 1644511149
transform 1 0 30176 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_332
timestamp 1644511149
transform 1 0 31648 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_341
timestamp 1644511149
transform 1 0 32476 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_353
timestamp 1644511149
transform 1 0 33580 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_360
timestamp 1644511149
transform 1 0 34224 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_368
timestamp 1644511149
transform 1 0 34960 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_380
timestamp 1644511149
transform 1 0 36064 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_392
timestamp 1644511149
transform 1 0 37168 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_404
timestamp 1644511149
transform 1 0 38272 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_416
timestamp 1644511149
transform 1 0 39376 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_421
timestamp 1644511149
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_433
timestamp 1644511149
transform 1 0 40940 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_439
timestamp 1644511149
transform 1 0 41492 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_443
timestamp 1644511149
transform 1 0 41860 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1644511149
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_134
timestamp 1644511149
transform 1 0 13432 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_146
timestamp 1644511149
transform 1 0 14536 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_152
timestamp 1644511149
transform 1 0 15088 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_160
timestamp 1644511149
transform 1 0 15824 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_173
timestamp 1644511149
transform 1 0 17020 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_185
timestamp 1644511149
transform 1 0 18124 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_207
timestamp 1644511149
transform 1 0 20148 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1644511149
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1644511149
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_241
timestamp 1644511149
transform 1 0 23276 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_250
timestamp 1644511149
transform 1 0 24104 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_262
timestamp 1644511149
transform 1 0 25208 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_270
timestamp 1644511149
transform 1 0 25944 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_274
timestamp 1644511149
transform 1 0 26312 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_298
timestamp 1644511149
transform 1 0 28520 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_312
timestamp 1644511149
transform 1 0 29808 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_332
timestamp 1644511149
transform 1 0 31648 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_343
timestamp 1644511149
transform 1 0 32660 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_352
timestamp 1644511149
transform 1 0 33488 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_372
timestamp 1644511149
transform 1 0 35328 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_384
timestamp 1644511149
transform 1 0 36432 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_405
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_417
timestamp 1644511149
transform 1 0 39468 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_444
timestamp 1644511149
transform 1 0 41952 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_449
timestamp 1644511149
transform 1 0 42412 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1644511149
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1644511149
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_148
timestamp 1644511149
transform 1 0 14720 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_156
timestamp 1644511149
transform 1 0 15456 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_164
timestamp 1644511149
transform 1 0 16192 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_172
timestamp 1644511149
transform 1 0 16928 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_184
timestamp 1644511149
transform 1 0 18032 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_192
timestamp 1644511149
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_212
timestamp 1644511149
transform 1 0 20608 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_222
timestamp 1644511149
transform 1 0 21528 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_230
timestamp 1644511149
transform 1 0 22264 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_238
timestamp 1644511149
transform 1 0 23000 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_248
timestamp 1644511149
transform 1 0 23920 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_256
timestamp 1644511149
transform 1 0 24656 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_268
timestamp 1644511149
transform 1 0 25760 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_272
timestamp 1644511149
transform 1 0 26128 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_276
timestamp 1644511149
transform 1 0 26496 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_280
timestamp 1644511149
transform 1 0 26864 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_295
timestamp 1644511149
transform 1 0 28244 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_304
timestamp 1644511149
transform 1 0 29072 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_315
timestamp 1644511149
transform 1 0 30084 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_321
timestamp 1644511149
transform 1 0 30636 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_332
timestamp 1644511149
transform 1 0 31648 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_336
timestamp 1644511149
transform 1 0 32016 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_340
timestamp 1644511149
transform 1 0 32384 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_360
timestamp 1644511149
transform 1 0 34224 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_377
timestamp 1644511149
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_389
timestamp 1644511149
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_401
timestamp 1644511149
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1644511149
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1644511149
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_421
timestamp 1644511149
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_433
timestamp 1644511149
transform 1 0 40940 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_437
timestamp 1644511149
transform 1 0 41308 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_441
timestamp 1644511149
transform 1 0 41676 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_449
timestamp 1644511149
transform 1 0 42412 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_9
timestamp 1644511149
transform 1 0 1932 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_13
timestamp 1644511149
transform 1 0 2300 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_25
timestamp 1644511149
transform 1 0 3404 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_37
timestamp 1644511149
transform 1 0 4508 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_49
timestamp 1644511149
transform 1 0 5612 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1644511149
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_121
timestamp 1644511149
transform 1 0 12236 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_127
timestamp 1644511149
transform 1 0 12788 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_139
timestamp 1644511149
transform 1 0 13892 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_47_150
timestamp 1644511149
transform 1 0 14904 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_156
timestamp 1644511149
transform 1 0 15456 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_164
timestamp 1644511149
transform 1 0 16192 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_177
timestamp 1644511149
transform 1 0 17388 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_188
timestamp 1644511149
transform 1 0 18400 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_196
timestamp 1644511149
transform 1 0 19136 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_204
timestamp 1644511149
transform 1 0 19872 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_211
timestamp 1644511149
transform 1 0 20516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1644511149
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_233
timestamp 1644511149
transform 1 0 22540 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_239
timestamp 1644511149
transform 1 0 23092 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_47_263
timestamp 1644511149
transform 1 0 25300 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_269
timestamp 1644511149
transform 1 0 25852 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_275
timestamp 1644511149
transform 1 0 26404 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1644511149
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_300
timestamp 1644511149
transform 1 0 28704 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_312
timestamp 1644511149
transform 1 0 29808 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_320
timestamp 1644511149
transform 1 0 30544 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_332
timestamp 1644511149
transform 1 0 31648 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_341
timestamp 1644511149
transform 1 0 32476 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_347
timestamp 1644511149
transform 1 0 33028 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_356
timestamp 1644511149
transform 1 0 33856 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_364
timestamp 1644511149
transform 1 0 34592 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_369
timestamp 1644511149
transform 1 0 35052 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_381
timestamp 1644511149
transform 1 0 36156 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_389
timestamp 1644511149
transform 1 0 36892 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_405
timestamp 1644511149
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_417
timestamp 1644511149
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_429
timestamp 1644511149
transform 1 0 40572 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_47_440
timestamp 1644511149
transform 1 0 41584 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_449
timestamp 1644511149
transform 1 0 42412 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_24
timestamp 1644511149
transform 1 0 3312 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_109
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_121
timestamp 1644511149
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_136
timestamp 1644511149
transform 1 0 13616 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_148
timestamp 1644511149
transform 1 0 14720 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_160
timestamp 1644511149
transform 1 0 15824 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_171
timestamp 1644511149
transform 1 0 16836 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_178
timestamp 1644511149
transform 1 0 17480 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_190
timestamp 1644511149
transform 1 0 18584 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_217
timestamp 1644511149
transform 1 0 21068 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_221
timestamp 1644511149
transform 1 0 21436 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_226
timestamp 1644511149
transform 1 0 21896 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_237
timestamp 1644511149
transform 1 0 22908 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1644511149
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1644511149
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_257
timestamp 1644511149
transform 1 0 24748 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_265
timestamp 1644511149
transform 1 0 25484 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_285
timestamp 1644511149
transform 1 0 27324 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_289
timestamp 1644511149
transform 1 0 27692 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_294
timestamp 1644511149
transform 1 0 28152 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_304
timestamp 1644511149
transform 1 0 29072 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_312
timestamp 1644511149
transform 1 0 29808 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_336
timestamp 1644511149
transform 1 0 32016 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_348
timestamp 1644511149
transform 1 0 33120 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_360
timestamp 1644511149
transform 1 0 34224 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_365
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_377
timestamp 1644511149
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_389
timestamp 1644511149
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_401
timestamp 1644511149
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1644511149
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1644511149
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_421
timestamp 1644511149
transform 1 0 39836 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_425
timestamp 1644511149
transform 1 0 40204 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_447
timestamp 1644511149
transform 1 0 42228 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_9
timestamp 1644511149
transform 1 0 1932 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_21
timestamp 1644511149
transform 1 0 3036 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_33
timestamp 1644511149
transform 1 0 4140 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_45
timestamp 1644511149
transform 1 0 5244 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_53
timestamp 1644511149
transform 1 0 5980 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_135
timestamp 1644511149
transform 1 0 13524 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_139
timestamp 1644511149
transform 1 0 13892 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_150
timestamp 1644511149
transform 1 0 14904 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_158
timestamp 1644511149
transform 1 0 15640 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_164
timestamp 1644511149
transform 1 0 16192 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_180
timestamp 1644511149
transform 1 0 17664 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_192
timestamp 1644511149
transform 1 0 18768 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_198
timestamp 1644511149
transform 1 0 19320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_203
timestamp 1644511149
transform 1 0 19780 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_211
timestamp 1644511149
transform 1 0 20516 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1644511149
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1644511149
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_225
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_231
timestamp 1644511149
transform 1 0 22356 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_239
timestamp 1644511149
transform 1 0 23092 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_246
timestamp 1644511149
transform 1 0 23736 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_255
timestamp 1644511149
transform 1 0 24564 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_267
timestamp 1644511149
transform 1 0 25668 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_274
timestamp 1644511149
transform 1 0 26312 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_49_284
timestamp 1644511149
transform 1 0 27232 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_292
timestamp 1644511149
transform 1 0 27968 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_301
timestamp 1644511149
transform 1 0 28796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_313
timestamp 1644511149
transform 1 0 29900 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_321
timestamp 1644511149
transform 1 0 30636 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_332
timestamp 1644511149
transform 1 0 31648 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_349
timestamp 1644511149
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_361
timestamp 1644511149
transform 1 0 34316 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_366
timestamp 1644511149
transform 1 0 34776 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_378
timestamp 1644511149
transform 1 0 35880 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_390
timestamp 1644511149
transform 1 0 36984 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_402
timestamp 1644511149
transform 1 0 38088 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_414
timestamp 1644511149
transform 1 0 39192 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_426
timestamp 1644511149
transform 1 0 40296 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_438
timestamp 1644511149
transform 1 0 41400 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_443
timestamp 1644511149
transform 1 0 41860 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1644511149
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_449
timestamp 1644511149
transform 1 0 42412 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1644511149
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_131
timestamp 1644511149
transform 1 0 13156 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_149
timestamp 1644511149
transform 1 0 14812 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_163
timestamp 1644511149
transform 1 0 16100 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_170
timestamp 1644511149
transform 1 0 16744 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_190
timestamp 1644511149
transform 1 0 18584 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_205
timestamp 1644511149
transform 1 0 19964 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_209
timestamp 1644511149
transform 1 0 20332 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_226
timestamp 1644511149
transform 1 0 21896 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_232
timestamp 1644511149
transform 1 0 22448 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_239
timestamp 1644511149
transform 1 0 23092 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_247
timestamp 1644511149
transform 1 0 23828 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1644511149
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_263
timestamp 1644511149
transform 1 0 25300 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_272
timestamp 1644511149
transform 1 0 26128 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_284
timestamp 1644511149
transform 1 0 27232 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_292
timestamp 1644511149
transform 1 0 27968 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_304
timestamp 1644511149
transform 1 0 29072 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_314
timestamp 1644511149
transform 1 0 29992 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_334
timestamp 1644511149
transform 1 0 31832 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_50_358
timestamp 1644511149
transform 1 0 34040 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_381
timestamp 1644511149
transform 1 0 36156 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_393
timestamp 1644511149
transform 1 0 37260 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_403
timestamp 1644511149
transform 1 0 38180 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_407
timestamp 1644511149
transform 1 0 38548 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_414
timestamp 1644511149
transform 1 0 39192 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_427
timestamp 1644511149
transform 1 0 40388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_439
timestamp 1644511149
transform 1 0 41492 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_447
timestamp 1644511149
transform 1 0 42228 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1644511149
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1644511149
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_129
timestamp 1644511149
transform 1 0 12972 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_134
timestamp 1644511149
transform 1 0 13432 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_147
timestamp 1644511149
transform 1 0 14628 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_154
timestamp 1644511149
transform 1 0 15272 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1644511149
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_177
timestamp 1644511149
transform 1 0 17388 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_181
timestamp 1644511149
transform 1 0 17756 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_185
timestamp 1644511149
transform 1 0 18124 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_205
timestamp 1644511149
transform 1 0 19964 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_51_216
timestamp 1644511149
transform 1 0 20976 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_233
timestamp 1644511149
transform 1 0 22540 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_51_257
timestamp 1644511149
transform 1 0 24748 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_51_271
timestamp 1644511149
transform 1 0 26036 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1644511149
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_284
timestamp 1644511149
transform 1 0 27232 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_293
timestamp 1644511149
transform 1 0 28060 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_313
timestamp 1644511149
transform 1 0 29900 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_325
timestamp 1644511149
transform 1 0 31004 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_333
timestamp 1644511149
transform 1 0 31740 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_346
timestamp 1644511149
transform 1 0 32936 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_356
timestamp 1644511149
transform 1 0 33856 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_367
timestamp 1644511149
transform 1 0 34868 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_371
timestamp 1644511149
transform 1 0 35236 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_388
timestamp 1644511149
transform 1 0 36800 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_412
timestamp 1644511149
transform 1 0 39008 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_432
timestamp 1644511149
transform 1 0 40848 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_443
timestamp 1644511149
transform 1 0 41860 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1644511149
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_449
timestamp 1644511149
transform 1 0 42412 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_146
timestamp 1644511149
transform 1 0 14536 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_153
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_157
timestamp 1644511149
transform 1 0 15548 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_163
timestamp 1644511149
transform 1 0 16100 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_175
timestamp 1644511149
transform 1 0 17204 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_182
timestamp 1644511149
transform 1 0 17848 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1644511149
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_197
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_209
timestamp 1644511149
transform 1 0 20332 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_216
timestamp 1644511149
transform 1 0 20976 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_226
timestamp 1644511149
transform 1 0 21896 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_236
timestamp 1644511149
transform 1 0 22816 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_243
timestamp 1644511149
transform 1 0 23460 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1644511149
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_261
timestamp 1644511149
transform 1 0 25116 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_267
timestamp 1644511149
transform 1 0 25668 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_284
timestamp 1644511149
transform 1 0 27232 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_291
timestamp 1644511149
transform 1 0 27876 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_297
timestamp 1644511149
transform 1 0 28428 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_302
timestamp 1644511149
transform 1 0 28888 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_321
timestamp 1644511149
transform 1 0 30636 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_338
timestamp 1644511149
transform 1 0 32200 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_346
timestamp 1644511149
transform 1 0 32936 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_358
timestamp 1644511149
transform 1 0 34040 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_370
timestamp 1644511149
transform 1 0 35144 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_378
timestamp 1644511149
transform 1 0 35880 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_385
timestamp 1644511149
transform 1 0 36524 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_393
timestamp 1644511149
transform 1 0 37260 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_401
timestamp 1644511149
transform 1 0 37996 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_410
timestamp 1644511149
transform 1 0 38824 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_418
timestamp 1644511149
transform 1 0 39560 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_421
timestamp 1644511149
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_433
timestamp 1644511149
transform 1 0 40940 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_437
timestamp 1644511149
transform 1 0 41308 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_441
timestamp 1644511149
transform 1 0 41676 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_449
timestamp 1644511149
transform 1 0 42412 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1644511149
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1644511149
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_39
timestamp 1644511149
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1644511149
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1644511149
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_53_151
timestamp 1644511149
transform 1 0 14996 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_53_162
timestamp 1644511149
transform 1 0 16008 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_179
timestamp 1644511149
transform 1 0 17572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_191
timestamp 1644511149
transform 1 0 18676 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_203
timestamp 1644511149
transform 1 0 19780 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_211
timestamp 1644511149
transform 1 0 20516 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_220
timestamp 1644511149
transform 1 0 21344 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_228
timestamp 1644511149
transform 1 0 22080 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_240
timestamp 1644511149
transform 1 0 23184 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_245
timestamp 1644511149
transform 1 0 23644 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_251
timestamp 1644511149
transform 1 0 24196 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_256
timestamp 1644511149
transform 1 0 24656 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_274
timestamp 1644511149
transform 1 0 26312 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_53_288
timestamp 1644511149
transform 1 0 27600 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_296
timestamp 1644511149
transform 1 0 28336 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_301
timestamp 1644511149
transform 1 0 28796 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_309
timestamp 1644511149
transform 1 0 29532 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_314
timestamp 1644511149
transform 1 0 29992 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_323
timestamp 1644511149
transform 1 0 30820 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_331
timestamp 1644511149
transform 1 0 31556 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1644511149
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_342
timestamp 1644511149
transform 1 0 32568 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_354
timestamp 1644511149
transform 1 0 33672 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_367
timestamp 1644511149
transform 1 0 34868 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_378
timestamp 1644511149
transform 1 0 35880 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_390
timestamp 1644511149
transform 1 0 36984 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_399
timestamp 1644511149
transform 1 0 37812 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_407
timestamp 1644511149
transform 1 0 38548 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_419
timestamp 1644511149
transform 1 0 39652 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_426
timestamp 1644511149
transform 1 0 40296 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_430
timestamp 1644511149
transform 1 0 40664 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_434
timestamp 1644511149
transform 1 0 41032 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1644511149
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1644511149
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_449
timestamp 1644511149
transform 1 0 42412 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1644511149
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1644511149
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_157
timestamp 1644511149
transform 1 0 15548 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_171
timestamp 1644511149
transform 1 0 16836 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_182
timestamp 1644511149
transform 1 0 17848 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1644511149
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1644511149
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_205
timestamp 1644511149
transform 1 0 19964 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_215
timestamp 1644511149
transform 1 0 20884 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_235
timestamp 1644511149
transform 1 0 22724 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_247
timestamp 1644511149
transform 1 0 23828 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1644511149
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_261
timestamp 1644511149
transform 1 0 25116 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_269
timestamp 1644511149
transform 1 0 25852 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_279
timestamp 1644511149
transform 1 0 26772 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_299
timestamp 1644511149
transform 1 0 28612 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1644511149
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_313
timestamp 1644511149
transform 1 0 29900 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_318
timestamp 1644511149
transform 1 0 30360 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_327
timestamp 1644511149
transform 1 0 31188 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_335
timestamp 1644511149
transform 1 0 31924 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_346
timestamp 1644511149
transform 1 0 32936 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_360
timestamp 1644511149
transform 1 0 34224 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_375
timestamp 1644511149
transform 1 0 35604 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_383
timestamp 1644511149
transform 1 0 36340 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_394
timestamp 1644511149
transform 1 0 37352 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_398
timestamp 1644511149
transform 1 0 37720 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_409
timestamp 1644511149
transform 1 0 38732 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_417
timestamp 1644511149
transform 1 0 39468 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_421
timestamp 1644511149
transform 1 0 39836 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_425
timestamp 1644511149
transform 1 0 40204 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_447
timestamp 1644511149
transform 1 0 42228 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1644511149
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1644511149
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_39
timestamp 1644511149
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1644511149
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1644511149
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1644511149
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1644511149
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_191
timestamp 1644511149
transform 1 0 18676 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_200
timestamp 1644511149
transform 1 0 19504 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_206
timestamp 1644511149
transform 1 0 20056 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_210
timestamp 1644511149
transform 1 0 20424 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_220
timestamp 1644511149
transform 1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_237
timestamp 1644511149
transform 1 0 22908 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_243
timestamp 1644511149
transform 1 0 23460 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_264
timestamp 1644511149
transform 1 0 25392 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_275
timestamp 1644511149
transform 1 0 26404 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1644511149
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_284
timestamp 1644511149
transform 1 0 27232 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_296
timestamp 1644511149
transform 1 0 28336 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_303
timestamp 1644511149
transform 1 0 28980 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_323
timestamp 1644511149
transform 1 0 30820 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_331
timestamp 1644511149
transform 1 0 31556 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1644511149
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_345
timestamp 1644511149
transform 1 0 32844 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_353
timestamp 1644511149
transform 1 0 33580 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_372
timestamp 1644511149
transform 1 0 35328 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_380
timestamp 1644511149
transform 1 0 36064 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_388
timestamp 1644511149
transform 1 0 36800 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_409
timestamp 1644511149
transform 1 0 38732 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_418
timestamp 1644511149
transform 1 0 39560 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_438
timestamp 1644511149
transform 1 0 41400 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_446
timestamp 1644511149
transform 1 0 42136 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_449
timestamp 1644511149
transform 1 0 42412 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1644511149
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_149
timestamp 1644511149
transform 1 0 14812 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_155
timestamp 1644511149
transform 1 0 15364 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_167
timestamp 1644511149
transform 1 0 16468 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_174
timestamp 1644511149
transform 1 0 17112 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_185
timestamp 1644511149
transform 1 0 18124 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_192
timestamp 1644511149
transform 1 0 18768 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_207
timestamp 1644511149
transform 1 0 20148 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_214
timestamp 1644511149
transform 1 0 20792 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_221
timestamp 1644511149
transform 1 0 21436 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_229
timestamp 1644511149
transform 1 0 22172 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_248
timestamp 1644511149
transform 1 0 23920 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_261
timestamp 1644511149
transform 1 0 25116 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_275
timestamp 1644511149
transform 1 0 26404 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_286
timestamp 1644511149
transform 1 0 27416 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_293
timestamp 1644511149
transform 1 0 28060 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_305
timestamp 1644511149
transform 1 0 29164 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_317
timestamp 1644511149
transform 1 0 30268 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_325
timestamp 1644511149
transform 1 0 31004 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_333
timestamp 1644511149
transform 1 0 31740 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_343
timestamp 1644511149
transform 1 0 32660 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_353
timestamp 1644511149
transform 1 0 33580 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_361
timestamp 1644511149
transform 1 0 34316 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_369
timestamp 1644511149
transform 1 0 35052 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_381
timestamp 1644511149
transform 1 0 36156 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_389
timestamp 1644511149
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_410
timestamp 1644511149
transform 1 0 38824 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_418
timestamp 1644511149
transform 1 0 39560 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_421
timestamp 1644511149
transform 1 0 39836 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_425
timestamp 1644511149
transform 1 0 40204 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_447
timestamp 1644511149
transform 1 0 42228 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1644511149
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1644511149
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1644511149
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1644511149
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_149
timestamp 1644511149
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1644511149
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_172
timestamp 1644511149
transform 1 0 16928 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_184
timestamp 1644511149
transform 1 0 18032 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_190
timestamp 1644511149
transform 1 0 18584 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_199
timestamp 1644511149
transform 1 0 19412 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_207
timestamp 1644511149
transform 1 0 20148 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_220
timestamp 1644511149
transform 1 0 21344 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_230
timestamp 1644511149
transform 1 0 22264 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_236
timestamp 1644511149
transform 1 0 22816 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_241
timestamp 1644511149
transform 1 0 23276 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_248
timestamp 1644511149
transform 1 0 23920 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_256
timestamp 1644511149
transform 1 0 24656 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_262
timestamp 1644511149
transform 1 0 25208 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_269
timestamp 1644511149
transform 1 0 25852 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_276
timestamp 1644511149
transform 1 0 26496 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_303
timestamp 1644511149
transform 1 0 28980 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_315
timestamp 1644511149
transform 1 0 30084 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_327
timestamp 1644511149
transform 1 0 31188 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1644511149
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_342
timestamp 1644511149
transform 1 0 32568 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_350
timestamp 1644511149
transform 1 0 33304 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_362
timestamp 1644511149
transform 1 0 34408 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_374
timestamp 1644511149
transform 1 0 35512 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_386
timestamp 1644511149
transform 1 0 36616 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_406
timestamp 1644511149
transform 1 0 38456 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_417
timestamp 1644511149
transform 1 0 39468 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_444
timestamp 1644511149
transform 1 0 41952 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_449
timestamp 1644511149
transform 1 0 42412 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1644511149
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1644511149
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_157
timestamp 1644511149
transform 1 0 15548 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_165
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_173
timestamp 1644511149
transform 1 0 17020 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_192
timestamp 1644511149
transform 1 0 18768 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_205
timestamp 1644511149
transform 1 0 19964 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_209
timestamp 1644511149
transform 1 0 20332 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_229
timestamp 1644511149
transform 1 0 22172 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_241
timestamp 1644511149
transform 1 0 23276 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_249
timestamp 1644511149
transform 1 0 24012 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_265
timestamp 1644511149
transform 1 0 25484 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_273
timestamp 1644511149
transform 1 0 26220 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_277
timestamp 1644511149
transform 1 0 26588 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_286
timestamp 1644511149
transform 1 0 27416 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_293
timestamp 1644511149
transform 1 0 28060 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_305
timestamp 1644511149
transform 1 0 29164 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_318
timestamp 1644511149
transform 1 0 30360 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_330
timestamp 1644511149
transform 1 0 31464 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_334
timestamp 1644511149
transform 1 0 31832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_351
timestamp 1644511149
transform 1 0 33396 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1644511149
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_369
timestamp 1644511149
transform 1 0 35052 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_374
timestamp 1644511149
transform 1 0 35512 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_383
timestamp 1644511149
transform 1 0 36340 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_387
timestamp 1644511149
transform 1 0 36708 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_392
timestamp 1644511149
transform 1 0 37168 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_399
timestamp 1644511149
transform 1 0 37812 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_403
timestamp 1644511149
transform 1 0 38180 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_411
timestamp 1644511149
transform 1 0 38916 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1644511149
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_437
timestamp 1644511149
transform 1 0 41308 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_444
timestamp 1644511149
transform 1 0 41952 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_450
timestamp 1644511149
transform 1 0 42504 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1644511149
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1644511149
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1644511149
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1644511149
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1644511149
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_143
timestamp 1644511149
transform 1 0 14260 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_150
timestamp 1644511149
transform 1 0 14904 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_158
timestamp 1644511149
transform 1 0 15640 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_166
timestamp 1644511149
transform 1 0 16376 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_173
timestamp 1644511149
transform 1 0 17020 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_181
timestamp 1644511149
transform 1 0 17756 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_190
timestamp 1644511149
transform 1 0 18584 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_194
timestamp 1644511149
transform 1 0 18952 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_203
timestamp 1644511149
transform 1 0 19780 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_218
timestamp 1644511149
transform 1 0 21160 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_235
timestamp 1644511149
transform 1 0 22724 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_250
timestamp 1644511149
transform 1 0 24104 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_262
timestamp 1644511149
transform 1 0 25208 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_271
timestamp 1644511149
transform 1 0 26036 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1644511149
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_284
timestamp 1644511149
transform 1 0 27232 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_296
timestamp 1644511149
transform 1 0 28336 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_308
timestamp 1644511149
transform 1 0 29440 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_312
timestamp 1644511149
transform 1 0 29808 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_319
timestamp 1644511149
transform 1 0 30452 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1644511149
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1644511149
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_344
timestamp 1644511149
transform 1 0 32752 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_353
timestamp 1644511149
transform 1 0 33580 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_360
timestamp 1644511149
transform 1 0 34224 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_59_382
timestamp 1644511149
transform 1 0 36248 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_390
timestamp 1644511149
transform 1 0 36984 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_401
timestamp 1644511149
transform 1 0 37996 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_414
timestamp 1644511149
transform 1 0 39192 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_422
timestamp 1644511149
transform 1 0 39928 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_444
timestamp 1644511149
transform 1 0 41952 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_449
timestamp 1644511149
transform 1 0 42412 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1644511149
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_162
timestamp 1644511149
transform 1 0 16008 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_176
timestamp 1644511149
transform 1 0 17296 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_184
timestamp 1644511149
transform 1 0 18032 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_192
timestamp 1644511149
transform 1 0 18768 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_205
timestamp 1644511149
transform 1 0 19964 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_217
timestamp 1644511149
transform 1 0 21068 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_60_241
timestamp 1644511149
transform 1 0 23276 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_249
timestamp 1644511149
transform 1 0 24012 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_260
timestamp 1644511149
transform 1 0 25024 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_264
timestamp 1644511149
transform 1 0 25392 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_273
timestamp 1644511149
transform 1 0 26220 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_285
timestamp 1644511149
transform 1 0 27324 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_297
timestamp 1644511149
transform 1 0 28428 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_305
timestamp 1644511149
transform 1 0 29164 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_325
timestamp 1644511149
transform 1 0 31004 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_333
timestamp 1644511149
transform 1 0 31740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_340
timestamp 1644511149
transform 1 0 32384 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_354
timestamp 1644511149
transform 1 0 33672 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_362
timestamp 1644511149
transform 1 0 34408 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_373
timestamp 1644511149
transform 1 0 35420 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_385
timestamp 1644511149
transform 1 0 36524 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_402
timestamp 1644511149
transform 1 0 38088 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_410
timestamp 1644511149
transform 1 0 38824 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_418
timestamp 1644511149
transform 1 0 39560 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_424
timestamp 1644511149
transform 1 0 40112 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_433
timestamp 1644511149
transform 1 0 40940 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_440
timestamp 1644511149
transform 1 0 41584 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_447
timestamp 1644511149
transform 1 0 42228 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_30
timestamp 1644511149
transform 1 0 3864 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_46
timestamp 1644511149
transform 1 0 5336 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1644511149
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_145
timestamp 1644511149
transform 1 0 14444 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_150
timestamp 1644511149
transform 1 0 14904 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_158
timestamp 1644511149
transform 1 0 15640 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_164
timestamp 1644511149
transform 1 0 16192 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_175
timestamp 1644511149
transform 1 0 17204 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_182
timestamp 1644511149
transform 1 0 17848 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_194
timestamp 1644511149
transform 1 0 18952 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_206
timestamp 1644511149
transform 1 0 20056 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_218
timestamp 1644511149
transform 1 0 21160 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_233
timestamp 1644511149
transform 1 0 22540 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_238
timestamp 1644511149
transform 1 0 23000 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_249
timestamp 1644511149
transform 1 0 24012 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_256
timestamp 1644511149
transform 1 0 24656 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_61_269
timestamp 1644511149
transform 1 0 25852 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_277
timestamp 1644511149
transform 1 0 26588 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_288
timestamp 1644511149
transform 1 0 27600 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_296
timestamp 1644511149
transform 1 0 28336 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_313
timestamp 1644511149
transform 1 0 29900 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_324
timestamp 1644511149
transform 1 0 30912 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_344
timestamp 1644511149
transform 1 0 32752 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_350
timestamp 1644511149
transform 1 0 33304 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_367
timestamp 1644511149
transform 1 0 34868 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_378
timestamp 1644511149
transform 1 0 35880 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_390
timestamp 1644511149
transform 1 0 36984 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_417
timestamp 1644511149
transform 1 0 39468 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_437
timestamp 1644511149
transform 1 0 41308 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_444
timestamp 1644511149
transform 1 0 41952 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_449
timestamp 1644511149
transform 1 0 42412 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_9
timestamp 1644511149
transform 1 0 1932 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_13
timestamp 1644511149
transform 1 0 2300 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_20
timestamp 1644511149
transform 1 0 2944 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_45
timestamp 1644511149
transform 1 0 5244 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_57
timestamp 1644511149
transform 1 0 6348 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_69
timestamp 1644511149
transform 1 0 7452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_81
timestamp 1644511149
transform 1 0 8556 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_157
timestamp 1644511149
transform 1 0 15548 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_166
timestamp 1644511149
transform 1 0 16376 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_170
timestamp 1644511149
transform 1 0 16744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_176
timestamp 1644511149
transform 1 0 17296 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_186
timestamp 1644511149
transform 1 0 18216 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_194
timestamp 1644511149
transform 1 0 18952 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_200
timestamp 1644511149
transform 1 0 19504 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_212
timestamp 1644511149
transform 1 0 20608 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_224
timestamp 1644511149
transform 1 0 21712 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_230
timestamp 1644511149
transform 1 0 22264 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_247
timestamp 1644511149
transform 1 0 23828 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1644511149
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_259
timestamp 1644511149
transform 1 0 24932 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_271
timestamp 1644511149
transform 1 0 26036 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_278
timestamp 1644511149
transform 1 0 26680 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_290
timestamp 1644511149
transform 1 0 27784 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_302
timestamp 1644511149
transform 1 0 28888 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_62_312
timestamp 1644511149
transform 1 0 29808 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_325
timestamp 1644511149
transform 1 0 31004 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_337
timestamp 1644511149
transform 1 0 32108 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_345
timestamp 1644511149
transform 1 0 32844 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_352
timestamp 1644511149
transform 1 0 33488 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_360
timestamp 1644511149
transform 1 0 34224 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_373
timestamp 1644511149
transform 1 0 35420 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_381
timestamp 1644511149
transform 1 0 36156 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_398
timestamp 1644511149
transform 1 0 37720 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_406
timestamp 1644511149
transform 1 0 38456 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_414
timestamp 1644511149
transform 1 0 39192 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_421
timestamp 1644511149
transform 1 0 39836 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_425
timestamp 1644511149
transform 1 0 40204 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_447
timestamp 1644511149
transform 1 0 42228 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_63_12
timestamp 1644511149
transform 1 0 2208 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_18
timestamp 1644511149
transform 1 0 2760 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_28
timestamp 1644511149
transform 1 0 3680 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_44
timestamp 1644511149
transform 1 0 5152 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_52
timestamp 1644511149
transform 1 0 5888 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_141
timestamp 1644511149
transform 1 0 14076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_146
timestamp 1644511149
transform 1 0 14536 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_154
timestamp 1644511149
transform 1 0 15272 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_181
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_185
timestamp 1644511149
transform 1 0 18124 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_191
timestamp 1644511149
transform 1 0 18676 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_203
timestamp 1644511149
transform 1 0 19780 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_207
timestamp 1644511149
transform 1 0 20148 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_211
timestamp 1644511149
transform 1 0 20516 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_219
timestamp 1644511149
transform 1 0 21252 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1644511149
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_225
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_231
timestamp 1644511149
transform 1 0 22356 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_236
timestamp 1644511149
transform 1 0 22816 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_246
timestamp 1644511149
transform 1 0 23736 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_260
timestamp 1644511149
transform 1 0 25024 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_269
timestamp 1644511149
transform 1 0 25852 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_276
timestamp 1644511149
transform 1 0 26496 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_293
timestamp 1644511149
transform 1 0 28060 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_298
timestamp 1644511149
transform 1 0 28520 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_305
timestamp 1644511149
transform 1 0 29164 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_314
timestamp 1644511149
transform 1 0 29992 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_326
timestamp 1644511149
transform 1 0 31096 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_331
timestamp 1644511149
transform 1 0 31556 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1644511149
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_350
timestamp 1644511149
transform 1 0 33304 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_362
timestamp 1644511149
transform 1 0 34408 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_63_386
timestamp 1644511149
transform 1 0 36616 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_401
timestamp 1644511149
transform 1 0 37996 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_410
timestamp 1644511149
transform 1 0 38824 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_419
timestamp 1644511149
transform 1 0 39652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_431
timestamp 1644511149
transform 1 0 40756 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_439
timestamp 1644511149
transform 1 0 41492 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_443
timestamp 1644511149
transform 1 0 41860 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1644511149
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_449
timestamp 1644511149
transform 1 0 42412 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_24
timestamp 1644511149
transform 1 0 3312 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_45
timestamp 1644511149
transform 1 0 5244 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_57
timestamp 1644511149
transform 1 0 6348 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_69
timestamp 1644511149
transform 1 0 7452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_81
timestamp 1644511149
transform 1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_172
timestamp 1644511149
transform 1 0 16928 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_176
timestamp 1644511149
transform 1 0 17296 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_185
timestamp 1644511149
transform 1 0 18124 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_192
timestamp 1644511149
transform 1 0 18768 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_213
timestamp 1644511149
transform 1 0 20700 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_233
timestamp 1644511149
transform 1 0 22540 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1644511149
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1644511149
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_256
timestamp 1644511149
transform 1 0 24656 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_260
timestamp 1644511149
transform 1 0 25024 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_269
timestamp 1644511149
transform 1 0 25852 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_273
timestamp 1644511149
transform 1 0 26220 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_290
timestamp 1644511149
transform 1 0 27784 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_298
timestamp 1644511149
transform 1 0 28520 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_304
timestamp 1644511149
transform 1 0 29072 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_316
timestamp 1644511149
transform 1 0 30176 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_320
timestamp 1644511149
transform 1 0 30544 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_327
timestamp 1644511149
transform 1 0 31188 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_339
timestamp 1644511149
transform 1 0 32292 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_345
timestamp 1644511149
transform 1 0 32844 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_353
timestamp 1644511149
transform 1 0 33580 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_360
timestamp 1644511149
transform 1 0 34224 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_377
timestamp 1644511149
transform 1 0 35788 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_384
timestamp 1644511149
transform 1 0 36432 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_400
timestamp 1644511149
transform 1 0 37904 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_408
timestamp 1644511149
transform 1 0 38640 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_416
timestamp 1644511149
transform 1 0 39376 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_424
timestamp 1644511149
transform 1 0 40112 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_436
timestamp 1644511149
transform 1 0 41216 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_443
timestamp 1644511149
transform 1 0 41860 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_3
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_65_9
timestamp 1644511149
transform 1 0 1932 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_15
timestamp 1644511149
transform 1 0 2484 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_37
timestamp 1644511149
transform 1 0 4508 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_49
timestamp 1644511149
transform 1 0 5612 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_93
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1644511149
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_122
timestamp 1644511149
transform 1 0 12328 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_134
timestamp 1644511149
transform 1 0 13432 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_146
timestamp 1644511149
transform 1 0 14536 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_158
timestamp 1644511149
transform 1 0 15640 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_166
timestamp 1644511149
transform 1 0 16376 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_65_169
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_65_191
timestamp 1644511149
transform 1 0 18676 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_203
timestamp 1644511149
transform 1 0 19780 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_215
timestamp 1644511149
transform 1 0 20884 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1644511149
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_241
timestamp 1644511149
transform 1 0 23276 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_65_253
timestamp 1644511149
transform 1 0 24380 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_259
timestamp 1644511149
transform 1 0 24932 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_276
timestamp 1644511149
transform 1 0 26496 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_281
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_289
timestamp 1644511149
transform 1 0 27692 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_308
timestamp 1644511149
transform 1 0 29440 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_328
timestamp 1644511149
transform 1 0 31280 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_65_344
timestamp 1644511149
transform 1 0 32752 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_350
timestamp 1644511149
transform 1 0 33304 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_367
timestamp 1644511149
transform 1 0 34868 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_379
timestamp 1644511149
transform 1 0 35972 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_65_386
timestamp 1644511149
transform 1 0 36616 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_65_393
timestamp 1644511149
transform 1 0 37260 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_401
timestamp 1644511149
transform 1 0 37996 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_406
timestamp 1644511149
transform 1 0 38456 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_416
timestamp 1644511149
transform 1 0 39376 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_436
timestamp 1644511149
transform 1 0 41216 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_443
timestamp 1644511149
transform 1 0 41860 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1644511149
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_449
timestamp 1644511149
transform 1 0 42412 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_66_3
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_66_9
timestamp 1644511149
transform 1 0 1932 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_15
timestamp 1644511149
transform 1 0 2484 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_19
timestamp 1644511149
transform 1 0 2852 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1644511149
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_32
timestamp 1644511149
transform 1 0 4048 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_44
timestamp 1644511149
transform 1 0 5152 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_56
timestamp 1644511149
transform 1 0 6256 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_68
timestamp 1644511149
transform 1 0 7360 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_80
timestamp 1644511149
transform 1 0 8464 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_91
timestamp 1644511149
transform 1 0 9476 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_103
timestamp 1644511149
transform 1 0 10580 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_118
timestamp 1644511149
transform 1 0 11960 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_130
timestamp 1644511149
transform 1 0 13064 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_138
timestamp 1644511149
transform 1 0 13800 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_153
timestamp 1644511149
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_165
timestamp 1644511149
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_177
timestamp 1644511149
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1644511149
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1644511149
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_197
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_209
timestamp 1644511149
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_221
timestamp 1644511149
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_233
timestamp 1644511149
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1644511149
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1644511149
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_253
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_263
timestamp 1644511149
transform 1 0 25300 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_66_274
timestamp 1644511149
transform 1 0 26312 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_286
timestamp 1644511149
transform 1 0 27416 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_298
timestamp 1644511149
transform 1 0 28520 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_306
timestamp 1644511149
transform 1 0 29256 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_309
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_313
timestamp 1644511149
transform 1 0 29900 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_317
timestamp 1644511149
transform 1 0 30268 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_321
timestamp 1644511149
transform 1 0 30636 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_327
timestamp 1644511149
transform 1 0 31188 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_338
timestamp 1644511149
transform 1 0 32200 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_342
timestamp 1644511149
transform 1 0 32568 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_359
timestamp 1644511149
transform 1 0 34132 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1644511149
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_365
timestamp 1644511149
transform 1 0 34684 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_373
timestamp 1644511149
transform 1 0 35420 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_390
timestamp 1644511149
transform 1 0 36984 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_66_412
timestamp 1644511149
transform 1 0 39008 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_421
timestamp 1644511149
transform 1 0 39836 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_425
timestamp 1644511149
transform 1 0 40204 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_447
timestamp 1644511149
transform 1 0 42228 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_6
timestamp 1644511149
transform 1 0 1656 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_13
timestamp 1644511149
transform 1 0 2300 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_25
timestamp 1644511149
transform 1 0 3404 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_32
timestamp 1644511149
transform 1 0 4048 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_38
timestamp 1644511149
transform 1 0 4600 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_42
timestamp 1644511149
transform 1 0 4968 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_54
timestamp 1644511149
transform 1 0 6072 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_95
timestamp 1644511149
transform 1 0 9844 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_108
timestamp 1644511149
transform 1 0 11040 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_125
timestamp 1644511149
transform 1 0 12604 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_132
timestamp 1644511149
transform 1 0 13248 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_144
timestamp 1644511149
transform 1 0 14352 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_156
timestamp 1644511149
transform 1 0 15456 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_181
timestamp 1644511149
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_193
timestamp 1644511149
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_205
timestamp 1644511149
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1644511149
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1644511149
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_225
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_237
timestamp 1644511149
transform 1 0 22908 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_244
timestamp 1644511149
transform 1 0 23552 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_256
timestamp 1644511149
transform 1 0 24656 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_268
timestamp 1644511149
transform 1 0 25760 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_281
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_293
timestamp 1644511149
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_305
timestamp 1644511149
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_317
timestamp 1644511149
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1644511149
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1644511149
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_337
timestamp 1644511149
transform 1 0 32108 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_348
timestamp 1644511149
transform 1 0 33120 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_355
timestamp 1644511149
transform 1 0 33764 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_367
timestamp 1644511149
transform 1 0 34868 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_374
timestamp 1644511149
transform 1 0 35512 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_378
timestamp 1644511149
transform 1 0 35880 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_383
timestamp 1644511149
transform 1 0 36340 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1644511149
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_393
timestamp 1644511149
transform 1 0 37260 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_399
timestamp 1644511149
transform 1 0 37812 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_403
timestamp 1644511149
transform 1 0 38180 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_415
timestamp 1644511149
transform 1 0 39284 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_419
timestamp 1644511149
transform 1 0 39652 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_444
timestamp 1644511149
transform 1 0 41952 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_449
timestamp 1644511149
transform 1 0 42412 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_24
timestamp 1644511149
transform 1 0 3312 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_32
timestamp 1644511149
transform 1 0 4048 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_68_59
timestamp 1644511149
transform 1 0 6532 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_71
timestamp 1644511149
transform 1 0 7636 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1644511149
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_68_91
timestamp 1644511149
transform 1 0 9476 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_103
timestamp 1644511149
transform 1 0 10580 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_116
timestamp 1644511149
transform 1 0 11776 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_122
timestamp 1644511149
transform 1 0 12328 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_126
timestamp 1644511149
transform 1 0 12696 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1644511149
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1644511149
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_144
timestamp 1644511149
transform 1 0 14352 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_156
timestamp 1644511149
transform 1 0 15456 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_168
timestamp 1644511149
transform 1 0 16560 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_180
timestamp 1644511149
transform 1 0 17664 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_192
timestamp 1644511149
transform 1 0 18768 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_197
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_209
timestamp 1644511149
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_221
timestamp 1644511149
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_233
timestamp 1644511149
transform 1 0 22540 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_238
timestamp 1644511149
transform 1 0 23000 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1644511149
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1644511149
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_253
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_265
timestamp 1644511149
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_280
timestamp 1644511149
transform 1 0 26864 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_292
timestamp 1644511149
transform 1 0 27968 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_304
timestamp 1644511149
transform 1 0 29072 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_309
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_321
timestamp 1644511149
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_333
timestamp 1644511149
transform 1 0 31740 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_341
timestamp 1644511149
transform 1 0 32476 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_68_346
timestamp 1644511149
transform 1 0 32936 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_354
timestamp 1644511149
transform 1 0 33672 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_359
timestamp 1644511149
transform 1 0 34132 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1644511149
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_368
timestamp 1644511149
transform 1 0 34960 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_379
timestamp 1644511149
transform 1 0 35972 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_386
timestamp 1644511149
transform 1 0 36616 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_398
timestamp 1644511149
transform 1 0 37720 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_410
timestamp 1644511149
transform 1 0 38824 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_416
timestamp 1644511149
transform 1 0 39376 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_421
timestamp 1644511149
transform 1 0 39836 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_425
timestamp 1644511149
transform 1 0 40204 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_432
timestamp 1644511149
transform 1 0 40848 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_439
timestamp 1644511149
transform 1 0 41492 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_446
timestamp 1644511149
transform 1 0 42136 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_450
timestamp 1644511149
transform 1 0 42504 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_69_3
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_27
timestamp 1644511149
transform 1 0 3588 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_34
timestamp 1644511149
transform 1 0 4232 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_41
timestamp 1644511149
transform 1 0 4876 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_47
timestamp 1644511149
transform 1 0 5428 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1644511149
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1644511149
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_60
timestamp 1644511149
transform 1 0 6624 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_72
timestamp 1644511149
transform 1 0 7728 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_69_84
timestamp 1644511149
transform 1 0 8832 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_108
timestamp 1644511149
transform 1 0 11040 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_113
timestamp 1644511149
transform 1 0 11500 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_135
timestamp 1644511149
transform 1 0 13524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_69_162
timestamp 1644511149
transform 1 0 16008 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_69_169
timestamp 1644511149
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_181
timestamp 1644511149
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_193
timestamp 1644511149
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_69_205
timestamp 1644511149
transform 1 0 19964 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_211
timestamp 1644511149
transform 1 0 20516 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1644511149
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_228
timestamp 1644511149
transform 1 0 22080 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_240
timestamp 1644511149
transform 1 0 23184 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_262
timestamp 1644511149
transform 1 0 25208 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1644511149
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1644511149
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_302
timestamp 1644511149
transform 1 0 28888 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_309
timestamp 1644511149
transform 1 0 29532 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_321
timestamp 1644511149
transform 1 0 30636 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_69_332
timestamp 1644511149
transform 1 0 31648 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_358
timestamp 1644511149
transform 1 0 34040 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_366
timestamp 1644511149
transform 1 0 34776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_388
timestamp 1644511149
transform 1 0 36800 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_393
timestamp 1644511149
transform 1 0 37260 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_401
timestamp 1644511149
transform 1 0 37996 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_69_406
timestamp 1644511149
transform 1 0 38456 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_414
timestamp 1644511149
transform 1 0 39192 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_419
timestamp 1644511149
transform 1 0 39652 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_444
timestamp 1644511149
transform 1 0 41952 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_449
timestamp 1644511149
transform 1 0 42412 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_24
timestamp 1644511149
transform 1 0 3312 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_70_29
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_35
timestamp 1644511149
transform 1 0 4324 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_60
timestamp 1644511149
transform 1 0 6624 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_72
timestamp 1644511149
transform 1 0 7728 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_89
timestamp 1644511149
transform 1 0 9292 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_96
timestamp 1644511149
transform 1 0 9936 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_103
timestamp 1644511149
transform 1 0 10580 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_128
timestamp 1644511149
transform 1 0 12880 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_132
timestamp 1644511149
transform 1 0 13248 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_136
timestamp 1644511149
transform 1 0 13616 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_162
timestamp 1644511149
transform 1 0 16008 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_174
timestamp 1644511149
transform 1 0 17112 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_186
timestamp 1644511149
transform 1 0 18216 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_194
timestamp 1644511149
transform 1 0 18952 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_197
timestamp 1644511149
transform 1 0 19228 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_205
timestamp 1644511149
transform 1 0 19964 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_228
timestamp 1644511149
transform 1 0 22080 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_235
timestamp 1644511149
transform 1 0 22724 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_242
timestamp 1644511149
transform 1 0 23368 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_250
timestamp 1644511149
transform 1 0 24104 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_274
timestamp 1644511149
transform 1 0 26312 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_299
timestamp 1644511149
transform 1 0 28612 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1644511149
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_330
timestamp 1644511149
transform 1 0 31464 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_338
timestamp 1644511149
transform 1 0 32200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_360
timestamp 1644511149
transform 1 0 34224 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_365
timestamp 1644511149
transform 1 0 34684 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_369
timestamp 1644511149
transform 1 0 35052 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_391
timestamp 1644511149
transform 1 0 37076 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_416
timestamp 1644511149
transform 1 0 39376 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_421
timestamp 1644511149
transform 1 0 39836 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_425
timestamp 1644511149
transform 1 0 40204 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_447
timestamp 1644511149
transform 1 0 42228 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_3
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_13
timestamp 1644511149
transform 1 0 2300 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_20
timestamp 1644511149
transform 1 0 2944 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_71_50
timestamp 1644511149
transform 1 0 5704 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1644511149
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_69
timestamp 1644511149
transform 1 0 7452 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_77
timestamp 1644511149
transform 1 0 8188 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_83
timestamp 1644511149
transform 1 0 8740 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_85
timestamp 1644511149
transform 1 0 8924 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_97
timestamp 1644511149
transform 1 0 10028 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_71_108
timestamp 1644511149
transform 1 0 11040 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_113
timestamp 1644511149
transform 1 0 11500 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_136
timestamp 1644511149
transform 1 0 13616 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_144
timestamp 1644511149
transform 1 0 14352 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_151
timestamp 1644511149
transform 1 0 14996 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_163
timestamp 1644511149
transform 1 0 16100 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1644511149
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_169
timestamp 1644511149
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_181
timestamp 1644511149
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_193
timestamp 1644511149
transform 1 0 18860 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_71_197
timestamp 1644511149
transform 1 0 19228 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_205
timestamp 1644511149
transform 1 0 19964 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_71_210
timestamp 1644511149
transform 1 0 20424 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_222
timestamp 1644511149
transform 1 0 21528 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_71_246
timestamp 1644511149
transform 1 0 23736 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_71_253
timestamp 1644511149
transform 1 0 24380 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_261
timestamp 1644511149
transform 1 0 25116 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_71_272
timestamp 1644511149
transform 1 0 26128 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_284
timestamp 1644511149
transform 1 0 27232 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_296
timestamp 1644511149
transform 1 0 28336 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_312
timestamp 1644511149
transform 1 0 29808 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_324
timestamp 1644511149
transform 1 0 30912 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_328
timestamp 1644511149
transform 1 0 31280 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_332
timestamp 1644511149
transform 1 0 31648 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_337
timestamp 1644511149
transform 1 0 32108 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_341
timestamp 1644511149
transform 1 0 32476 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_345
timestamp 1644511149
transform 1 0 32844 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_353
timestamp 1644511149
transform 1 0 33580 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_357
timestamp 1644511149
transform 1 0 33948 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_363
timestamp 1644511149
transform 1 0 34500 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_386
timestamp 1644511149
transform 1 0 36616 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_71_393
timestamp 1644511149
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_405
timestamp 1644511149
transform 1 0 38364 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_409
timestamp 1644511149
transform 1 0 38732 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_416
timestamp 1644511149
transform 1 0 39376 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_421
timestamp 1644511149
transform 1 0 39836 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_444
timestamp 1644511149
transform 1 0 41952 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_449
timestamp 1644511149
transform 1 0 42412 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 42872 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 42872 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 42872 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 42872 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 42872 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 42872 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 42872 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 42872 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 42872 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 42872 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 42872 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 42872 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 42872 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 42872 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 42872 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 42872 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 42872 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 42872 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 42872 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 42872 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 42872 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 42872 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 42872 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 42872 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 42872 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 42872 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 42872 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 42872 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 42872 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 42872 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 42872 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 42872 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 42872 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 42872 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 42872 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 42872 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 42872 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 42872 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 42872 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 42872 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 42872 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 42872 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 42872 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 42872 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 42872 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 42872 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 42872 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 42872 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 42872 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 42872 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 42872 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 42872 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 42872 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 42872 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 42872 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 42872 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 42872 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 42872 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 42872 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 42872 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 42872 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 42872 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 42872 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 42872 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 42872 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 42872 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 42872 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 42872 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 42872 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 42872 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 42872 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 42872 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 3680 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 8832 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 13984 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 19136 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 24288 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 29440 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 34592 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 39744 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _0951_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10212 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _0952_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  _0953_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0954_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 41492 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0955_
timestamp 1644511149
transform 1 0 20240 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0956_
timestamp 1644511149
transform 1 0 41400 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0957_
timestamp 1644511149
transform -1 0 4048 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0958_
timestamp 1644511149
transform 1 0 41400 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0959_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8740 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0960_
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0961_
timestamp 1644511149
transform -1 0 4324 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0962_
timestamp 1644511149
transform 1 0 29256 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0963_
timestamp 1644511149
transform 1 0 41860 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0964_
timestamp 1644511149
transform -1 0 41584 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0965_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10212 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _0966_
timestamp 1644511149
transform -1 0 11776 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0967_
timestamp 1644511149
transform -1 0 5704 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0968_
timestamp 1644511149
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0969_
timestamp 1644511149
transform -1 0 2300 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0970_
timestamp 1644511149
transform 1 0 39100 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp 1644511149
transform -1 0 2208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0972_
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0973_
timestamp 1644511149
transform 1 0 41308 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0974_
timestamp 1644511149
transform -1 0 41032 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0975_
timestamp 1644511149
transform -1 0 11040 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0976_
timestamp 1644511149
transform 1 0 26588 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0977_
timestamp 1644511149
transform 1 0 41584 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0978_
timestamp 1644511149
transform -1 0 11040 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0979_
timestamp 1644511149
transform -1 0 2392 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0980_
timestamp 1644511149
transform 1 0 41400 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0981_
timestamp 1644511149
transform 1 0 4692 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0982_
timestamp 1644511149
transform 1 0 41400 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0983_
timestamp 1644511149
transform -1 0 3036 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0984_
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0985_
timestamp 1644511149
transform -1 0 2208 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0986_
timestamp 1644511149
transform -1 0 2208 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0987_
timestamp 1644511149
transform 1 0 9200 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0988_
timestamp 1644511149
transform 1 0 37812 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0989_
timestamp 1644511149
transform -1 0 2208 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0990_
timestamp 1644511149
transform 1 0 10856 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0991_
timestamp 1644511149
transform -1 0 35972 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0992_
timestamp 1644511149
transform -1 0 10304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0993_
timestamp 1644511149
transform 1 0 41308 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0994_
timestamp 1644511149
transform 1 0 41400 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0995_
timestamp 1644511149
transform 1 0 22724 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0996_
timestamp 1644511149
transform -1 0 5888 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  _0997_
timestamp 1644511149
transform 1 0 4048 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0998_
timestamp 1644511149
transform 1 0 21804 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0999_
timestamp 1644511149
transform -1 0 4324 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1000_
timestamp 1644511149
transform -1 0 4232 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1001_
timestamp 1644511149
transform 1 0 40940 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1002_
timestamp 1644511149
transform 1 0 12420 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1003_
timestamp 1644511149
transform 1 0 4140 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1004_
timestamp 1644511149
transform 1 0 31372 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1005_
timestamp 1644511149
transform -1 0 11776 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1006_
timestamp 1644511149
transform 1 0 37812 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1007_
timestamp 1644511149
transform 1 0 13064 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1008_
timestamp 1644511149
transform -1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1009_
timestamp 1644511149
transform -1 0 3680 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_2  _1010_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34684 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1011_
timestamp 1644511149
transform -1 0 4876 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1012_
timestamp 1644511149
transform 1 0 41308 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1013_
timestamp 1644511149
transform -1 0 40848 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1014_
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1015_
timestamp 1644511149
transform -1 0 5244 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1016_
timestamp 1644511149
transform 1 0 41676 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1017_
timestamp 1644511149
transform 1 0 41584 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1018_
timestamp 1644511149
transform -1 0 41768 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1019_
timestamp 1644511149
transform -1 0 2208 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1020_
timestamp 1644511149
transform -1 0 2300 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1021_
timestamp 1644511149
transform -1 0 5336 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1022_
timestamp 1644511149
transform -1 0 2300 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1023_
timestamp 1644511149
transform 1 0 41308 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1024_
timestamp 1644511149
transform -1 0 2208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1025_
timestamp 1644511149
transform 1 0 41308 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1026_
timestamp 1644511149
transform 1 0 23276 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1027_
timestamp 1644511149
transform 1 0 5520 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _1028_
timestamp 1644511149
transform 1 0 6072 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1029_
timestamp 1644511149
transform -1 0 5796 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1030_
timestamp 1644511149
transform -1 0 15364 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1031_
timestamp 1644511149
transform 1 0 34684 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1032_
timestamp 1644511149
transform -1 0 20700 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1033_
timestamp 1644511149
transform 1 0 33856 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1034_
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1035_
timestamp 1644511149
transform 1 0 41308 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1036_
timestamp 1644511149
transform 1 0 39928 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1037_
timestamp 1644511149
transform 1 0 25944 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1038_
timestamp 1644511149
transform -1 0 2944 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1039_
timestamp 1644511149
transform 1 0 41308 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1040_
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1041_
timestamp 1644511149
transform 1 0 36340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1042_
timestamp 1644511149
transform -1 0 2300 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1043_
timestamp 1644511149
transform -1 0 32936 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1044_
timestamp 1644511149
transform -1 0 18676 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1045_
timestamp 1644511149
transform -1 0 2944 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _1046_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6164 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _1047_
timestamp 1644511149
transform 1 0 23552 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1048_
timestamp 1644511149
transform 1 0 41584 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1049_
timestamp 1644511149
transform 1 0 27784 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1050_
timestamp 1644511149
transform -1 0 2944 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1051_
timestamp 1644511149
transform -1 0 35972 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1052_
timestamp 1644511149
transform -1 0 5796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1053_
timestamp 1644511149
transform -1 0 2852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1054_
timestamp 1644511149
transform 1 0 39100 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1055_
timestamp 1644511149
transform 1 0 39100 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1056_
timestamp 1644511149
transform 1 0 40848 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1057_
timestamp 1644511149
transform 1 0 3312 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1058_
timestamp 1644511149
transform 1 0 10488 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1059_
timestamp 1644511149
transform -1 0 41400 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1060_
timestamp 1644511149
transform 1 0 37168 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1061_
timestamp 1644511149
transform -1 0 12236 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1062_
timestamp 1644511149
transform -1 0 12880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1063_
timestamp 1644511149
transform 1 0 41492 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1064_
timestamp 1644511149
transform 1 0 10948 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1065_
timestamp 1644511149
transform -1 0 2944 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1066_
timestamp 1644511149
transform 1 0 41400 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1067_
timestamp 1644511149
transform -1 0 41676 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1068_
timestamp 1644511149
transform 1 0 41768 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1069_
timestamp 1644511149
transform -1 0 9476 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1070_
timestamp 1644511149
transform 1 0 10948 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1071_
timestamp 1644511149
transform 1 0 10304 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1072_
timestamp 1644511149
transform -1 0 2392 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1073_
timestamp 1644511149
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1074_
timestamp 1644511149
transform 1 0 13340 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1075_
timestamp 1644511149
transform -1 0 2300 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1076_
timestamp 1644511149
transform -1 0 11684 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1077_
timestamp 1644511149
transform 1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1078_
timestamp 1644511149
transform -1 0 40940 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1079_
timestamp 1644511149
transform 1 0 41952 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1080_
timestamp 1644511149
transform -1 0 16928 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1081_
timestamp 1644511149
transform -1 0 3036 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1082_
timestamp 1644511149
transform 1 0 22632 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1083_
timestamp 1644511149
transform 1 0 38180 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1084_
timestamp 1644511149
transform -1 0 8280 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1085_
timestamp 1644511149
transform 1 0 25944 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1086_
timestamp 1644511149
transform 1 0 27508 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1087_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25484 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__nor4_1  _1088_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24196 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1089_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24472 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1090_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 24380 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_2  _1091_
timestamp 1644511149
transform -1 0 26496 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1092_
timestamp 1644511149
transform -1 0 34960 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1093_
timestamp 1644511149
transform 1 0 25024 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1094_
timestamp 1644511149
transform 1 0 25208 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1095_
timestamp 1644511149
transform 1 0 24472 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2b_1  _1096_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27692 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1097_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27048 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1098_
timestamp 1644511149
transform 1 0 27324 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1099_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28612 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1100_
timestamp 1644511149
transform 1 0 30360 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1101_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25760 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1102_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26772 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1103_
timestamp 1644511149
transform 1 0 27784 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1104_
timestamp 1644511149
transform -1 0 28796 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1105_
timestamp 1644511149
transform -1 0 29808 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1106_
timestamp 1644511149
transform -1 0 27232 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _1107_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 27324 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1108_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28152 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _1109_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 26036 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1110_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 24656 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1111_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 24104 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1112_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 27140 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1113_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__o22ai_1  _1114_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1115_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28152 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1116_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29532 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1117_
timestamp 1644511149
transform 1 0 30636 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1118_
timestamp 1644511149
transform 1 0 30728 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1119_
timestamp 1644511149
transform 1 0 28612 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1120_
timestamp 1644511149
transform -1 0 29072 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1121_
timestamp 1644511149
transform 1 0 26680 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1122_
timestamp 1644511149
transform -1 0 23460 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _1123_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 25668 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1124_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1125_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 28888 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _1126_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 29992 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1127_
timestamp 1644511149
transform 1 0 30728 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1128_
timestamp 1644511149
transform -1 0 30452 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1129_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 30360 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1130_
timestamp 1644511149
transform -1 0 28980 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1131_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 26036 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1132_
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1133_
timestamp 1644511149
transform 1 0 28888 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1134_
timestamp 1644511149
transform 1 0 26588 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1135_
timestamp 1644511149
transform 1 0 23000 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1136_
timestamp 1644511149
transform 1 0 22448 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1137_
timestamp 1644511149
transform -1 0 23920 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o22ai_1  _1138_
timestamp 1644511149
transform 1 0 26036 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1139_
timestamp 1644511149
transform 1 0 30728 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1140_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1141_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30360 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _1142_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1143_
timestamp 1644511149
transform 1 0 30636 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1144_
timestamp 1644511149
transform 1 0 30452 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1145_
timestamp 1644511149
transform -1 0 28796 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _1146_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 29256 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1147_
timestamp 1644511149
transform 1 0 29624 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _1148_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1149_
timestamp 1644511149
transform 1 0 28612 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1150_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29164 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _1151_
timestamp 1644511149
transform 1 0 24288 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1152_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1153_
timestamp 1644511149
transform 1 0 26404 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1154_
timestamp 1644511149
transform 1 0 27232 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or3_2  _1155_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25208 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _1156_
timestamp 1644511149
transform -1 0 26036 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _1157_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30728 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _1158_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25300 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1159_
timestamp 1644511149
transform -1 0 35052 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _1160_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30636 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1161_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 33028 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_2  _1162_
timestamp 1644511149
transform -1 0 32844 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1163_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24840 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1164_
timestamp 1644511149
transform 1 0 30084 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1165_
timestamp 1644511149
transform 1 0 30728 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1166_
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1167_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31924 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1168_
timestamp 1644511149
transform -1 0 34224 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1169_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 33764 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1170_
timestamp 1644511149
transform 1 0 33212 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1171_
timestamp 1644511149
transform 1 0 34224 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1172_
timestamp 1644511149
transform 1 0 33580 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1173_
timestamp 1644511149
transform -1 0 35052 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1174_
timestamp 1644511149
transform 1 0 34960 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1175_
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1176_
timestamp 1644511149
transform -1 0 35144 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1177_
timestamp 1644511149
transform 1 0 35604 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__xor2_1  _1178_
timestamp 1644511149
transform 1 0 35236 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1179_
timestamp 1644511149
transform 1 0 35972 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1180_
timestamp 1644511149
transform 1 0 35604 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1181_
timestamp 1644511149
transform -1 0 37076 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1182_
timestamp 1644511149
transform -1 0 35144 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1183_
timestamp 1644511149
transform 1 0 24748 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1184_
timestamp 1644511149
transform -1 0 24932 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1185_
timestamp 1644511149
transform 1 0 25208 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1186_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25300 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1187_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 26588 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1188_
timestamp 1644511149
transform 1 0 30084 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1189_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 31648 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1190_
timestamp 1644511149
transform 1 0 29900 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _1191_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1192_
timestamp 1644511149
transform 1 0 24840 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1193_
timestamp 1644511149
transform 1 0 28428 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1194_
timestamp 1644511149
transform 1 0 29992 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1195_
timestamp 1644511149
transform 1 0 35420 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1196_
timestamp 1644511149
transform -1 0 35144 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1197_
timestamp 1644511149
transform 1 0 35788 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1198_
timestamp 1644511149
transform 1 0 36800 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _1199_
timestamp 1644511149
transform 1 0 33304 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1200_
timestamp 1644511149
transform 1 0 36708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1201_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 34684 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1202_
timestamp 1644511149
transform -1 0 37996 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _1203_
timestamp 1644511149
transform -1 0 35328 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1204_
timestamp 1644511149
transform -1 0 34040 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1205_
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1206_
timestamp 1644511149
transform 1 0 30912 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _1207_
timestamp 1644511149
transform 1 0 32476 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1208_
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1209_
timestamp 1644511149
transform -1 0 36156 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1210_
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1211_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1212_
timestamp 1644511149
transform 1 0 35328 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1213_
timestamp 1644511149
transform 1 0 37352 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1214_
timestamp 1644511149
transform 1 0 34868 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1215_
timestamp 1644511149
transform -1 0 33856 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1216_
timestamp 1644511149
transform 1 0 32936 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1217_
timestamp 1644511149
transform 1 0 33580 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1218_
timestamp 1644511149
transform 1 0 36524 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1219_
timestamp 1644511149
transform -1 0 36708 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1220_
timestamp 1644511149
transform 1 0 32844 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1221_
timestamp 1644511149
transform 1 0 31924 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1222_
timestamp 1644511149
transform 1 0 30452 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1223_
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1224_
timestamp 1644511149
transform 1 0 37444 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1225_
timestamp 1644511149
transform 1 0 35696 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1226_
timestamp 1644511149
transform 1 0 35696 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1227_
timestamp 1644511149
transform 1 0 35052 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1228_
timestamp 1644511149
transform 1 0 35604 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1229_
timestamp 1644511149
transform 1 0 34500 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1230_
timestamp 1644511149
transform 1 0 32568 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1231_
timestamp 1644511149
transform 1 0 31372 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1232_
timestamp 1644511149
transform 1 0 33580 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1233_
timestamp 1644511149
transform -1 0 34132 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1234_
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1235_
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1236_
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1237_
timestamp 1644511149
transform 1 0 34684 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1238_
timestamp 1644511149
transform -1 0 37720 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1239_
timestamp 1644511149
transform 1 0 35972 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1240_
timestamp 1644511149
transform 1 0 35696 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1241_
timestamp 1644511149
transform -1 0 35788 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1242_
timestamp 1644511149
transform 1 0 36156 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1243_
timestamp 1644511149
transform 1 0 36248 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1244_
timestamp 1644511149
transform 1 0 38456 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1245_
timestamp 1644511149
transform -1 0 38180 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1246_
timestamp 1644511149
transform -1 0 38088 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1247_
timestamp 1644511149
transform -1 0 15456 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1248_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15088 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1249_
timestamp 1644511149
transform -1 0 17664 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1250_
timestamp 1644511149
transform 1 0 18768 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1251_
timestamp 1644511149
transform 1 0 20792 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1252_
timestamp 1644511149
transform 1 0 21528 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1253_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22356 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1254_
timestamp 1644511149
transform 1 0 38456 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1255_
timestamp 1644511149
transform -1 0 38088 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1256_
timestamp 1644511149
transform 1 0 37444 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1257_
timestamp 1644511149
transform -1 0 41032 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1258_
timestamp 1644511149
transform -1 0 38364 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1259_
timestamp 1644511149
transform -1 0 39100 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1260_
timestamp 1644511149
transform -1 0 37812 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1261_
timestamp 1644511149
transform -1 0 40480 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1262_
timestamp 1644511149
transform -1 0 39376 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1263_
timestamp 1644511149
transform 1 0 38916 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1264_
timestamp 1644511149
transform -1 0 39560 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1265_
timestamp 1644511149
transform 1 0 38824 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1266_
timestamp 1644511149
transform -1 0 39652 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1267_
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1268_
timestamp 1644511149
transform 1 0 20240 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1269_
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _1270_
timestamp 1644511149
transform -1 0 15916 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1271_
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1272_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 16192 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1273_
timestamp 1644511149
transform 1 0 12696 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1274_
timestamp 1644511149
transform -1 0 14536 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1275_
timestamp 1644511149
transform 1 0 15180 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1276_
timestamp 1644511149
transform 1 0 16836 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1277_
timestamp 1644511149
transform 1 0 18584 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1278_
timestamp 1644511149
transform 1 0 15364 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1279_
timestamp 1644511149
transform -1 0 19136 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1280_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17572 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1281_
timestamp 1644511149
transform 1 0 15272 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__or3_1  _1282_
timestamp 1644511149
transform 1 0 15640 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1283_
timestamp 1644511149
transform -1 0 17296 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1284_
timestamp 1644511149
transform 1 0 12144 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1285_
timestamp 1644511149
transform 1 0 26220 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1286_
timestamp 1644511149
transform 1 0 37536 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1287_
timestamp 1644511149
transform -1 0 38732 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_1  _1288_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 37260 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1289_
timestamp 1644511149
transform -1 0 38456 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nor3b_1  _1290_
timestamp 1644511149
transform 1 0 36616 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1291_
timestamp 1644511149
transform 1 0 26036 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1292_
timestamp 1644511149
transform -1 0 27232 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1293_
timestamp 1644511149
transform 1 0 26128 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1294_
timestamp 1644511149
transform -1 0 27232 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1295_
timestamp 1644511149
transform 1 0 19964 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1296_
timestamp 1644511149
transform -1 0 20148 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1297_
timestamp 1644511149
transform 1 0 16100 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1298_
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1299_
timestamp 1644511149
transform -1 0 16652 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_2  _1300_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16100 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1301_
timestamp 1644511149
transform -1 0 17204 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1302_
timestamp 1644511149
transform 1 0 17664 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _1303_
timestamp 1644511149
transform 1 0 18216 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1304_
timestamp 1644511149
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1305_
timestamp 1644511149
transform -1 0 17388 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1306_
timestamp 1644511149
transform -1 0 17572 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1307_
timestamp 1644511149
transform 1 0 17112 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1308_
timestamp 1644511149
transform 1 0 20516 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1309_
timestamp 1644511149
transform 1 0 19504 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1310_
timestamp 1644511149
transform -1 0 20516 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1311_
timestamp 1644511149
transform -1 0 16284 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1312_
timestamp 1644511149
transform -1 0 15732 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1313_
timestamp 1644511149
transform -1 0 15916 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1314_
timestamp 1644511149
transform 1 0 14812 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1315_
timestamp 1644511149
transform 1 0 17756 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1316_
timestamp 1644511149
transform -1 0 18676 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1317_
timestamp 1644511149
transform -1 0 18584 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1318_
timestamp 1644511149
transform 1 0 17940 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1319_
timestamp 1644511149
transform -1 0 21252 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1320_
timestamp 1644511149
transform -1 0 19504 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1321_
timestamp 1644511149
transform 1 0 19596 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1322_
timestamp 1644511149
transform -1 0 21344 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1323_
timestamp 1644511149
transform -1 0 19504 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1324_
timestamp 1644511149
transform 1 0 19504 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1325_
timestamp 1644511149
transform 1 0 19044 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1326_
timestamp 1644511149
transform 1 0 21620 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1327_
timestamp 1644511149
transform -1 0 20608 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1328_
timestamp 1644511149
transform -1 0 18308 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1329_
timestamp 1644511149
transform 1 0 18032 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1330_
timestamp 1644511149
transform -1 0 17664 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1331_
timestamp 1644511149
transform 1 0 14720 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1332_
timestamp 1644511149
transform 1 0 14904 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1333_
timestamp 1644511149
transform -1 0 18124 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1334_
timestamp 1644511149
transform 1 0 31280 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1335_
timestamp 1644511149
transform -1 0 24840 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1336_
timestamp 1644511149
transform 1 0 32292 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1337_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 38456 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _1338_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 37168 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _1339_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 37996 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1340_
timestamp 1644511149
transform 1 0 39100 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1341_
timestamp 1644511149
transform 1 0 32752 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1342_
timestamp 1644511149
transform -1 0 29992 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1343_
timestamp 1644511149
transform 1 0 30544 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _1344_
timestamp 1644511149
transform 1 0 31556 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _1345_
timestamp 1644511149
transform -1 0 34868 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1346_
timestamp 1644511149
transform 1 0 32108 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _1347_
timestamp 1644511149
transform 1 0 33028 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1348_
timestamp 1644511149
transform 1 0 28520 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1349_
timestamp 1644511149
transform 1 0 29900 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1350_
timestamp 1644511149
transform 1 0 29624 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1351_
timestamp 1644511149
transform 1 0 29992 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1352_
timestamp 1644511149
transform 1 0 28520 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1353_
timestamp 1644511149
transform -1 0 28796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1354_
timestamp 1644511149
transform -1 0 29164 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1355_
timestamp 1644511149
transform -1 0 29072 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1356_
timestamp 1644511149
transform 1 0 28244 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1357_
timestamp 1644511149
transform 1 0 30728 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1358_
timestamp 1644511149
transform -1 0 31188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1359_
timestamp 1644511149
transform -1 0 32844 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _1360_
timestamp 1644511149
transform 1 0 32108 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1361_
timestamp 1644511149
transform -1 0 33764 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1362_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31556 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1363_
timestamp 1644511149
transform 1 0 32384 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1364_
timestamp 1644511149
transform 1 0 32660 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1365_
timestamp 1644511149
transform 1 0 32936 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1366_
timestamp 1644511149
transform -1 0 34224 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1367_
timestamp 1644511149
transform 1 0 32936 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1368_
timestamp 1644511149
transform 1 0 33120 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1369_
timestamp 1644511149
transform 1 0 33856 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1370_
timestamp 1644511149
transform -1 0 33580 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1371_
timestamp 1644511149
transform 1 0 31832 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1372_
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1373_
timestamp 1644511149
transform 1 0 33948 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1374_
timestamp 1644511149
transform 1 0 29900 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1375_
timestamp 1644511149
transform 1 0 29808 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1376_
timestamp 1644511149
transform -1 0 32752 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1377_
timestamp 1644511149
transform 1 0 30636 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1378_
timestamp 1644511149
transform 1 0 30820 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1379_
timestamp 1644511149
transform -1 0 30912 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1380_
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1381_
timestamp 1644511149
transform -1 0 31188 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1382_
timestamp 1644511149
transform 1 0 31372 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1383_
timestamp 1644511149
transform -1 0 31556 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1384_
timestamp 1644511149
transform 1 0 29716 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1385_
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1386_
timestamp 1644511149
transform -1 0 31556 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1387_
timestamp 1644511149
transform -1 0 30820 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1388_
timestamp 1644511149
transform 1 0 32292 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1389_
timestamp 1644511149
transform 1 0 33304 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1390_
timestamp 1644511149
transform -1 0 32936 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1391_
timestamp 1644511149
transform 1 0 32660 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1392_
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1393_
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1394_
timestamp 1644511149
transform 1 0 35696 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1395_
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1396_
timestamp 1644511149
transform -1 0 33856 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1397_
timestamp 1644511149
transform -1 0 34868 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1398_
timestamp 1644511149
transform -1 0 34776 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1399_
timestamp 1644511149
transform 1 0 35236 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1400_
timestamp 1644511149
transform -1 0 37352 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1401_
timestamp 1644511149
transform 1 0 35512 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1402_
timestamp 1644511149
transform 1 0 36248 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1403_
timestamp 1644511149
transform -1 0 38732 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1404_
timestamp 1644511149
transform -1 0 36800 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1405_
timestamp 1644511149
transform 1 0 36524 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1406_
timestamp 1644511149
transform 1 0 38364 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1407_
timestamp 1644511149
transform -1 0 37996 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1408_
timestamp 1644511149
transform -1 0 38180 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1409_
timestamp 1644511149
transform 1 0 37812 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1410_
timestamp 1644511149
transform 1 0 38640 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1411_
timestamp 1644511149
transform 1 0 39836 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1412_
timestamp 1644511149
transform -1 0 38456 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1413_
timestamp 1644511149
transform 1 0 37904 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1414_
timestamp 1644511149
transform 1 0 39100 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1415_
timestamp 1644511149
transform 1 0 38824 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1416_
timestamp 1644511149
transform -1 0 40296 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1417_
timestamp 1644511149
transform -1 0 36340 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1418_
timestamp 1644511149
transform -1 0 35512 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1419_
timestamp 1644511149
transform 1 0 35512 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1420_
timestamp 1644511149
transform 1 0 37536 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1421_
timestamp 1644511149
transform 1 0 36800 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1422_
timestamp 1644511149
transform 1 0 37536 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1423_
timestamp 1644511149
transform -1 0 38916 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1424_
timestamp 1644511149
transform 1 0 38548 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1425_
timestamp 1644511149
transform -1 0 38824 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1426_
timestamp 1644511149
transform -1 0 40112 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1427_
timestamp 1644511149
transform -1 0 37720 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1428_
timestamp 1644511149
transform -1 0 39192 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1429_
timestamp 1644511149
transform -1 0 38456 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1430_
timestamp 1644511149
transform -1 0 39652 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1431_
timestamp 1644511149
transform -1 0 39376 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1432_
timestamp 1644511149
transform 1 0 38732 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1433_
timestamp 1644511149
transform -1 0 40112 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1434_
timestamp 1644511149
transform -1 0 38824 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1435_
timestamp 1644511149
transform -1 0 38456 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1436_
timestamp 1644511149
transform -1 0 38180 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1437_
timestamp 1644511149
transform -1 0 36616 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1438_
timestamp 1644511149
transform 1 0 35972 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1439_
timestamp 1644511149
transform 1 0 35880 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1440_
timestamp 1644511149
transform -1 0 36892 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1441_
timestamp 1644511149
transform -1 0 36156 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1442_
timestamp 1644511149
transform 1 0 35604 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1443_
timestamp 1644511149
transform -1 0 23828 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1444_
timestamp 1644511149
transform 1 0 21712 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1445_
timestamp 1644511149
transform 1 0 21252 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1446_
timestamp 1644511149
transform -1 0 22632 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1447_
timestamp 1644511149
transform 1 0 22080 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1448_
timestamp 1644511149
transform -1 0 23276 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1449_
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1450_
timestamp 1644511149
transform -1 0 22908 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1451_
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1452_
timestamp 1644511149
transform -1 0 23184 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1453_
timestamp 1644511149
transform 1 0 22908 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1454_
timestamp 1644511149
transform 1 0 23552 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1455_
timestamp 1644511149
transform 1 0 22632 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1456_
timestamp 1644511149
transform 1 0 22816 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1457_
timestamp 1644511149
transform -1 0 23920 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1458_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 25300 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1459_
timestamp 1644511149
transform -1 0 19964 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1460_
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1461_
timestamp 1644511149
transform 1 0 22724 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1462_
timestamp 1644511149
transform -1 0 28888 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _1463_
timestamp 1644511149
transform 1 0 21344 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1464_
timestamp 1644511149
transform -1 0 23644 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1465_
timestamp 1644511149
transform -1 0 20056 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1466_
timestamp 1644511149
transform 1 0 22724 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1467_
timestamp 1644511149
transform -1 0 20700 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _1468_
timestamp 1644511149
transform -1 0 20792 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1469_
timestamp 1644511149
transform 1 0 20424 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1470_
timestamp 1644511149
transform -1 0 22080 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21boi_1  _1471_
timestamp 1644511149
transform -1 0 21896 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1472_
timestamp 1644511149
transform -1 0 14904 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1473_
timestamp 1644511149
transform 1 0 17848 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1474_
timestamp 1644511149
transform 1 0 17848 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1475_
timestamp 1644511149
transform -1 0 18860 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1476_
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1477_
timestamp 1644511149
transform 1 0 20056 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1478_
timestamp 1644511149
transform 1 0 18492 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1479_
timestamp 1644511149
transform 1 0 19596 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1480_
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1481_
timestamp 1644511149
transform -1 0 20240 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1482_
timestamp 1644511149
transform 1 0 14536 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1483_
timestamp 1644511149
transform -1 0 19780 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1484_
timestamp 1644511149
transform 1 0 18032 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1485_
timestamp 1644511149
transform 1 0 20792 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1486_
timestamp 1644511149
transform -1 0 22080 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1487_
timestamp 1644511149
transform -1 0 13616 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1488_
timestamp 1644511149
transform -1 0 19504 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1489_
timestamp 1644511149
transform -1 0 22264 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1490_
timestamp 1644511149
transform -1 0 20424 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1491_
timestamp 1644511149
transform 1 0 13432 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1492_
timestamp 1644511149
transform -1 0 18032 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21boi_1  _1493_
timestamp 1644511149
transform -1 0 18492 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1494_
timestamp 1644511149
transform 1 0 17572 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1495_
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1496_
timestamp 1644511149
transform -1 0 20240 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1497_
timestamp 1644511149
transform -1 0 18584 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1498_
timestamp 1644511149
transform -1 0 21160 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1499_
timestamp 1644511149
transform 1 0 14812 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1500_
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1501_
timestamp 1644511149
transform 1 0 15916 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1502_
timestamp 1644511149
transform -1 0 16560 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1503_
timestamp 1644511149
transform 1 0 13248 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1504_
timestamp 1644511149
transform -1 0 17112 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1505_
timestamp 1644511149
transform 1 0 13340 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1506_
timestamp 1644511149
transform 1 0 18216 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1507_
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1508_
timestamp 1644511149
transform -1 0 16560 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1509_
timestamp 1644511149
transform 1 0 15456 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1510_
timestamp 1644511149
transform 1 0 15732 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _1511_
timestamp 1644511149
transform 1 0 17664 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1512_
timestamp 1644511149
transform -1 0 17112 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1513_
timestamp 1644511149
transform -1 0 17296 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1514_
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_2  _1515_
timestamp 1644511149
transform -1 0 17020 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1516_
timestamp 1644511149
transform 1 0 16468 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1517_
timestamp 1644511149
transform -1 0 29072 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _1518_
timestamp 1644511149
transform -1 0 23092 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1519_
timestamp 1644511149
transform 1 0 17388 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1520_
timestamp 1644511149
transform 1 0 17480 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1521_
timestamp 1644511149
transform -1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1522_
timestamp 1644511149
transform 1 0 15456 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1523_
timestamp 1644511149
transform -1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1524_
timestamp 1644511149
transform -1 0 15640 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1525_
timestamp 1644511149
transform -1 0 14720 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1526_
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1527_
timestamp 1644511149
transform -1 0 13064 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1528_
timestamp 1644511149
transform -1 0 14536 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1529_
timestamp 1644511149
transform -1 0 13616 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1530_
timestamp 1644511149
transform 1 0 13340 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1531_
timestamp 1644511149
transform 1 0 13248 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1532_
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1533_
timestamp 1644511149
transform 1 0 13156 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1534_
timestamp 1644511149
transform 1 0 14720 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _1535_
timestamp 1644511149
transform 1 0 14352 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1536_
timestamp 1644511149
transform -1 0 15824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1537_
timestamp 1644511149
transform -1 0 15732 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1538_
timestamp 1644511149
transform 1 0 18768 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1539_
timestamp 1644511149
transform -1 0 16008 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1540_
timestamp 1644511149
transform 1 0 15456 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1541_
timestamp 1644511149
transform 1 0 14352 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1542_
timestamp 1644511149
transform 1 0 17572 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1543_
timestamp 1644511149
transform -1 0 17296 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1544_
timestamp 1644511149
transform 1 0 15548 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_2  _1545_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15180 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__o31a_1  _1546_
timestamp 1644511149
transform -1 0 15824 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1547_
timestamp 1644511149
transform -1 0 25300 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1548_
timestamp 1644511149
transform -1 0 25668 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1549_
timestamp 1644511149
transform 1 0 23920 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1550_
timestamp 1644511149
transform 1 0 20792 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1551_
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_2  _1552_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 24656 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1553_
timestamp 1644511149
transform 1 0 23276 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1554_
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1555_
timestamp 1644511149
transform 1 0 16192 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1556_
timestamp 1644511149
transform 1 0 16928 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_1  _1557_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17020 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1558_
timestamp 1644511149
transform 1 0 20884 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1559_
timestamp 1644511149
transform -1 0 15180 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1560_
timestamp 1644511149
transform -1 0 16008 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1561_
timestamp 1644511149
transform -1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1562_
timestamp 1644511149
transform -1 0 14444 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1563_
timestamp 1644511149
transform -1 0 14996 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1564_
timestamp 1644511149
transform -1 0 16928 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1565_
timestamp 1644511149
transform 1 0 14536 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _1566_
timestamp 1644511149
transform -1 0 16652 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1567_
timestamp 1644511149
transform 1 0 15364 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1568_
timestamp 1644511149
transform -1 0 13616 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1569_
timestamp 1644511149
transform -1 0 15640 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1570_
timestamp 1644511149
transform 1 0 15180 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1571_
timestamp 1644511149
transform 1 0 14352 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1572_
timestamp 1644511149
transform -1 0 14812 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1573_
timestamp 1644511149
transform -1 0 13432 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1574_
timestamp 1644511149
transform 1 0 12512 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1575_
timestamp 1644511149
transform 1 0 15916 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1576_
timestamp 1644511149
transform -1 0 13616 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1577_
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _1578_
timestamp 1644511149
transform -1 0 16192 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1579_
timestamp 1644511149
transform 1 0 16744 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1580_
timestamp 1644511149
transform 1 0 16468 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1581_
timestamp 1644511149
transform -1 0 16928 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1582_
timestamp 1644511149
transform -1 0 14904 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1583_
timestamp 1644511149
transform 1 0 14444 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1584_
timestamp 1644511149
transform 1 0 14444 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1585_
timestamp 1644511149
transform 1 0 16192 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1586_
timestamp 1644511149
transform -1 0 17388 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1587_
timestamp 1644511149
transform -1 0 15456 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1588_
timestamp 1644511149
transform 1 0 17204 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1589_
timestamp 1644511149
transform 1 0 17756 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1590_
timestamp 1644511149
transform -1 0 15272 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1591_
timestamp 1644511149
transform -1 0 23828 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1592_
timestamp 1644511149
transform -1 0 15180 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1593_
timestamp 1644511149
transform 1 0 14260 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _1594_
timestamp 1644511149
transform 1 0 25024 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1595_
timestamp 1644511149
transform 1 0 24748 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1596_
timestamp 1644511149
transform 1 0 15640 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1597_
timestamp 1644511149
transform 1 0 17572 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1598_
timestamp 1644511149
transform -1 0 17848 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1599_
timestamp 1644511149
transform -1 0 17112 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1600_
timestamp 1644511149
transform 1 0 15088 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1601_
timestamp 1644511149
transform -1 0 16192 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1602_
timestamp 1644511149
transform -1 0 24656 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _1603_
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1604_
timestamp 1644511149
transform -1 0 17204 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1605_
timestamp 1644511149
transform -1 0 14536 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1606_
timestamp 1644511149
transform -1 0 13432 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1607_
timestamp 1644511149
transform -1 0 14628 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1608_
timestamp 1644511149
transform -1 0 14720 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _1609_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1610_
timestamp 1644511149
transform 1 0 22172 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1611_
timestamp 1644511149
transform -1 0 16928 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1612_
timestamp 1644511149
transform -1 0 19504 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1613_
timestamp 1644511149
transform 1 0 20056 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1614_
timestamp 1644511149
transform -1 0 22080 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _1615_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__o31a_1  _1616_
timestamp 1644511149
transform 1 0 17940 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1617_
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1618_
timestamp 1644511149
transform -1 0 17296 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1619_
timestamp 1644511149
transform -1 0 15640 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_1  _1620_
timestamp 1644511149
transform -1 0 14904 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1621_
timestamp 1644511149
transform -1 0 14904 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1622_
timestamp 1644511149
transform -1 0 16192 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1623_
timestamp 1644511149
transform -1 0 17204 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1624_
timestamp 1644511149
transform -1 0 14536 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1625_
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1626_
timestamp 1644511149
transform -1 0 16376 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _1627_
timestamp 1644511149
transform 1 0 15548 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1628_
timestamp 1644511149
transform -1 0 15916 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1629_
timestamp 1644511149
transform 1 0 16836 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1630_
timestamp 1644511149
transform 1 0 17664 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1631_
timestamp 1644511149
transform -1 0 17756 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1632_
timestamp 1644511149
transform -1 0 18124 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1633_
timestamp 1644511149
transform 1 0 18216 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1634_
timestamp 1644511149
transform -1 0 18768 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1635_
timestamp 1644511149
transform 1 0 17572 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1636_
timestamp 1644511149
transform 1 0 18124 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1637_
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1638_
timestamp 1644511149
transform 1 0 16376 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o221ai_1  _1639_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18124 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1640_
timestamp 1644511149
transform 1 0 19044 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1641_
timestamp 1644511149
transform 1 0 19320 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1642_
timestamp 1644511149
transform 1 0 19780 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1643_
timestamp 1644511149
transform 1 0 17848 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1644_
timestamp 1644511149
transform -1 0 19964 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1645_
timestamp 1644511149
transform 1 0 18492 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1646_
timestamp 1644511149
transform 1 0 18676 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1647_
timestamp 1644511149
transform 1 0 17664 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1648_
timestamp 1644511149
transform 1 0 18216 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1649_
timestamp 1644511149
transform -1 0 20792 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1650_
timestamp 1644511149
transform -1 0 21436 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1651_
timestamp 1644511149
transform 1 0 20700 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1652_
timestamp 1644511149
transform 1 0 20148 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1653_
timestamp 1644511149
transform -1 0 22264 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1654_
timestamp 1644511149
transform -1 0 21160 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1655_
timestamp 1644511149
transform 1 0 20424 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1656_
timestamp 1644511149
transform -1 0 23460 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1657_
timestamp 1644511149
transform 1 0 21344 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1658_
timestamp 1644511149
transform 1 0 20516 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1659_
timestamp 1644511149
transform 1 0 20792 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1660_
timestamp 1644511149
transform -1 0 20884 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1661_
timestamp 1644511149
transform 1 0 19504 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1662_
timestamp 1644511149
transform -1 0 21344 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1663_
timestamp 1644511149
transform -1 0 25208 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _1664_
timestamp 1644511149
transform 1 0 25760 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _1665_
timestamp 1644511149
transform 1 0 25668 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1666_
timestamp 1644511149
transform -1 0 25024 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1667_
timestamp 1644511149
transform -1 0 24656 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1668_
timestamp 1644511149
transform 1 0 24104 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1669_
timestamp 1644511149
transform -1 0 24012 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1670_
timestamp 1644511149
transform -1 0 23000 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_1  _1671_
timestamp 1644511149
transform -1 0 22724 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1672_
timestamp 1644511149
transform -1 0 22816 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1673_
timestamp 1644511149
transform 1 0 23368 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1674_
timestamp 1644511149
transform -1 0 24380 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1675_
timestamp 1644511149
transform -1 0 22264 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1676_
timestamp 1644511149
transform -1 0 26496 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1677_
timestamp 1644511149
transform -1 0 23736 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1678_
timestamp 1644511149
transform -1 0 23644 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1679_
timestamp 1644511149
transform -1 0 20516 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1680_
timestamp 1644511149
transform 1 0 25392 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1681_
timestamp 1644511149
transform 1 0 24748 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1682_
timestamp 1644511149
transform -1 0 24932 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1683_
timestamp 1644511149
transform -1 0 25852 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1684_
timestamp 1644511149
transform 1 0 25852 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1685_
timestamp 1644511149
transform -1 0 26680 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1686_
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1687_
timestamp 1644511149
transform -1 0 27600 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1688_
timestamp 1644511149
transform -1 0 26220 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1689_
timestamp 1644511149
transform -1 0 27232 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1690_
timestamp 1644511149
transform -1 0 27232 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1691_
timestamp 1644511149
transform 1 0 23460 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o221ai_1  _1692_
timestamp 1644511149
transform 1 0 25208 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1693_
timestamp 1644511149
transform 1 0 26588 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1694_
timestamp 1644511149
transform -1 0 26036 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1695_
timestamp 1644511149
transform 1 0 25484 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1696_
timestamp 1644511149
transform 1 0 23368 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1697_
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1698_
timestamp 1644511149
transform 1 0 25576 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1699_
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1700_
timestamp 1644511149
transform 1 0 23000 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1701_
timestamp 1644511149
transform 1 0 23644 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1702_
timestamp 1644511149
transform 1 0 26220 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1703_
timestamp 1644511149
transform 1 0 27784 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1704_
timestamp 1644511149
transform -1 0 27416 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1705_
timestamp 1644511149
transform 1 0 26312 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1706_
timestamp 1644511149
transform 1 0 26956 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1707_
timestamp 1644511149
transform -1 0 28060 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1708_
timestamp 1644511149
transform 1 0 25760 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1709_
timestamp 1644511149
transform -1 0 27232 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1710_
timestamp 1644511149
transform 1 0 25484 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1711_
timestamp 1644511149
transform 1 0 25668 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1712_
timestamp 1644511149
transform 1 0 27600 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1713_
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1714_
timestamp 1644511149
transform -1 0 26772 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1715_
timestamp 1644511149
transform 1 0 23644 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1716_
timestamp 1644511149
transform 1 0 30452 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _1717_
timestamp 1644511149
transform 1 0 30728 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__o21bai_1  _1718_
timestamp 1644511149
transform 1 0 30084 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1719_
timestamp 1644511149
transform 1 0 30912 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1720_
timestamp 1644511149
transform 1 0 32016 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1721_
timestamp 1644511149
transform -1 0 30176 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1722_
timestamp 1644511149
transform 1 0 28888 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1723_
timestamp 1644511149
transform -1 0 28244 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1724_
timestamp 1644511149
transform -1 0 30084 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _1725_
timestamp 1644511149
transform 1 0 28520 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1726_
timestamp 1644511149
transform -1 0 29900 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1727_
timestamp 1644511149
transform -1 0 28796 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1728_
timestamp 1644511149
transform -1 0 28520 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1729_
timestamp 1644511149
transform 1 0 27784 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1730_
timestamp 1644511149
transform -1 0 29992 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1731_
timestamp 1644511149
transform -1 0 28060 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1732_
timestamp 1644511149
transform -1 0 29072 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1733_
timestamp 1644511149
transform 1 0 28520 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1734_
timestamp 1644511149
transform -1 0 29072 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _1735_
timestamp 1644511149
transform 1 0 28336 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1736_
timestamp 1644511149
transform -1 0 29624 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1737_
timestamp 1644511149
transform -1 0 28704 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1738_
timestamp 1644511149
transform -1 0 29808 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1739_
timestamp 1644511149
transform -1 0 29808 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1740_
timestamp 1644511149
transform 1 0 33304 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1741_
timestamp 1644511149
transform -1 0 27600 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1742_
timestamp 1644511149
transform 1 0 26588 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1743_
timestamp 1644511149
transform -1 0 33580 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1744_
timestamp 1644511149
transform -1 0 31832 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1745_
timestamp 1644511149
transform -1 0 33028 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1746_
timestamp 1644511149
transform 1 0 31188 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1747_
timestamp 1644511149
transform -1 0 32936 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1748_
timestamp 1644511149
transform 1 0 32292 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1749_
timestamp 1644511149
transform -1 0 34224 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1750_
timestamp 1644511149
transform -1 0 32660 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1751_
timestamp 1644511149
transform 1 0 31096 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1752_
timestamp 1644511149
transform -1 0 23000 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1753_
timestamp 1644511149
transform -1 0 22908 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1754_
timestamp 1644511149
transform -1 0 25944 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1755_
timestamp 1644511149
transform 1 0 25944 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1756_
timestamp 1644511149
transform -1 0 27416 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1757_
timestamp 1644511149
transform -1 0 23736 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1758_
timestamp 1644511149
transform -1 0 23092 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _1759_
timestamp 1644511149
transform -1 0 25116 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1760_
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1761_
timestamp 1644511149
transform -1 0 25944 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1762_
timestamp 1644511149
transform 1 0 25484 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1763_
timestamp 1644511149
transform 1 0 25024 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1764_
timestamp 1644511149
transform -1 0 26312 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1765_
timestamp 1644511149
transform 1 0 25944 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1766_
timestamp 1644511149
transform 1 0 25852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1767_
timestamp 1644511149
transform 1 0 25852 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1768_
timestamp 1644511149
transform -1 0 27232 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1769_
timestamp 1644511149
transform -1 0 25484 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1770_
timestamp 1644511149
transform 1 0 24104 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1771_
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1772_
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1773_
timestamp 1644511149
transform -1 0 23000 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_1  _1774_
timestamp 1644511149
transform -1 0 21712 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1775_
timestamp 1644511149
transform 1 0 22080 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1776_
timestamp 1644511149
transform 1 0 20516 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1777_
timestamp 1644511149
transform 1 0 23368 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1778_
timestamp 1644511149
transform -1 0 21896 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1779_
timestamp 1644511149
transform -1 0 21252 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1780_
timestamp 1644511149
transform 1 0 20976 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1781_
timestamp 1644511149
transform 1 0 19964 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1782_
timestamp 1644511149
transform 1 0 20240 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1783_
timestamp 1644511149
transform -1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1784_
timestamp 1644511149
transform 1 0 19504 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_4  _1785_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23828 0 -1 32640
box -38 -48 1602 592
use sky130_fd_sc_hd__xor2_1  _1786_
timestamp 1644511149
transform 1 0 21988 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1787_
timestamp 1644511149
transform -1 0 23828 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1788_
timestamp 1644511149
transform -1 0 23276 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1789_
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1790_
timestamp 1644511149
transform -1 0 20976 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1791_
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1792_
timestamp 1644511149
transform 1 0 20148 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1793_
timestamp 1644511149
transform -1 0 21160 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1794_
timestamp 1644511149
transform 1 0 20700 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1795_
timestamp 1644511149
transform 1 0 19596 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1796_
timestamp 1644511149
transform 1 0 19228 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1797_
timestamp 1644511149
transform -1 0 20056 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1798_
timestamp 1644511149
transform -1 0 18492 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1799_
timestamp 1644511149
transform 1 0 17848 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1800_
timestamp 1644511149
transform -1 0 32200 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1801_
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1802_
timestamp 1644511149
transform -1 0 32568 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1803_
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1804_
timestamp 1644511149
transform 1 0 30636 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1805_
timestamp 1644511149
transform -1 0 31648 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1806_
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1807_
timestamp 1644511149
transform 1 0 32108 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1808_
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1809_
timestamp 1644511149
transform 1 0 32568 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1810_
timestamp 1644511149
transform 1 0 33948 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1811_
timestamp 1644511149
transform -1 0 33856 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1812_
timestamp 1644511149
transform -1 0 32384 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1813_
timestamp 1644511149
transform -1 0 34132 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1814_
timestamp 1644511149
transform -1 0 33488 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1815_
timestamp 1644511149
transform 1 0 28796 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1816_
timestamp 1644511149
transform -1 0 29164 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1817_
timestamp 1644511149
transform 1 0 29992 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1818_
timestamp 1644511149
transform 1 0 30912 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1819_
timestamp 1644511149
transform 1 0 28336 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _1820_
timestamp 1644511149
transform -1 0 28796 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1821_
timestamp 1644511149
transform 1 0 26128 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1822_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 38732 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1823_
timestamp 1644511149
transform 1 0 36800 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1824_
timestamp 1644511149
transform 1 0 38824 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1825_
timestamp 1644511149
transform 1 0 33396 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1826_
timestamp 1644511149
transform 1 0 29348 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1827_
timestamp 1644511149
transform 1 0 31280 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1828_
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1829_
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1830_
timestamp 1644511149
transform 1 0 36340 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1831_
timestamp 1644511149
transform 1 0 31464 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1832_
timestamp 1644511149
transform -1 0 31004 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1833_
timestamp 1644511149
transform -1 0 31464 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1834_
timestamp 1644511149
transform 1 0 27324 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1835_
timestamp 1644511149
transform 1 0 37720 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1836_
timestamp 1644511149
transform 1 0 37536 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1837_
timestamp 1644511149
transform 1 0 27232 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1838_
timestamp 1644511149
transform -1 0 29072 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1839_
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1840_
timestamp 1644511149
transform 1 0 16836 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1841_
timestamp 1644511149
transform 1 0 21068 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1842_
timestamp 1644511149
transform 1 0 14720 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1843_
timestamp 1644511149
transform 1 0 14720 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1844_
timestamp 1644511149
transform 1 0 17296 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1845_
timestamp 1644511149
transform 1 0 19872 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1846_
timestamp 1644511149
transform -1 0 21344 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1847_
timestamp 1644511149
transform 1 0 14260 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1848_
timestamp 1644511149
transform 1 0 18308 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1849_
timestamp 1644511149
transform 1 0 29808 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1850_
timestamp 1644511149
transform 1 0 27968 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1851_
timestamp 1644511149
transform -1 0 34132 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1852_
timestamp 1644511149
transform -1 0 34868 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1853_
timestamp 1644511149
transform -1 0 34868 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1854_
timestamp 1644511149
transform -1 0 33396 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1855_
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1856_
timestamp 1644511149
transform 1 0 28428 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1857_
timestamp 1644511149
transform 1 0 29348 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1858_
timestamp 1644511149
transform 1 0 30728 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1859_
timestamp 1644511149
transform 1 0 32568 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1860_
timestamp 1644511149
transform 1 0 33856 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1861_
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1862_
timestamp 1644511149
transform -1 0 36800 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1863_
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1864_
timestamp 1644511149
transform 1 0 37536 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1865_
timestamp 1644511149
transform 1 0 39376 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1866_
timestamp 1644511149
transform 1 0 39928 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1867_
timestamp 1644511149
transform 1 0 34776 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1868_
timestamp 1644511149
transform -1 0 38088 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1869_
timestamp 1644511149
transform 1 0 39836 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1870_
timestamp 1644511149
transform 1 0 39836 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1871_
timestamp 1644511149
transform 1 0 39744 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1872_
timestamp 1644511149
transform -1 0 39008 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1873_
timestamp 1644511149
transform 1 0 35512 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1874_
timestamp 1644511149
transform 1 0 35144 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1875_
timestamp 1644511149
transform 1 0 22448 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1876_
timestamp 1644511149
transform -1 0 25760 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1877_
timestamp 1644511149
transform 1 0 23000 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1878_
timestamp 1644511149
transform 1 0 23276 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1879_
timestamp 1644511149
transform 1 0 23000 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1880_
timestamp 1644511149
transform 1 0 24288 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1881_
timestamp 1644511149
transform 1 0 22356 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1882_
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1883_
timestamp 1644511149
transform 1 0 20884 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1884_
timestamp 1644511149
transform 1 0 22356 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1885_
timestamp 1644511149
transform 1 0 18952 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1886_
timestamp 1644511149
transform 1 0 19596 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1887_
timestamp 1644511149
transform 1 0 19320 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1888_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20240 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1889_
timestamp 1644511149
transform 1 0 22448 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1890_
timestamp 1644511149
transform 1 0 22448 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1891_
timestamp 1644511149
transform 1 0 21988 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1892_
timestamp 1644511149
transform 1 0 19320 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1893_
timestamp 1644511149
transform 1 0 22540 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1894_
timestamp 1644511149
transform 1 0 22448 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1895_
timestamp 1644511149
transform 1 0 12880 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1896_
timestamp 1644511149
transform -1 0 15548 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1897_
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1898_
timestamp 1644511149
transform 1 0 17756 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1899_
timestamp 1644511149
transform 1 0 12880 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1900_
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1901_
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1902_
timestamp 1644511149
transform -1 0 12972 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1903_
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1904_
timestamp 1644511149
transform 1 0 14076 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1905_
timestamp 1644511149
transform -1 0 18768 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1906_
timestamp 1644511149
transform 1 0 14352 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1907_
timestamp 1644511149
transform 1 0 12880 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1908_
timestamp 1644511149
transform 1 0 12144 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1909_
timestamp 1644511149
transform 1 0 11868 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1910_
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1911_
timestamp 1644511149
transform 1 0 14444 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1912_
timestamp 1644511149
transform -1 0 18584 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1913_
timestamp 1644511149
transform 1 0 11684 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1914_
timestamp 1644511149
transform 1 0 12052 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1915_
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1916_
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1917_
timestamp 1644511149
transform 1 0 15456 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1918_
timestamp 1644511149
transform 1 0 17204 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1919_
timestamp 1644511149
transform -1 0 20700 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1920_
timestamp 1644511149
transform -1 0 19964 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1921_
timestamp 1644511149
transform 1 0 17204 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1922_
timestamp 1644511149
transform -1 0 22172 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1923_
timestamp 1644511149
transform 1 0 20424 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1924_
timestamp 1644511149
transform -1 0 22724 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1925_
timestamp 1644511149
transform 1 0 21804 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1926_
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1927_
timestamp 1644511149
transform 1 0 21068 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1928_
timestamp 1644511149
transform 1 0 25024 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1929_
timestamp 1644511149
transform 1 0 26312 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1930_
timestamp 1644511149
transform -1 0 24748 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1931_
timestamp 1644511149
transform 1 0 22448 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1932_
timestamp 1644511149
transform -1 0 28980 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1933_
timestamp 1644511149
transform -1 0 27232 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1934_
timestamp 1644511149
transform -1 0 28612 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1935_
timestamp 1644511149
transform 1 0 30360 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1936_
timestamp 1644511149
transform 1 0 28428 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1937_
timestamp 1644511149
transform 1 0 29624 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1938_
timestamp 1644511149
transform 1 0 30544 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1939_
timestamp 1644511149
transform -1 0 34868 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1940_
timestamp 1644511149
transform -1 0 36708 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1941_
timestamp 1644511149
transform 1 0 30820 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1942_
timestamp 1644511149
transform 1 0 23644 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1943_
timestamp 1644511149
transform 1 0 26036 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1944_
timestamp 1644511149
transform -1 0 27324 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1945_
timestamp 1644511149
transform 1 0 23828 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1946_
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1947_
timestamp 1644511149
transform 1 0 19596 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1948_
timestamp 1644511149
transform -1 0 20148 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1949_
timestamp 1644511149
transform 1 0 23092 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1950_
timestamp 1644511149
transform 1 0 21344 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1951_
timestamp 1644511149
transform 1 0 19504 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1952_
timestamp 1644511149
transform 1 0 17388 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1953_
timestamp 1644511149
transform 1 0 32752 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1954_
timestamp 1644511149
transform 1 0 31648 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1955_
timestamp 1644511149
transform 1 0 32200 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1956_
timestamp 1644511149
transform 1 0 29072 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1957_
timestamp 1644511149
transform -1 0 29348 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1958_
timestamp 1644511149
transform -1 0 27232 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1959_
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1960_
timestamp 1644511149
transform 1 0 27416 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1961_
timestamp 1644511149
transform 1 0 26680 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1962_
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1963_
timestamp 1644511149
transform 1 0 26036 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1964_
timestamp 1644511149
transform 1 0 25300 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1965_
timestamp 1644511149
transform 1 0 25392 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1966_
timestamp 1644511149
transform 1 0 35236 0 -1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1967_
timestamp 1644511149
transform -1 0 35236 0 -1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1968_
timestamp 1644511149
transform 1 0 34868 0 1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1969_
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1970_
timestamp 1644511149
transform 1 0 32752 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1971_
timestamp 1644511149
transform 1 0 33856 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1972_
timestamp 1644511149
transform -1 0 26312 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1973__6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 7544 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1974__7
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1975__8
timestamp 1644511149
transform -1 0 18400 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1976__9
timestamp 1644511149
transform 1 0 1472 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1977__10
timestamp 1644511149
transform -1 0 40112 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1978__11
timestamp 1644511149
transform 1 0 9200 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1979__12
timestamp 1644511149
transform -1 0 42228 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1980__13
timestamp 1644511149
transform 1 0 4416 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1981__14
timestamp 1644511149
transform -1 0 41032 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1982__15
timestamp 1644511149
transform 1 0 39376 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1983__16
timestamp 1644511149
transform -1 0 40940 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1984__17
timestamp 1644511149
transform -1 0 19872 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1985__18
timestamp 1644511149
transform -1 0 35512 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1986__19
timestamp 1644511149
transform 1 0 4048 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1987__20
timestamp 1644511149
transform -1 0 23644 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1988__21
timestamp 1644511149
transform -1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1989__22
timestamp 1644511149
transform -1 0 42228 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1990__23
timestamp 1644511149
transform 1 0 41584 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1991__24
timestamp 1644511149
transform -1 0 6624 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1992__25
timestamp 1644511149
transform 1 0 39376 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1993__26
timestamp 1644511149
transform 1 0 2576 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1994__27
timestamp 1644511149
transform 1 0 41584 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1995__28
timestamp 1644511149
transform -1 0 27232 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1996__29
timestamp 1644511149
transform -1 0 11776 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1997__30
timestamp 1644511149
transform 1 0 41584 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1998__31
timestamp 1644511149
transform 1 0 2668 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1999__32
timestamp 1644511149
transform 1 0 38456 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2000__33
timestamp 1644511149
transform -1 0 1932 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2001__34
timestamp 1644511149
transform -1 0 38088 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2002__35
timestamp 1644511149
transform -1 0 5336 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2003__36
timestamp 1644511149
transform -1 0 41032 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2004__37
timestamp 1644511149
transform 1 0 39100 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2005__38
timestamp 1644511149
transform -1 0 38732 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2006__39
timestamp 1644511149
transform -1 0 29808 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2007__40
timestamp 1644511149
transform -1 0 6624 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2008__41
timestamp 1644511149
transform 1 0 2576 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2009__42
timestamp 1644511149
transform 1 0 41584 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2010__43
timestamp 1644511149
transform -1 0 20424 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2011__44
timestamp 1644511149
transform 1 0 39100 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2012__45
timestamp 1644511149
transform -1 0 2300 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2013__46
timestamp 1644511149
transform 1 0 15456 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2014__47
timestamp 1644511149
transform -1 0 2300 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2015__48
timestamp 1644511149
transform 1 0 41584 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2016__49
timestamp 1644511149
transform -1 0 2208 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2017__50
timestamp 1644511149
transform 1 0 36340 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2018__51
timestamp 1644511149
transform -1 0 2300 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2019__52
timestamp 1644511149
transform -1 0 28060 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2020__53
timestamp 1644511149
transform 1 0 39376 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2021__54
timestamp 1644511149
transform 1 0 22908 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2022__55
timestamp 1644511149
transform -1 0 32844 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2023__56
timestamp 1644511149
transform -1 0 2300 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2024__57
timestamp 1644511149
transform 1 0 33672 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2025__58
timestamp 1644511149
transform -1 0 15088 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2026__59
timestamp 1644511149
transform 1 0 41584 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2027__60
timestamp 1644511149
transform -1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2028__61
timestamp 1644511149
transform -1 0 1932 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2029__62
timestamp 1644511149
transform -1 0 1932 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2030__63
timestamp 1644511149
transform -1 0 41216 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2031__64
timestamp 1644511149
transform 1 0 41676 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2032__65
timestamp 1644511149
transform -1 0 42228 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2033__66
timestamp 1644511149
transform -1 0 14352 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2034__67
timestamp 1644511149
transform 1 0 39376 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2035__68
timestamp 1644511149
transform 1 0 22264 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2036__69
timestamp 1644511149
transform 1 0 34500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2037__70
timestamp 1644511149
transform -1 0 14996 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2038__71
timestamp 1644511149
transform -1 0 22172 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2039__72
timestamp 1644511149
transform 1 0 40664 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2040__73
timestamp 1644511149
transform -1 0 1932 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2041__74
timestamp 1644511149
transform 1 0 40020 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2042__75
timestamp 1644511149
transform 1 0 10764 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2043__76
timestamp 1644511149
transform -1 0 4508 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2044__77
timestamp 1644511149
transform -1 0 10120 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2045__78
timestamp 1644511149
transform -1 0 2024 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2046__79
timestamp 1644511149
transform -1 0 40756 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2047__80
timestamp 1644511149
transform 1 0 41584 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2048__81
timestamp 1644511149
transform -1 0 41032 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2049__82
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2050__83
timestamp 1644511149
transform 1 0 9660 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2051__84
timestamp 1644511149
transform 1 0 36524 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2052__85
timestamp 1644511149
transform 1 0 10764 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2053__86
timestamp 1644511149
transform 1 0 31372 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2054__87
timestamp 1644511149
transform 1 0 12972 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2055__88
timestamp 1644511149
transform -1 0 40940 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2056__89
timestamp 1644511149
transform -1 0 4048 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2057__90
timestamp 1644511149
transform -1 0 4692 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2058__91
timestamp 1644511149
transform -1 0 22724 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2059__92
timestamp 1644511149
transform 1 0 23092 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2060__93
timestamp 1644511149
transform -1 0 41216 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2061__94
timestamp 1644511149
transform -1 0 40940 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2062__95
timestamp 1644511149
transform 1 0 25852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2063__96
timestamp 1644511149
transform 1 0 36524 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2064__97
timestamp 1644511149
transform 1 0 41584 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2065__98
timestamp 1644511149
transform -1 0 4048 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2066__99
timestamp 1644511149
transform -1 0 35880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2067__100
timestamp 1644511149
transform -1 0 1932 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2068__101
timestamp 1644511149
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2069__102
timestamp 1644511149
transform 1 0 9016 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2070__103
timestamp 1644511149
transform -1 0 1932 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2071__104
timestamp 1644511149
transform -1 0 1932 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2072__105
timestamp 1644511149
transform -1 0 1656 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2073_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7176 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2074_
timestamp 1644511149
transform 1 0 1656 0 -1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2075_
timestamp 1644511149
transform 1 0 18124 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2076_
timestamp 1644511149
transform 1 0 1748 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2077_
timestamp 1644511149
transform 1 0 39836 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2078_
timestamp 1644511149
transform -1 0 11040 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2079_
timestamp 1644511149
transform -1 0 41952 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2080_
timestamp 1644511149
transform -1 0 5612 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2081_
timestamp 1644511149
transform 1 0 40296 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2082_
timestamp 1644511149
transform 1 0 40296 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2083_
timestamp 1644511149
transform 1 0 40296 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2084_
timestamp 1644511149
transform 1 0 19504 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2085_
timestamp 1644511149
transform 1 0 34868 0 -1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2086_
timestamp 1644511149
transform 1 0 4692 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2087_
timestamp 1644511149
transform 1 0 23276 0 -1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2088_
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2089_
timestamp 1644511149
transform -1 0 41952 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2090_
timestamp 1644511149
transform -1 0 42228 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2091_
timestamp 1644511149
transform -1 0 6532 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2092_
timestamp 1644511149
transform 1 0 40296 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2093_
timestamp 1644511149
transform -1 0 3312 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2094_
timestamp 1644511149
transform -1 0 42228 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2095_
timestamp 1644511149
transform 1 0 26956 0 -1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2096_
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2097_
timestamp 1644511149
transform -1 0 42228 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2098_
timestamp 1644511149
transform -1 0 3312 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2099_
timestamp 1644511149
transform 1 0 39560 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2100_
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2101_
timestamp 1644511149
transform 1 0 37536 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2102_
timestamp 1644511149
transform 1 0 4692 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2103_
timestamp 1644511149
transform 1 0 40296 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2104_
timestamp 1644511149
transform 1 0 40020 0 -1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2105_
timestamp 1644511149
transform 1 0 37444 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2106_
timestamp 1644511149
transform 1 0 29532 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2107_
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2108_
timestamp 1644511149
transform -1 0 4508 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2109_
timestamp 1644511149
transform -1 0 41952 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2110_
timestamp 1644511149
transform 1 0 20148 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2111_
timestamp 1644511149
transform 1 0 40020 0 -1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2112_
timestamp 1644511149
transform 1 0 1932 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2113_
timestamp 1644511149
transform 1 0 16100 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2114_
timestamp 1644511149
transform 1 0 1932 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2115_
timestamp 1644511149
transform -1 0 41952 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2116_
timestamp 1644511149
transform 1 0 12144 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2117_
timestamp 1644511149
transform 1 0 11776 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2118_
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2119_
timestamp 1644511149
transform 1 0 40296 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2120_
timestamp 1644511149
transform -1 0 5704 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2121_
timestamp 1644511149
transform 1 0 40020 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2122_
timestamp 1644511149
transform 1 0 40020 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2123_
timestamp 1644511149
transform 1 0 40204 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2124_
timestamp 1644511149
transform 1 0 1840 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2125_
timestamp 1644511149
transform -1 0 37076 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2126_
timestamp 1644511149
transform 1 0 1932 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2127_
timestamp 1644511149
transform 1 0 27784 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2128_
timestamp 1644511149
transform 1 0 40296 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2129_
timestamp 1644511149
transform 1 0 23460 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2130_
timestamp 1644511149
transform 1 0 32292 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2131_
timestamp 1644511149
transform 1 0 1932 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2132_
timestamp 1644511149
transform 1 0 34684 0 -1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2133_
timestamp 1644511149
transform 1 0 14260 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2134_
timestamp 1644511149
transform -1 0 42228 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2135_
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2136_
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2137_
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2138_
timestamp 1644511149
transform 1 0 40296 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2139_
timestamp 1644511149
transform -1 0 42228 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2140_
timestamp 1644511149
transform -1 0 41952 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2141_
timestamp 1644511149
transform 1 0 14076 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2142_
timestamp 1644511149
transform 1 0 40020 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2143_
timestamp 1644511149
transform 1 0 22632 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2144_
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2145_
timestamp 1644511149
transform 1 0 14076 0 -1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2146_
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2147_
timestamp 1644511149
transform -1 0 41952 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2148_
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2149_
timestamp 1644511149
transform 1 0 40296 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2150_
timestamp 1644511149
transform 1 0 10948 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2151_
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2152_
timestamp 1644511149
transform 1 0 9016 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2153_
timestamp 1644511149
transform 1 0 1748 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2154_
timestamp 1644511149
transform 1 0 40020 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2155_
timestamp 1644511149
transform -1 0 42228 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2156_
timestamp 1644511149
transform 1 0 40296 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2157_
timestamp 1644511149
transform -1 0 5060 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2158_
timestamp 1644511149
transform -1 0 13524 0 -1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2159_
timestamp 1644511149
transform 1 0 37444 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2160_
timestamp 1644511149
transform 1 0 11316 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2161_
timestamp 1644511149
transform 1 0 32108 0 -1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2162_
timestamp 1644511149
transform -1 0 13616 0 -1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2163_
timestamp 1644511149
transform 1 0 40020 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2164_
timestamp 1644511149
transform -1 0 3312 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2165_
timestamp 1644511149
transform 1 0 3956 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2166_
timestamp 1644511149
transform 1 0 21804 0 -1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2167_
timestamp 1644511149
transform 1 0 24380 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2168_
timestamp 1644511149
transform 1 0 40296 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2169_
timestamp 1644511149
transform 1 0 40020 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2170_
timestamp 1644511149
transform 1 0 26680 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2171_
timestamp 1644511149
transform 1 0 36984 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2172_
timestamp 1644511149
transform -1 0 42228 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2173_
timestamp 1644511149
transform 1 0 3772 0 -1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2174_
timestamp 1644511149
transform 1 0 34868 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2175_
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2176_
timestamp 1644511149
transform 1 0 38456 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2177_
timestamp 1644511149
transform 1 0 9108 0 -1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2178_
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2179_
timestamp 1644511149
transform 1 0 1656 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2180_
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i
timestamp 1644511149
transform -1 0 28244 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_0_0_wb_clk_i
timestamp 1644511149
transform -1 0 20976 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_1_0_wb_clk_i
timestamp 1644511149
transform -1 0 20516 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_2_0_wb_clk_i
timestamp 1644511149
transform -1 0 27876 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 29900 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_4_0_wb_clk_i
timestamp 1644511149
transform 1 0 21528 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_5_0_wb_clk_i
timestamp 1644511149
transform -1 0 22816 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_6_0_wb_clk_i
timestamp 1644511149
transform 1 0 31280 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_7_0_wb_clk_i
timestamp 1644511149
transform 1 0 31556 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_0_0_wb_clk_i
timestamp 1644511149
transform -1 0 19964 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_2_0_wb_clk_i
timestamp 1644511149
transform -1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 21620 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_4_0_wb_clk_i
timestamp 1644511149
transform -1 0 26496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_5_0_wb_clk_i
timestamp 1644511149
transform 1 0 31188 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_6_0_wb_clk_i
timestamp 1644511149
transform -1 0 28336 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_7_0_wb_clk_i
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_8_0_wb_clk_i
timestamp 1644511149
transform -1 0 19780 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_9_0_wb_clk_i
timestamp 1644511149
transform 1 0 22724 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_10_0_wb_clk_i
timestamp 1644511149
transform -1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_11_0_wb_clk_i
timestamp 1644511149
transform 1 0 22908 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_12_0_wb_clk_i
timestamp 1644511149
transform -1 0 30544 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_13_0_wb_clk_i
timestamp 1644511149
transform 1 0 33212 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_14_0_wb_clk_i
timestamp 1644511149
transform -1 0 30360 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_15_0_wb_clk_i
timestamp 1644511149
transform 1 0 33304 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24840 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2
timestamp 1644511149
transform 1 0 28336 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1644511149
transform -1 0 26404 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  input1
timestamp 1644511149
transform 1 0 1748 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1644511149
transform 1 0 24748 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input3
timestamp 1644511149
transform -1 0 42228 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1644511149
transform 1 0 7820 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 1644511149
transform -1 0 41952 0 -1 7616
box -38 -48 406 592
<< labels >>
rlabel metal3 s 0 40808 800 40928 6 active
port 0 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 24490 43200 24546 44000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 18 43200 74 44000 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 43200 36728 44000 36848 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 16762 43200 16818 44000 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 43200 38768 44000 38888 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 43200 3408 44000 3528 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 9034 43200 9090 44000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 10966 43200 11022 44000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 io_in[20]
port 13 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 io_in[21]
port 14 nsew signal input
rlabel metal3 s 43200 13608 44000 13728 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 8390 43200 8446 44000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 5814 43200 5870 44000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 43200 9528 44000 9648 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 43810 43200 43866 44000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 43200 17008 44000 17128 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 39448 800 39568 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 33506 43200 33562 44000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 38658 43200 38714 44000 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 43200 27208 44000 27328 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 39302 43200 39358 44000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 25134 43200 25190 44000 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 43200 26528 44000 26648 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 43200 42168 44000 42288 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 43200 29248 44000 29368 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 7746 43200 7802 44000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 io_oeb[0]
port 39 nsew signal tristate
rlabel metal3 s 0 14968 800 15088 6 io_oeb[10]
port 40 nsew signal tristate
rlabel metal3 s 43200 25168 44000 25288 6 io_oeb[11]
port 41 nsew signal tristate
rlabel metal3 s 43200 12928 44000 13048 6 io_oeb[12]
port 42 nsew signal tristate
rlabel metal3 s 43200 12248 44000 12368 6 io_oeb[13]
port 43 nsew signal tristate
rlabel metal3 s 0 4088 800 4208 6 io_oeb[14]
port 44 nsew signal tristate
rlabel metal2 s 12254 43200 12310 44000 6 io_oeb[15]
port 45 nsew signal tristate
rlabel metal3 s 43200 2048 44000 2168 6 io_oeb[16]
port 46 nsew signal tristate
rlabel metal2 s 11610 0 11666 800 6 io_oeb[17]
port 47 nsew signal tristate
rlabel metal2 s 32218 43200 32274 44000 6 io_oeb[18]
port 48 nsew signal tristate
rlabel metal2 s 12898 43200 12954 44000 6 io_oeb[19]
port 49 nsew signal tristate
rlabel metal2 s 34794 0 34850 800 6 io_oeb[1]
port 50 nsew signal tristate
rlabel metal3 s 43200 19048 44000 19168 6 io_oeb[20]
port 51 nsew signal tristate
rlabel metal2 s 1950 43200 2006 44000 6 io_oeb[21]
port 52 nsew signal tristate
rlabel metal2 s 4526 0 4582 800 6 io_oeb[22]
port 53 nsew signal tristate
rlabel metal2 s 21914 43200 21970 44000 6 io_oeb[23]
port 54 nsew signal tristate
rlabel metal2 s 23202 43200 23258 44000 6 io_oeb[24]
port 55 nsew signal tristate
rlabel metal2 s 41878 0 41934 800 6 io_oeb[25]
port 56 nsew signal tristate
rlabel metal3 s 43200 34688 44000 34808 6 io_oeb[26]
port 57 nsew signal tristate
rlabel metal2 s 26422 43200 26478 44000 6 io_oeb[27]
port 58 nsew signal tristate
rlabel metal2 s 37370 0 37426 800 6 io_oeb[28]
port 59 nsew signal tristate
rlabel metal3 s 43200 28568 44000 28688 6 io_oeb[29]
port 60 nsew signal tristate
rlabel metal2 s 36726 43200 36782 44000 6 io_oeb[2]
port 61 nsew signal tristate
rlabel metal2 s 2594 43200 2650 44000 6 io_oeb[30]
port 62 nsew signal tristate
rlabel metal2 s 36082 0 36138 800 6 io_oeb[31]
port 63 nsew signal tristate
rlabel metal3 s 0 21768 800 21888 6 io_oeb[32]
port 64 nsew signal tristate
rlabel metal2 s 43166 0 43222 800 6 io_oeb[33]
port 65 nsew signal tristate
rlabel metal2 s 9678 43200 9734 44000 6 io_oeb[34]
port 66 nsew signal tristate
rlabel metal3 s 0 19728 800 19848 6 io_oeb[35]
port 67 nsew signal tristate
rlabel metal3 s 0 10208 800 10328 6 io_oeb[36]
port 68 nsew signal tristate
rlabel metal3 s 0 16328 800 16448 6 io_oeb[37]
port 69 nsew signal tristate
rlabel metal2 s 22558 0 22614 800 6 io_oeb[3]
port 70 nsew signal tristate
rlabel metal3 s 43200 8 44000 128 6 io_oeb[4]
port 71 nsew signal tristate
rlabel metal3 s 0 28568 800 28688 6 io_oeb[5]
port 72 nsew signal tristate
rlabel metal3 s 43200 15648 44000 15768 6 io_oeb[6]
port 73 nsew signal tristate
rlabel metal2 s 11610 43200 11666 44000 6 io_oeb[7]
port 74 nsew signal tristate
rlabel metal2 s 3882 0 3938 800 6 io_oeb[8]
port 75 nsew signal tristate
rlabel metal2 s 9678 0 9734 800 6 io_oeb[9]
port 76 nsew signal tristate
rlabel metal3 s 43200 41488 44000 41608 6 io_out[0]
port 77 nsew signal tristate
rlabel metal3 s 43200 23808 44000 23928 6 io_out[10]
port 78 nsew signal tristate
rlabel metal3 s 0 2048 800 2168 6 io_out[11]
port 79 nsew signal tristate
rlabel metal3 s 0 6808 800 6928 6 io_out[12]
port 80 nsew signal tristate
rlabel metal2 s 35438 0 35494 800 6 io_out[13]
port 81 nsew signal tristate
rlabel metal3 s 43200 35368 44000 35488 6 io_out[14]
port 82 nsew signal tristate
rlabel metal3 s 0 36728 800 36848 6 io_out[15]
port 83 nsew signal tristate
rlabel metal3 s 43200 23128 44000 23248 6 io_out[16]
port 84 nsew signal tristate
rlabel metal2 s 40590 43200 40646 44000 6 io_out[17]
port 85 nsew signal tristate
rlabel metal2 s 41234 0 41290 800 6 io_out[18]
port 86 nsew signal tristate
rlabel metal3 s 0 21088 800 21208 6 io_out[19]
port 87 nsew signal tristate
rlabel metal2 s 29642 43200 29698 44000 6 io_out[1]
port 88 nsew signal tristate
rlabel metal2 s 36082 43200 36138 44000 6 io_out[20]
port 89 nsew signal tristate
rlabel metal3 s 0 36048 800 36168 6 io_out[21]
port 90 nsew signal tristate
rlabel metal2 s 28354 0 28410 800 6 io_out[22]
port 91 nsew signal tristate
rlabel metal3 s 43200 19728 44000 19848 6 io_out[23]
port 92 nsew signal tristate
rlabel metal2 s 23846 0 23902 800 6 io_out[24]
port 93 nsew signal tristate
rlabel metal2 s 32862 43200 32918 44000 6 io_out[25]
port 94 nsew signal tristate
rlabel metal3 s 0 4768 800 4888 6 io_out[26]
port 95 nsew signal tristate
rlabel metal2 s 34150 43200 34206 44000 6 io_out[27]
port 96 nsew signal tristate
rlabel metal2 s 15474 0 15530 800 6 io_out[28]
port 97 nsew signal tristate
rlabel metal3 s 43200 688 44000 808 6 io_out[29]
port 98 nsew signal tristate
rlabel metal2 s 6458 0 6514 800 6 io_out[2]
port 99 nsew signal tristate
rlabel metal3 s 0 5448 800 5568 6 io_out[30]
port 100 nsew signal tristate
rlabel metal3 s 0 12248 800 12368 6 io_out[31]
port 101 nsew signal tristate
rlabel metal3 s 0 41488 800 41608 6 io_out[32]
port 102 nsew signal tristate
rlabel metal3 s 43200 6128 44000 6248 6 io_out[33]
port 103 nsew signal tristate
rlabel metal3 s 43200 36048 44000 36168 6 io_out[34]
port 104 nsew signal tristate
rlabel metal3 s 43200 33328 44000 33448 6 io_out[35]
port 105 nsew signal tristate
rlabel metal2 s 14186 43200 14242 44000 6 io_out[36]
port 106 nsew signal tristate
rlabel metal3 s 43200 39448 44000 39568 6 io_out[37]
port 107 nsew signal tristate
rlabel metal3 s 0 38088 800 38208 6 io_out[3]
port 108 nsew signal tristate
rlabel metal3 s 43200 25848 44000 25968 6 io_out[4]
port 109 nsew signal tristate
rlabel metal2 s 20626 43200 20682 44000 6 io_out[5]
port 110 nsew signal tristate
rlabel metal2 s 42522 43200 42578 44000 6 io_out[6]
port 111 nsew signal tristate
rlabel metal3 s 0 17688 800 17808 6 io_out[7]
port 112 nsew signal tristate
rlabel metal2 s 16762 0 16818 800 6 io_out[8]
port 113 nsew signal tristate
rlabel metal3 s 0 13608 800 13728 6 io_out[9]
port 114 nsew signal tristate
rlabel metal3 s 43200 6808 44000 6928 6 la1_data_in[0]
port 115 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 la1_data_in[10]
port 116 nsew signal input
rlabel metal3 s 43200 5448 44000 5568 6 la1_data_in[11]
port 117 nsew signal input
rlabel metal3 s 0 33328 800 33448 6 la1_data_in[12]
port 118 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 la1_data_in[13]
port 119 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 la1_data_in[14]
port 120 nsew signal input
rlabel metal2 s 14830 43200 14886 44000 6 la1_data_in[15]
port 121 nsew signal input
rlabel metal2 s 27710 43200 27766 44000 6 la1_data_in[16]
port 122 nsew signal input
rlabel metal2 s 21270 43200 21326 44000 6 la1_data_in[17]
port 123 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 la1_data_in[18]
port 124 nsew signal input
rlabel metal2 s 15474 43200 15530 44000 6 la1_data_in[19]
port 125 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 la1_data_in[1]
port 126 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 la1_data_in[20]
port 127 nsew signal input
rlabel metal2 s 43166 43200 43222 44000 6 la1_data_in[21]
port 128 nsew signal input
rlabel metal3 s 43200 7488 44000 7608 6 la1_data_in[22]
port 129 nsew signal input
rlabel metal3 s 0 688 800 808 6 la1_data_in[23]
port 130 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 la1_data_in[24]
port 131 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 la1_data_in[25]
port 132 nsew signal input
rlabel metal3 s 43200 2728 44000 2848 6 la1_data_in[26]
port 133 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 la1_data_in[27]
port 134 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 la1_data_in[28]
port 135 nsew signal input
rlabel metal2 s 662 43200 718 44000 6 la1_data_in[29]
port 136 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 la1_data_in[2]
port 137 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 la1_data_in[30]
port 138 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 la1_data_in[31]
port 139 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 la1_data_in[3]
port 140 nsew signal input
rlabel metal2 s 37370 43200 37426 44000 6 la1_data_in[4]
port 141 nsew signal input
rlabel metal3 s 43200 21768 44000 21888 6 la1_data_in[5]
port 142 nsew signal input
rlabel metal2 s 17406 43200 17462 44000 6 la1_data_in[6]
port 143 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 la1_data_in[7]
port 144 nsew signal input
rlabel metal2 s 18050 43200 18106 44000 6 la1_data_in[8]
port 145 nsew signal input
rlabel metal3 s 0 30608 800 30728 6 la1_data_in[9]
port 146 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 la1_data_out[0]
port 147 nsew signal tristate
rlabel metal3 s 43200 10208 44000 10328 6 la1_data_out[10]
port 148 nsew signal tristate
rlabel metal2 s 19982 0 20038 800 6 la1_data_out[11]
port 149 nsew signal tristate
rlabel metal3 s 43200 40128 44000 40248 6 la1_data_out[12]
port 150 nsew signal tristate
rlabel metal2 s 4526 43200 4582 44000 6 la1_data_out[13]
port 151 nsew signal tristate
rlabel metal2 s 23846 43200 23902 44000 6 la1_data_out[14]
port 152 nsew signal tristate
rlabel metal3 s 0 1368 800 1488 6 la1_data_out[15]
port 153 nsew signal tristate
rlabel metal3 s 43200 14968 44000 15088 6 la1_data_out[16]
port 154 nsew signal tristate
rlabel metal3 s 43200 31968 44000 32088 6 la1_data_out[17]
port 155 nsew signal tristate
rlabel metal2 s 5170 43200 5226 44000 6 la1_data_out[18]
port 156 nsew signal tristate
rlabel metal3 s 43200 22448 44000 22568 6 la1_data_out[19]
port 157 nsew signal tristate
rlabel metal3 s 0 40128 800 40248 6 la1_data_out[1]
port 158 nsew signal tristate
rlabel metal3 s 0 8848 800 8968 6 la1_data_out[20]
port 159 nsew signal tristate
rlabel metal3 s 43200 38088 44000 38208 6 la1_data_out[21]
port 160 nsew signal tristate
rlabel metal2 s 27066 43200 27122 44000 6 la1_data_out[22]
port 161 nsew signal tristate
rlabel metal2 s 10966 0 11022 800 6 la1_data_out[23]
port 162 nsew signal tristate
rlabel metal3 s 43200 16328 44000 16448 6 la1_data_out[24]
port 163 nsew signal tristate
rlabel metal3 s 0 3408 800 3528 6 la1_data_out[25]
port 164 nsew signal tristate
rlabel metal3 s 43200 4088 44000 4208 6 la1_data_out[26]
port 165 nsew signal tristate
rlabel metal3 s 0 42848 800 42968 6 la1_data_out[27]
port 166 nsew signal tristate
rlabel metal2 s 39302 0 39358 800 6 la1_data_out[28]
port 167 nsew signal tristate
rlabel metal2 s 5170 0 5226 800 6 la1_data_out[29]
port 168 nsew signal tristate
rlabel metal2 s 18694 0 18750 800 6 la1_data_out[2]
port 169 nsew signal tristate
rlabel metal3 s 43200 10888 44000 11008 6 la1_data_out[30]
port 170 nsew signal tristate
rlabel metal3 s 43200 42848 44000 42968 6 la1_data_out[31]
port 171 nsew signal tristate
rlabel metal3 s 0 8168 800 8288 6 la1_data_out[3]
port 172 nsew signal tristate
rlabel metal2 s 40590 0 40646 800 6 la1_data_out[4]
port 173 nsew signal tristate
rlabel metal2 s 3238 0 3294 800 6 la1_data_out[5]
port 174 nsew signal tristate
rlabel metal3 s 43200 18368 44000 18488 6 la1_data_out[6]
port 175 nsew signal tristate
rlabel metal2 s 662 0 718 800 6 la1_data_out[7]
port 176 nsew signal tristate
rlabel metal3 s 43200 32648 44000 32768 6 la1_data_out[8]
port 177 nsew signal tristate
rlabel metal2 s 41878 43200 41934 44000 6 la1_data_out[9]
port 178 nsew signal tristate
rlabel metal2 s 43810 0 43866 800 6 la1_oenb[0]
port 179 nsew signal input
rlabel metal2 s 39946 43200 40002 44000 6 la1_oenb[10]
port 180 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 la1_oenb[11]
port 181 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 la1_oenb[12]
port 182 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 la1_oenb[13]
port 183 nsew signal input
rlabel metal2 s 18 0 74 800 6 la1_oenb[14]
port 184 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 la1_oenb[15]
port 185 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 la1_oenb[16]
port 186 nsew signal input
rlabel metal2 s 3238 43200 3294 44000 6 la1_oenb[17]
port 187 nsew signal input
rlabel metal2 s 19982 43200 20038 44000 6 la1_oenb[18]
port 188 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 la1_oenb[19]
port 189 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 la1_oenb[1]
port 190 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 la1_oenb[20]
port 191 nsew signal input
rlabel metal2 s 28354 43200 28410 44000 6 la1_oenb[21]
port 192 nsew signal input
rlabel metal2 s 18694 43200 18750 44000 6 la1_oenb[22]
port 193 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 la1_oenb[23]
port 194 nsew signal input
rlabel metal2 s 35438 43200 35494 44000 6 la1_oenb[24]
port 195 nsew signal input
rlabel metal3 s 43200 8848 44000 8968 6 la1_oenb[25]
port 196 nsew signal input
rlabel metal3 s 0 34688 800 34808 6 la1_oenb[26]
port 197 nsew signal input
rlabel metal3 s 43200 31288 44000 31408 6 la1_oenb[27]
port 198 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 la1_oenb[28]
port 199 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 la1_oenb[29]
port 200 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 la1_oenb[2]
port 201 nsew signal input
rlabel metal3 s 43200 29928 44000 30048 6 la1_oenb[30]
port 202 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 la1_oenb[31]
port 203 nsew signal input
rlabel metal2 s 30930 43200 30986 44000 6 la1_oenb[3]
port 204 nsew signal input
rlabel metal2 s 30286 43200 30342 44000 6 la1_oenb[4]
port 205 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 la1_oenb[5]
port 206 nsew signal input
rlabel metal2 s 6458 43200 6514 44000 6 la1_oenb[6]
port 207 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 la1_oenb[7]
port 208 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 la1_oenb[8]
port 209 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 la1_oenb[9]
port 210 nsew signal input
rlabel metal4 s 4208 2128 4528 41392 6 vccd1
port 211 nsew power input
rlabel metal4 s 34928 2128 35248 41392 6 vccd1
port 211 nsew power input
rlabel metal4 s 19568 2128 19888 41392 6 vssd1
port 212 nsew ground input
rlabel metal3 s 43200 20408 44000 20528 6 wb_clk_i
port 213 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 44000 44000
<< end >>
