magic
tech sky130A
magscale 1 2
timestamp 1647517048
<< obsli1 >>
rect 1104 2159 44896 43537
<< obsm1 >>
rect 658 2128 45158 44124
<< metal2 >>
rect -10 45200 102 46000
rect 634 45200 746 46000
rect 1922 45200 2034 46000
rect 2566 45200 2678 46000
rect 3210 45200 3322 46000
rect 4498 45200 4610 46000
rect 5142 45200 5254 46000
rect 5786 45200 5898 46000
rect 7074 45200 7186 46000
rect 7718 45200 7830 46000
rect 8362 45200 8474 46000
rect 9650 45200 9762 46000
rect 10294 45200 10406 46000
rect 10938 45200 11050 46000
rect 12226 45200 12338 46000
rect 12870 45200 12982 46000
rect 13514 45200 13626 46000
rect 14802 45200 14914 46000
rect 15446 45200 15558 46000
rect 16090 45200 16202 46000
rect 17378 45200 17490 46000
rect 18022 45200 18134 46000
rect 18666 45200 18778 46000
rect 19954 45200 20066 46000
rect 20598 45200 20710 46000
rect 21242 45200 21354 46000
rect 22530 45200 22642 46000
rect 23174 45200 23286 46000
rect 23818 45200 23930 46000
rect 24462 45200 24574 46000
rect 25750 45200 25862 46000
rect 26394 45200 26506 46000
rect 27038 45200 27150 46000
rect 28326 45200 28438 46000
rect 28970 45200 29082 46000
rect 29614 45200 29726 46000
rect 30902 45200 31014 46000
rect 31546 45200 31658 46000
rect 32190 45200 32302 46000
rect 33478 45200 33590 46000
rect 34122 45200 34234 46000
rect 34766 45200 34878 46000
rect 36054 45200 36166 46000
rect 36698 45200 36810 46000
rect 37342 45200 37454 46000
rect 38630 45200 38742 46000
rect 39274 45200 39386 46000
rect 39918 45200 40030 46000
rect 41206 45200 41318 46000
rect 41850 45200 41962 46000
rect 42494 45200 42606 46000
rect 43782 45200 43894 46000
rect 44426 45200 44538 46000
rect 45070 45200 45182 46000
rect 45714 45200 45826 46000
rect -10 0 102 800
rect 634 0 746 800
rect 1278 0 1390 800
rect 1922 0 2034 800
rect 3210 0 3322 800
rect 3854 0 3966 800
rect 4498 0 4610 800
rect 5786 0 5898 800
rect 6430 0 6542 800
rect 7074 0 7186 800
rect 8362 0 8474 800
rect 9006 0 9118 800
rect 9650 0 9762 800
rect 10938 0 11050 800
rect 11582 0 11694 800
rect 12226 0 12338 800
rect 13514 0 13626 800
rect 14158 0 14270 800
rect 14802 0 14914 800
rect 16090 0 16202 800
rect 16734 0 16846 800
rect 17378 0 17490 800
rect 18666 0 18778 800
rect 19310 0 19422 800
rect 19954 0 20066 800
rect 21242 0 21354 800
rect 21886 0 21998 800
rect 22530 0 22642 800
rect 23174 0 23286 800
rect 24462 0 24574 800
rect 25106 0 25218 800
rect 25750 0 25862 800
rect 27038 0 27150 800
rect 27682 0 27794 800
rect 28326 0 28438 800
rect 29614 0 29726 800
rect 30258 0 30370 800
rect 30902 0 31014 800
rect 32190 0 32302 800
rect 32834 0 32946 800
rect 33478 0 33590 800
rect 34766 0 34878 800
rect 35410 0 35522 800
rect 36054 0 36166 800
rect 37342 0 37454 800
rect 37986 0 38098 800
rect 38630 0 38742 800
rect 39918 0 40030 800
rect 40562 0 40674 800
rect 41206 0 41318 800
rect 42494 0 42606 800
rect 43138 0 43250 800
rect 43782 0 43894 800
rect 45070 0 45182 800
rect 45714 0 45826 800
<< obsm2 >>
rect 802 45144 1866 45200
rect 2090 45144 2510 45200
rect 2734 45144 3154 45200
rect 3378 45144 4442 45200
rect 4666 45144 5086 45200
rect 5310 45144 5730 45200
rect 5954 45144 7018 45200
rect 7242 45144 7662 45200
rect 7886 45144 8306 45200
rect 8530 45144 9594 45200
rect 9818 45144 10238 45200
rect 10462 45144 10882 45200
rect 11106 45144 12170 45200
rect 12394 45144 12814 45200
rect 13038 45144 13458 45200
rect 13682 45144 14746 45200
rect 14970 45144 15390 45200
rect 15614 45144 16034 45200
rect 16258 45144 17322 45200
rect 17546 45144 17966 45200
rect 18190 45144 18610 45200
rect 18834 45144 19898 45200
rect 20122 45144 20542 45200
rect 20766 45144 21186 45200
rect 21410 45144 22474 45200
rect 22698 45144 23118 45200
rect 23342 45144 23762 45200
rect 23986 45144 24406 45200
rect 24630 45144 25694 45200
rect 25918 45144 26338 45200
rect 26562 45144 26982 45200
rect 27206 45144 28270 45200
rect 28494 45144 28914 45200
rect 29138 45144 29558 45200
rect 29782 45144 30846 45200
rect 31070 45144 31490 45200
rect 31714 45144 32134 45200
rect 32358 45144 33422 45200
rect 33646 45144 34066 45200
rect 34290 45144 34710 45200
rect 34934 45144 35998 45200
rect 36222 45144 36642 45200
rect 36866 45144 37286 45200
rect 37510 45144 38574 45200
rect 38798 45144 39218 45200
rect 39442 45144 39862 45200
rect 40086 45144 41150 45200
rect 41374 45144 41794 45200
rect 42018 45144 42438 45200
rect 42662 45144 43726 45200
rect 43950 45144 44370 45200
rect 44594 45144 45014 45200
rect 664 856 45152 45144
rect 802 31 1222 856
rect 1446 31 1866 856
rect 2090 31 3154 856
rect 3378 31 3798 856
rect 4022 31 4442 856
rect 4666 31 5730 856
rect 5954 31 6374 856
rect 6598 31 7018 856
rect 7242 31 8306 856
rect 8530 31 8950 856
rect 9174 31 9594 856
rect 9818 31 10882 856
rect 11106 31 11526 856
rect 11750 31 12170 856
rect 12394 31 13458 856
rect 13682 31 14102 856
rect 14326 31 14746 856
rect 14970 31 16034 856
rect 16258 31 16678 856
rect 16902 31 17322 856
rect 17546 31 18610 856
rect 18834 31 19254 856
rect 19478 31 19898 856
rect 20122 31 21186 856
rect 21410 31 21830 856
rect 22054 31 22474 856
rect 22698 31 23118 856
rect 23342 31 24406 856
rect 24630 31 25050 856
rect 25274 31 25694 856
rect 25918 31 26982 856
rect 27206 31 27626 856
rect 27850 31 28270 856
rect 28494 31 29558 856
rect 29782 31 30202 856
rect 30426 31 30846 856
rect 31070 31 32134 856
rect 32358 31 32778 856
rect 33002 31 33422 856
rect 33646 31 34710 856
rect 34934 31 35354 856
rect 35578 31 35998 856
rect 36222 31 37286 856
rect 37510 31 37930 856
rect 38154 31 38574 856
rect 38798 31 39862 856
rect 40086 31 40506 856
rect 40730 31 41150 856
rect 41374 31 42438 856
rect 42662 31 43082 856
rect 43306 31 43726 856
rect 43950 31 45014 856
<< metal3 >>
rect 0 45508 800 45748
rect 0 44828 800 45068
rect 45200 44828 46000 45068
rect 45200 44148 46000 44388
rect 0 43468 800 43708
rect 45200 43468 46000 43708
rect 0 42788 800 43028
rect 0 42108 800 42348
rect 45200 42108 46000 42348
rect 45200 41428 46000 41668
rect 0 40748 800 40988
rect 45200 40748 46000 40988
rect 0 40068 800 40308
rect 0 39388 800 39628
rect 45200 39388 46000 39628
rect 45200 38708 46000 38948
rect 0 38028 800 38268
rect 45200 38028 46000 38268
rect 0 37348 800 37588
rect 0 36668 800 36908
rect 45200 36668 46000 36908
rect 45200 35988 46000 36228
rect 0 35308 800 35548
rect 45200 35308 46000 35548
rect 0 34628 800 34868
rect 0 33948 800 34188
rect 45200 33948 46000 34188
rect 45200 33268 46000 33508
rect 0 32588 800 32828
rect 45200 32588 46000 32828
rect 0 31908 800 32148
rect 0 31228 800 31468
rect 45200 31228 46000 31468
rect 45200 30548 46000 30788
rect 0 29868 800 30108
rect 45200 29868 46000 30108
rect 0 29188 800 29428
rect 0 28508 800 28748
rect 45200 28508 46000 28748
rect 45200 27828 46000 28068
rect 0 27148 800 27388
rect 45200 27148 46000 27388
rect 0 26468 800 26708
rect 0 25788 800 26028
rect 45200 25788 46000 26028
rect 45200 25108 46000 25348
rect 0 24428 800 24668
rect 45200 24428 46000 24668
rect 0 23748 800 23988
rect 0 23068 800 23308
rect 45200 23068 46000 23308
rect 0 22388 800 22628
rect 45200 22388 46000 22628
rect 45200 21708 46000 21948
rect 0 21028 800 21268
rect 45200 21028 46000 21268
rect 0 20348 800 20588
rect 0 19668 800 19908
rect 45200 19668 46000 19908
rect 45200 18988 46000 19228
rect 0 18308 800 18548
rect 45200 18308 46000 18548
rect 0 17628 800 17868
rect 0 16948 800 17188
rect 45200 16948 46000 17188
rect 45200 16268 46000 16508
rect 0 15588 800 15828
rect 45200 15588 46000 15828
rect 0 14908 800 15148
rect 0 14228 800 14468
rect 45200 14228 46000 14468
rect 45200 13548 46000 13788
rect 0 12868 800 13108
rect 45200 12868 46000 13108
rect 0 12188 800 12428
rect 0 11508 800 11748
rect 45200 11508 46000 11748
rect 45200 10828 46000 11068
rect 0 10148 800 10388
rect 45200 10148 46000 10388
rect 0 9468 800 9708
rect 0 8788 800 9028
rect 45200 8788 46000 9028
rect 45200 8108 46000 8348
rect 0 7428 800 7668
rect 45200 7428 46000 7668
rect 0 6748 800 6988
rect 0 6068 800 6308
rect 45200 6068 46000 6308
rect 45200 5388 46000 5628
rect 0 4708 800 4948
rect 45200 4708 46000 4948
rect 0 4028 800 4268
rect 0 3348 800 3588
rect 45200 3348 46000 3588
rect 45200 2668 46000 2908
rect 0 1988 800 2228
rect 45200 1988 46000 2228
rect 0 1308 800 1548
rect 0 628 800 868
rect 45200 628 46000 868
rect 45200 -52 46000 188
<< obsm3 >>
rect 880 44748 45120 44981
rect 800 44468 45200 44748
rect 800 44068 45120 44468
rect 800 43788 45200 44068
rect 880 43388 45120 43788
rect 800 43108 45200 43388
rect 880 42708 45200 43108
rect 800 42428 45200 42708
rect 880 42028 45120 42428
rect 800 41748 45200 42028
rect 800 41348 45120 41748
rect 800 41068 45200 41348
rect 880 40668 45120 41068
rect 800 40388 45200 40668
rect 880 39988 45200 40388
rect 800 39708 45200 39988
rect 880 39308 45120 39708
rect 800 39028 45200 39308
rect 800 38628 45120 39028
rect 800 38348 45200 38628
rect 880 37948 45120 38348
rect 800 37668 45200 37948
rect 880 37268 45200 37668
rect 800 36988 45200 37268
rect 880 36588 45120 36988
rect 800 36308 45200 36588
rect 800 35908 45120 36308
rect 800 35628 45200 35908
rect 880 35228 45120 35628
rect 800 34948 45200 35228
rect 880 34548 45200 34948
rect 800 34268 45200 34548
rect 880 33868 45120 34268
rect 800 33588 45200 33868
rect 800 33188 45120 33588
rect 800 32908 45200 33188
rect 880 32508 45120 32908
rect 800 32228 45200 32508
rect 880 31828 45200 32228
rect 800 31548 45200 31828
rect 880 31148 45120 31548
rect 800 30868 45200 31148
rect 800 30468 45120 30868
rect 800 30188 45200 30468
rect 880 29788 45120 30188
rect 800 29508 45200 29788
rect 880 29108 45200 29508
rect 800 28828 45200 29108
rect 880 28428 45120 28828
rect 800 28148 45200 28428
rect 800 27748 45120 28148
rect 800 27468 45200 27748
rect 880 27068 45120 27468
rect 800 26788 45200 27068
rect 880 26388 45200 26788
rect 800 26108 45200 26388
rect 880 25708 45120 26108
rect 800 25428 45200 25708
rect 800 25028 45120 25428
rect 800 24748 45200 25028
rect 880 24348 45120 24748
rect 800 24068 45200 24348
rect 880 23668 45200 24068
rect 800 23388 45200 23668
rect 880 22988 45120 23388
rect 800 22708 45200 22988
rect 880 22308 45120 22708
rect 800 22028 45200 22308
rect 800 21628 45120 22028
rect 800 21348 45200 21628
rect 880 20948 45120 21348
rect 800 20668 45200 20948
rect 880 20268 45200 20668
rect 800 19988 45200 20268
rect 880 19588 45120 19988
rect 800 19308 45200 19588
rect 800 18908 45120 19308
rect 800 18628 45200 18908
rect 880 18228 45120 18628
rect 800 17948 45200 18228
rect 880 17548 45200 17948
rect 800 17268 45200 17548
rect 880 16868 45120 17268
rect 800 16588 45200 16868
rect 800 16188 45120 16588
rect 800 15908 45200 16188
rect 880 15508 45120 15908
rect 800 15228 45200 15508
rect 880 14828 45200 15228
rect 800 14548 45200 14828
rect 880 14148 45120 14548
rect 800 13868 45200 14148
rect 800 13468 45120 13868
rect 800 13188 45200 13468
rect 880 12788 45120 13188
rect 800 12508 45200 12788
rect 880 12108 45200 12508
rect 800 11828 45200 12108
rect 880 11428 45120 11828
rect 800 11148 45200 11428
rect 800 10748 45120 11148
rect 800 10468 45200 10748
rect 880 10068 45120 10468
rect 800 9788 45200 10068
rect 880 9388 45200 9788
rect 800 9108 45200 9388
rect 880 8708 45120 9108
rect 800 8428 45200 8708
rect 800 8028 45120 8428
rect 800 7748 45200 8028
rect 880 7348 45120 7748
rect 800 7068 45200 7348
rect 880 6668 45200 7068
rect 800 6388 45200 6668
rect 880 5988 45120 6388
rect 800 5708 45200 5988
rect 800 5308 45120 5708
rect 800 5028 45200 5308
rect 880 4628 45120 5028
rect 800 4348 45200 4628
rect 880 3948 45200 4348
rect 800 3668 45200 3948
rect 880 3268 45120 3668
rect 800 2988 45200 3268
rect 800 2588 45120 2988
rect 800 2308 45200 2588
rect 880 1908 45120 2308
rect 800 1628 45200 1908
rect 880 1228 45200 1628
rect 800 948 45200 1228
rect 880 548 45120 948
rect 800 268 45200 548
rect 800 35 45120 268
<< metal4 >>
rect 4208 2128 4528 43568
rect 19568 2128 19888 43568
rect 34928 2128 35248 43568
<< obsm4 >>
rect 24899 3979 34848 35597
rect 35328 3979 43181 35597
<< labels >>
rlabel metal3 s 0 42788 800 43028 6 active
port 1 nsew signal input
rlabel metal2 s 14158 0 14270 800 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 25750 45200 25862 46000 6 io_in[10]
port 3 nsew signal input
rlabel metal2 s -10 45200 102 46000 6 io_in[11]
port 4 nsew signal input
rlabel metal3 s 45200 38708 46000 38948 6 io_in[12]
port 5 nsew signal input
rlabel metal2 s 21886 0 21998 800 6 io_in[13]
port 6 nsew signal input
rlabel metal2 s 17378 45200 17490 46000 6 io_in[14]
port 7 nsew signal input
rlabel metal3 s 45200 40748 46000 40988 6 io_in[15]
port 8 nsew signal input
rlabel metal3 s 45200 3348 46000 3588 6 io_in[16]
port 9 nsew signal input
rlabel metal2 s 9650 45200 9762 46000 6 io_in[17]
port 10 nsew signal input
rlabel metal2 s 10938 45200 11050 46000 6 io_in[18]
port 11 nsew signal input
rlabel metal2 s 39918 0 40030 800 6 io_in[19]
port 12 nsew signal input
rlabel metal3 s 0 14908 800 15148 6 io_in[1]
port 13 nsew signal input
rlabel metal3 s 0 26468 800 26708 6 io_in[20]
port 14 nsew signal input
rlabel metal3 s 0 17628 800 17868 6 io_in[21]
port 15 nsew signal input
rlabel metal3 s 45200 14228 46000 14468 6 io_in[22]
port 16 nsew signal input
rlabel metal2 s 8362 45200 8474 46000 6 io_in[23]
port 17 nsew signal input
rlabel metal2 s 5786 45200 5898 46000 6 io_in[24]
port 18 nsew signal input
rlabel metal2 s 34766 0 34878 800 6 io_in[25]
port 19 nsew signal input
rlabel metal2 s 33478 0 33590 800 6 io_in[26]
port 20 nsew signal input
rlabel metal3 s 45200 10148 46000 10388 6 io_in[27]
port 21 nsew signal input
rlabel metal2 s 30258 0 30370 800 6 io_in[28]
port 22 nsew signal input
rlabel metal2 s 45714 45200 45826 46000 6 io_in[29]
port 23 nsew signal input
rlabel metal2 s 14802 0 14914 800 6 io_in[2]
port 24 nsew signal input
rlabel metal3 s 45200 18308 46000 18548 6 io_in[30]
port 25 nsew signal input
rlabel metal3 s 0 40748 800 40988 6 io_in[31]
port 26 nsew signal input
rlabel metal2 s 28326 0 28438 800 6 io_in[32]
port 27 nsew signal input
rlabel metal3 s 0 23748 800 23988 6 io_in[33]
port 28 nsew signal input
rlabel metal2 s 34766 45200 34878 46000 6 io_in[34]
port 29 nsew signal input
rlabel metal2 s 39918 45200 40030 46000 6 io_in[35]
port 30 nsew signal input
rlabel metal3 s 45200 28508 46000 28748 6 io_in[36]
port 31 nsew signal input
rlabel metal2 s 41206 45200 41318 46000 6 io_in[37]
port 32 nsew signal input
rlabel metal2 s 26394 45200 26506 46000 6 io_in[3]
port 33 nsew signal input
rlabel metal3 s 45200 27828 46000 28068 6 io_in[4]
port 34 nsew signal input
rlabel metal3 s 45200 44148 46000 44388 6 io_in[5]
port 35 nsew signal input
rlabel metal3 s 0 28508 800 28748 6 io_in[6]
port 36 nsew signal input
rlabel metal3 s 0 19668 800 19908 6 io_in[7]
port 37 nsew signal input
rlabel metal3 s 45200 30548 46000 30788 6 io_in[8]
port 38 nsew signal input
rlabel metal2 s 7718 45200 7830 46000 6 io_in[9]
port 39 nsew signal input
rlabel metal2 s 24462 0 24574 800 6 io_oeb[0]
port 40 nsew signal output
rlabel metal3 s 0 15588 800 15828 6 io_oeb[10]
port 41 nsew signal output
rlabel metal3 s 45200 25788 46000 26028 6 io_oeb[11]
port 42 nsew signal output
rlabel metal3 s 45200 13548 46000 13788 6 io_oeb[12]
port 43 nsew signal output
rlabel metal3 s 45200 12868 46000 13108 6 io_oeb[13]
port 44 nsew signal output
rlabel metal3 s 0 4028 800 4268 6 io_oeb[14]
port 45 nsew signal output
rlabel metal2 s 12870 45200 12982 46000 6 io_oeb[15]
port 46 nsew signal output
rlabel metal3 s 45200 1988 46000 2228 6 io_oeb[16]
port 47 nsew signal output
rlabel metal2 s 12226 0 12338 800 6 io_oeb[17]
port 48 nsew signal output
rlabel metal2 s 33478 45200 33590 46000 6 io_oeb[18]
port 49 nsew signal output
rlabel metal2 s 13514 45200 13626 46000 6 io_oeb[19]
port 50 nsew signal output
rlabel metal2 s 36054 0 36166 800 6 io_oeb[1]
port 51 nsew signal output
rlabel metal3 s 45200 19668 46000 19908 6 io_oeb[20]
port 52 nsew signal output
rlabel metal2 s 1922 45200 2034 46000 6 io_oeb[21]
port 53 nsew signal output
rlabel metal2 s 4498 0 4610 800 6 io_oeb[22]
port 54 nsew signal output
rlabel metal2 s 23174 45200 23286 46000 6 io_oeb[23]
port 55 nsew signal output
rlabel metal2 s 23818 45200 23930 46000 6 io_oeb[24]
port 56 nsew signal output
rlabel metal2 s 43782 0 43894 800 6 io_oeb[25]
port 57 nsew signal output
rlabel metal3 s 45200 35988 46000 36228 6 io_oeb[26]
port 58 nsew signal output
rlabel metal2 s 27038 45200 27150 46000 6 io_oeb[27]
port 59 nsew signal output
rlabel metal2 s 38630 0 38742 800 6 io_oeb[28]
port 60 nsew signal output
rlabel metal3 s 45200 29868 46000 30108 6 io_oeb[29]
port 61 nsew signal output
rlabel metal2 s 38630 45200 38742 46000 6 io_oeb[2]
port 62 nsew signal output
rlabel metal2 s 2566 45200 2678 46000 6 io_oeb[30]
port 63 nsew signal output
rlabel metal2 s 37986 0 38098 800 6 io_oeb[31]
port 64 nsew signal output
rlabel metal3 s 0 23068 800 23308 6 io_oeb[32]
port 65 nsew signal output
rlabel metal2 s 45070 0 45182 800 6 io_oeb[33]
port 66 nsew signal output
rlabel metal2 s 10294 45200 10406 46000 6 io_oeb[34]
port 67 nsew signal output
rlabel metal3 s 0 20348 800 20588 6 io_oeb[35]
port 68 nsew signal output
rlabel metal3 s 0 10148 800 10388 6 io_oeb[36]
port 69 nsew signal output
rlabel metal3 s 0 16948 800 17188 6 io_oeb[37]
port 70 nsew signal output
rlabel metal2 s 23174 0 23286 800 6 io_oeb[3]
port 71 nsew signal output
rlabel metal3 s 45200 -52 46000 188 6 io_oeb[4]
port 72 nsew signal output
rlabel metal3 s 0 29868 800 30108 6 io_oeb[5]
port 73 nsew signal output
rlabel metal3 s 45200 16268 46000 16508 6 io_oeb[6]
port 74 nsew signal output
rlabel metal2 s 12226 45200 12338 46000 6 io_oeb[7]
port 75 nsew signal output
rlabel metal2 s 3854 0 3966 800 6 io_oeb[8]
port 76 nsew signal output
rlabel metal2 s 9650 0 9762 800 6 io_oeb[9]
port 77 nsew signal output
rlabel metal3 s 45200 43468 46000 43708 6 io_out[0]
port 78 nsew signal output
rlabel metal3 s 45200 25108 46000 25348 6 io_out[10]
port 79 nsew signal output
rlabel metal3 s 0 1988 800 2228 6 io_out[11]
port 80 nsew signal output
rlabel metal3 s 0 6748 800 6988 6 io_out[12]
port 81 nsew signal output
rlabel metal2 s 37342 0 37454 800 6 io_out[13]
port 82 nsew signal output
rlabel metal3 s 45200 36668 46000 36908 6 io_out[14]
port 83 nsew signal output
rlabel metal3 s 0 38028 800 38268 6 io_out[15]
port 84 nsew signal output
rlabel metal3 s 45200 24428 46000 24668 6 io_out[16]
port 85 nsew signal output
rlabel metal2 s 42494 45200 42606 46000 6 io_out[17]
port 86 nsew signal output
rlabel metal2 s 43138 0 43250 800 6 io_out[18]
port 87 nsew signal output
rlabel metal3 s 0 22388 800 22628 6 io_out[19]
port 88 nsew signal output
rlabel metal2 s 30902 45200 31014 46000 6 io_out[1]
port 89 nsew signal output
rlabel metal2 s 37342 45200 37454 46000 6 io_out[20]
port 90 nsew signal output
rlabel metal3 s 0 37348 800 37588 6 io_out[21]
port 91 nsew signal output
rlabel metal2 s 29614 0 29726 800 6 io_out[22]
port 92 nsew signal output
rlabel metal3 s 45200 21028 46000 21268 6 io_out[23]
port 93 nsew signal output
rlabel metal2 s 25106 0 25218 800 6 io_out[24]
port 94 nsew signal output
rlabel metal2 s 34122 45200 34234 46000 6 io_out[25]
port 95 nsew signal output
rlabel metal3 s 0 4708 800 4948 6 io_out[26]
port 96 nsew signal output
rlabel metal2 s 36054 45200 36166 46000 6 io_out[27]
port 97 nsew signal output
rlabel metal2 s 16090 0 16202 800 6 io_out[28]
port 98 nsew signal output
rlabel metal3 s 45200 628 46000 868 6 io_out[29]
port 99 nsew signal output
rlabel metal2 s 6430 0 6542 800 6 io_out[2]
port 100 nsew signal output
rlabel metal3 s 0 6068 800 6308 6 io_out[30]
port 101 nsew signal output
rlabel metal3 s 0 12868 800 13108 6 io_out[31]
port 102 nsew signal output
rlabel metal3 s 0 43468 800 43708 6 io_out[32]
port 103 nsew signal output
rlabel metal3 s 45200 6068 46000 6308 6 io_out[33]
port 104 nsew signal output
rlabel metal3 s 45200 38028 46000 38268 6 io_out[34]
port 105 nsew signal output
rlabel metal3 s 45200 35308 46000 35548 6 io_out[35]
port 106 nsew signal output
rlabel metal2 s 14802 45200 14914 46000 6 io_out[36]
port 107 nsew signal output
rlabel metal3 s 45200 41428 46000 41668 6 io_out[37]
port 108 nsew signal output
rlabel metal3 s 0 40068 800 40308 6 io_out[3]
port 109 nsew signal output
rlabel metal3 s 45200 27148 46000 27388 6 io_out[4]
port 110 nsew signal output
rlabel metal2 s 21242 45200 21354 46000 6 io_out[5]
port 111 nsew signal output
rlabel metal2 s 44426 45200 44538 46000 6 io_out[6]
port 112 nsew signal output
rlabel metal3 s 0 18308 800 18548 6 io_out[7]
port 113 nsew signal output
rlabel metal2 s 17378 0 17490 800 6 io_out[8]
port 114 nsew signal output
rlabel metal3 s 0 14228 800 14468 6 io_out[9]
port 115 nsew signal output
rlabel metal3 s 45200 7428 46000 7668 6 la1_data_in[0]
port 116 nsew signal input
rlabel metal2 s 19954 0 20066 800 6 la1_data_in[10]
port 117 nsew signal input
rlabel metal3 s 45200 5388 46000 5628 6 la1_data_in[11]
port 118 nsew signal input
rlabel metal3 s 0 34628 800 34868 6 la1_data_in[12]
port 119 nsew signal input
rlabel metal2 s 30902 0 31014 800 6 la1_data_in[13]
port 120 nsew signal input
rlabel metal3 s 0 12188 800 12428 6 la1_data_in[14]
port 121 nsew signal input
rlabel metal2 s 15446 45200 15558 46000 6 la1_data_in[15]
port 122 nsew signal input
rlabel metal2 s 28970 45200 29082 46000 6 la1_data_in[16]
port 123 nsew signal input
rlabel metal2 s 22530 45200 22642 46000 6 la1_data_in[17]
port 124 nsew signal input
rlabel metal2 s 40562 0 40674 800 6 la1_data_in[18]
port 125 nsew signal input
rlabel metal2 s 16090 45200 16202 46000 6 la1_data_in[19]
port 126 nsew signal input
rlabel metal2 s 18666 0 18778 800 6 la1_data_in[1]
port 127 nsew signal input
rlabel metal3 s 0 33948 800 34188 6 la1_data_in[20]
port 128 nsew signal input
rlabel metal2 s 45070 45200 45182 46000 6 la1_data_in[21]
port 129 nsew signal input
rlabel metal3 s 45200 8108 46000 8348 6 la1_data_in[22]
port 130 nsew signal input
rlabel metal3 s 0 628 800 868 6 la1_data_in[23]
port 131 nsew signal input
rlabel metal2 s 13514 0 13626 800 6 la1_data_in[24]
port 132 nsew signal input
rlabel metal3 s 0 35308 800 35548 6 la1_data_in[25]
port 133 nsew signal input
rlabel metal3 s 45200 2668 46000 2908 6 la1_data_in[26]
port 134 nsew signal input
rlabel metal2 s 27038 0 27150 800 6 la1_data_in[27]
port 135 nsew signal input
rlabel metal3 s 0 31228 800 31468 6 la1_data_in[28]
port 136 nsew signal input
rlabel metal2 s 634 45200 746 46000 6 la1_data_in[29]
port 137 nsew signal input
rlabel metal2 s 10938 0 11050 800 6 la1_data_in[2]
port 138 nsew signal input
rlabel metal2 s 1278 0 1390 800 6 la1_data_in[30]
port 139 nsew signal input
rlabel metal2 s 35410 0 35522 800 6 la1_data_in[31]
port 140 nsew signal input
rlabel metal3 s 0 29188 800 29428 6 la1_data_in[3]
port 141 nsew signal input
rlabel metal2 s 39274 45200 39386 46000 6 la1_data_in[4]
port 142 nsew signal input
rlabel metal3 s 45200 22388 46000 22628 6 la1_data_in[5]
port 143 nsew signal input
rlabel metal2 s 18022 45200 18134 46000 6 la1_data_in[6]
port 144 nsew signal input
rlabel metal3 s 0 21028 800 21268 6 la1_data_in[7]
port 145 nsew signal input
rlabel metal2 s 18666 45200 18778 46000 6 la1_data_in[8]
port 146 nsew signal input
rlabel metal3 s 0 31908 800 32148 6 la1_data_in[9]
port 147 nsew signal input
rlabel metal2 s 7074 0 7186 800 6 la1_data_out[0]
port 148 nsew signal output
rlabel metal3 s 45200 10828 46000 11068 6 la1_data_out[10]
port 149 nsew signal output
rlabel metal2 s 21242 0 21354 800 6 la1_data_out[11]
port 150 nsew signal output
rlabel metal3 s 45200 42108 46000 42348 6 la1_data_out[12]
port 151 nsew signal output
rlabel metal2 s 4498 45200 4610 46000 6 la1_data_out[13]
port 152 nsew signal output
rlabel metal2 s 24462 45200 24574 46000 6 la1_data_out[14]
port 153 nsew signal output
rlabel metal3 s 0 1308 800 1548 6 la1_data_out[15]
port 154 nsew signal output
rlabel metal3 s 45200 15588 46000 15828 6 la1_data_out[16]
port 155 nsew signal output
rlabel metal3 s 45200 33268 46000 33508 6 la1_data_out[17]
port 156 nsew signal output
rlabel metal2 s 5142 45200 5254 46000 6 la1_data_out[18]
port 157 nsew signal output
rlabel metal3 s 45200 23068 46000 23308 6 la1_data_out[19]
port 158 nsew signal output
rlabel metal3 s 0 42108 800 42348 6 la1_data_out[1]
port 159 nsew signal output
rlabel metal3 s 0 9468 800 9708 6 la1_data_out[20]
port 160 nsew signal output
rlabel metal3 s 45200 39388 46000 39628 6 la1_data_out[21]
port 161 nsew signal output
rlabel metal2 s 28326 45200 28438 46000 6 la1_data_out[22]
port 162 nsew signal output
rlabel metal2 s 11582 0 11694 800 6 la1_data_out[23]
port 163 nsew signal output
rlabel metal3 s 45200 16948 46000 17188 6 la1_data_out[24]
port 164 nsew signal output
rlabel metal3 s 0 3348 800 3588 6 la1_data_out[25]
port 165 nsew signal output
rlabel metal3 s 45200 4708 46000 4948 6 la1_data_out[26]
port 166 nsew signal output
rlabel metal3 s 0 44828 800 45068 6 la1_data_out[27]
port 167 nsew signal output
rlabel metal2 s 41206 0 41318 800 6 la1_data_out[28]
port 168 nsew signal output
rlabel metal2 s 5786 0 5898 800 6 la1_data_out[29]
port 169 nsew signal output
rlabel metal2 s 19310 0 19422 800 6 la1_data_out[2]
port 170 nsew signal output
rlabel metal3 s 45200 11508 46000 11748 6 la1_data_out[30]
port 171 nsew signal output
rlabel metal3 s 45200 44828 46000 45068 6 la1_data_out[31]
port 172 nsew signal output
rlabel metal3 s 0 8788 800 9028 6 la1_data_out[3]
port 173 nsew signal output
rlabel metal2 s 42494 0 42606 800 6 la1_data_out[4]
port 174 nsew signal output
rlabel metal2 s 3210 0 3322 800 6 la1_data_out[5]
port 175 nsew signal output
rlabel metal3 s 45200 18988 46000 19228 6 la1_data_out[6]
port 176 nsew signal output
rlabel metal2 s 634 0 746 800 6 la1_data_out[7]
port 177 nsew signal output
rlabel metal3 s 45200 33948 46000 34188 6 la1_data_out[8]
port 178 nsew signal output
rlabel metal2 s 43782 45200 43894 46000 6 la1_data_out[9]
port 179 nsew signal output
rlabel metal2 s 45714 0 45826 800 6 la1_oenb[0]
port 180 nsew signal input
rlabel metal2 s 41850 45200 41962 46000 6 la1_oenb[10]
port 181 nsew signal input
rlabel metal3 s 0 25788 800 26028 6 la1_oenb[11]
port 182 nsew signal input
rlabel metal3 s 0 27148 800 27388 6 la1_oenb[12]
port 183 nsew signal input
rlabel metal2 s 27682 0 27794 800 6 la1_oenb[13]
port 184 nsew signal input
rlabel metal2 s -10 0 102 800 6 la1_oenb[14]
port 185 nsew signal input
rlabel metal2 s 32834 0 32946 800 6 la1_oenb[15]
port 186 nsew signal input
rlabel metal3 s 0 32588 800 32828 6 la1_oenb[16]
port 187 nsew signal input
rlabel metal2 s 3210 45200 3322 46000 6 la1_oenb[17]
port 188 nsew signal input
rlabel metal2 s 20598 45200 20710 46000 6 la1_oenb[18]
port 189 nsew signal input
rlabel metal3 s 0 24428 800 24668 6 la1_oenb[19]
port 190 nsew signal input
rlabel metal2 s 8362 0 8474 800 6 la1_oenb[1]
port 191 nsew signal input
rlabel metal2 s 1922 0 2034 800 6 la1_oenb[20]
port 192 nsew signal input
rlabel metal2 s 29614 45200 29726 46000 6 la1_oenb[21]
port 193 nsew signal input
rlabel metal2 s 19954 45200 20066 46000 6 la1_oenb[22]
port 194 nsew signal input
rlabel metal2 s 22530 0 22642 800 6 la1_oenb[23]
port 195 nsew signal input
rlabel metal2 s 36698 45200 36810 46000 6 la1_oenb[24]
port 196 nsew signal input
rlabel metal3 s 45200 8788 46000 9028 6 la1_oenb[25]
port 197 nsew signal input
rlabel metal3 s 0 36668 800 36908 6 la1_oenb[26]
port 198 nsew signal input
rlabel metal3 s 45200 32588 46000 32828 6 la1_oenb[27]
port 199 nsew signal input
rlabel metal2 s 9006 0 9118 800 6 la1_oenb[28]
port 200 nsew signal input
rlabel metal2 s 16734 0 16846 800 6 la1_oenb[29]
port 201 nsew signal input
rlabel metal3 s 0 7428 800 7668 6 la1_oenb[2]
port 202 nsew signal input
rlabel metal3 s 45200 31228 46000 31468 6 la1_oenb[30]
port 203 nsew signal input
rlabel metal2 s 25750 0 25862 800 6 la1_oenb[31]
port 204 nsew signal input
rlabel metal2 s 32190 45200 32302 46000 6 la1_oenb[3]
port 205 nsew signal input
rlabel metal2 s 31546 45200 31658 46000 6 la1_oenb[4]
port 206 nsew signal input
rlabel metal3 s 0 45508 800 45748 6 la1_oenb[5]
port 207 nsew signal input
rlabel metal2 s 7074 45200 7186 46000 6 la1_oenb[6]
port 208 nsew signal input
rlabel metal2 s 32190 0 32302 800 6 la1_oenb[7]
port 209 nsew signal input
rlabel metal3 s 0 11508 800 11748 6 la1_oenb[8]
port 210 nsew signal input
rlabel metal3 s 0 39388 800 39628 6 la1_oenb[9]
port 211 nsew signal input
rlabel metal4 s 4208 2128 4528 43568 6 vccd1
port 212 nsew power input
rlabel metal4 s 34928 2128 35248 43568 6 vccd1
port 212 nsew power input
rlabel metal4 s 19568 2128 19888 43568 6 vssd1
port 213 nsew ground input
rlabel metal3 s 45200 21708 46000 21948 6 wb_clk_i
port 214 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 46000 46000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3335800
string GDS_FILE /openlane/designs/wrapped_vga_clock/runs/RUN_2022.03.17_11.36.08/results/finishing/wrapped_vga_clock.magic.gds
string GDS_START 519986
<< end >>

