magic
tech sky130A
magscale 1 2
timestamp 1647517046
<< viali >>
rect 13185 43333 13219 43367
rect 14289 43333 14323 43367
rect 24593 43333 24627 43367
rect 27537 43333 27571 43367
rect 1869 43265 1903 43299
rect 2881 43265 2915 43299
rect 7849 43265 7883 43299
rect 12541 43265 12575 43299
rect 13093 43265 13127 43299
rect 2145 43197 2179 43231
rect 3801 43197 3835 43231
rect 3985 43197 4019 43231
rect 4261 43197 4295 43231
rect 14105 43197 14139 43231
rect 14565 43197 14599 43231
rect 23489 43197 23523 43231
rect 24409 43197 24443 43231
rect 24869 43197 24903 43231
rect 32321 43197 32355 43231
rect 32505 43197 32539 43231
rect 33517 43197 33551 43231
rect 2789 43061 2823 43095
rect 6561 43061 6595 43095
rect 8033 43061 8067 43095
rect 10977 43061 11011 43095
rect 11713 43061 11747 43095
rect 12449 43061 12483 43095
rect 20821 43061 20855 43095
rect 22661 43061 22695 43095
rect 27445 43061 27479 43095
rect 28089 43061 28123 43095
rect 30481 43061 30515 43095
rect 40049 43061 40083 43095
rect 42901 43061 42935 43095
rect 43821 43061 43855 43095
rect 2789 42721 2823 42755
rect 4353 42721 4387 42755
rect 6653 42721 6687 42755
rect 10333 42721 10367 42755
rect 11621 42721 11655 42755
rect 12449 42721 12483 42755
rect 14841 42721 14875 42755
rect 20821 42721 20855 42755
rect 21281 42721 21315 42755
rect 24869 42721 24903 42755
rect 27169 42721 27203 42755
rect 30481 42721 30515 42755
rect 30941 42721 30975 42755
rect 33149 42721 33183 42755
rect 37381 42721 37415 42755
rect 39957 42721 39991 42755
rect 41797 42721 41831 42755
rect 42349 42721 42383 42755
rect 43821 42721 43855 42755
rect 3249 42653 3283 42687
rect 4813 42653 4847 42687
rect 7113 42653 7147 42687
rect 9321 42653 9355 42687
rect 14381 42653 14415 42687
rect 16681 42653 16715 42687
rect 23857 42653 23891 42687
rect 24409 42653 24443 42687
rect 26709 42653 26743 42687
rect 33977 42653 34011 42687
rect 35449 42653 35483 42687
rect 36277 42653 36311 42687
rect 36737 42653 36771 42687
rect 3065 42585 3099 42619
rect 6469 42585 6503 42619
rect 9505 42585 9539 42619
rect 11805 42585 11839 42619
rect 14565 42585 14599 42619
rect 21005 42585 21039 42619
rect 24593 42585 24627 42619
rect 26893 42585 26927 42619
rect 30665 42585 30699 42619
rect 36921 42585 36955 42619
rect 40141 42585 40175 42619
rect 42533 42585 42567 42619
rect 10885 42313 10919 42347
rect 20913 42313 20947 42347
rect 27077 42313 27111 42347
rect 30665 42313 30699 42347
rect 33333 42313 33367 42347
rect 42717 42313 42751 42347
rect 2053 42245 2087 42279
rect 5457 42245 5491 42279
rect 6561 42245 6595 42279
rect 12173 42245 12207 42279
rect 16129 42245 16163 42279
rect 37473 42245 37507 42279
rect 38301 42245 38335 42279
rect 39957 42245 39991 42279
rect 4721 42177 4755 42211
rect 5549 42177 5583 42211
rect 9873 42177 9907 42211
rect 10793 42177 10827 42211
rect 11989 42177 12023 42211
rect 14289 42177 14323 42211
rect 20821 42177 20855 42211
rect 22661 42177 22695 42211
rect 26433 42177 26467 42211
rect 27169 42177 27203 42211
rect 27813 42177 27847 42211
rect 30573 42177 30607 42211
rect 33425 42177 33459 42211
rect 33977 42177 34011 42211
rect 36461 42177 36495 42211
rect 37381 42177 37415 42211
rect 42809 42177 42843 42211
rect 43453 42177 43487 42211
rect 43913 42177 43947 42211
rect 1869 42109 1903 42143
rect 2881 42109 2915 42143
rect 6377 42109 6411 42143
rect 7757 42109 7791 42143
rect 12909 42109 12943 42143
rect 14473 42109 14507 42143
rect 22845 42109 22879 42143
rect 23213 42109 23247 42143
rect 27997 42109 28031 42143
rect 28365 42109 28399 42143
rect 34161 42109 34195 42143
rect 34897 42109 34931 42143
rect 38117 42109 38151 42143
rect 4813 41973 4847 42007
rect 36369 41973 36403 42007
rect 43361 41973 43395 42007
rect 44005 41973 44039 42007
rect 3893 41769 3927 41803
rect 10057 41769 10091 41803
rect 14565 41769 14599 41803
rect 22753 41769 22787 41803
rect 23397 41769 23431 41803
rect 24501 41769 24535 41803
rect 28089 41769 28123 41803
rect 34805 41769 34839 41803
rect 37841 41769 37875 41803
rect 38393 41769 38427 41803
rect 39957 41769 39991 41803
rect 15117 41701 15151 41735
rect 2789 41633 2823 41667
rect 3249 41633 3283 41667
rect 5181 41633 5215 41667
rect 6377 41633 6411 41667
rect 6561 41633 6595 41667
rect 35449 41633 35483 41667
rect 35633 41633 35667 41667
rect 36093 41633 36127 41667
rect 42533 41633 42567 41667
rect 44005 41633 44039 41667
rect 44189 41633 44223 41667
rect 3985 41565 4019 41599
rect 10149 41565 10183 41599
rect 11529 41565 11563 41599
rect 12081 41565 12115 41599
rect 14473 41565 14507 41599
rect 22661 41565 22695 41599
rect 23305 41565 23339 41599
rect 24409 41565 24443 41599
rect 28181 41565 28215 41599
rect 34897 41565 34931 41599
rect 37933 41565 37967 41599
rect 39865 41565 39899 41599
rect 3065 41497 3099 41531
rect 10977 41497 11011 41531
rect 12909 41497 12943 41531
rect 2973 41225 3007 41259
rect 6469 41225 6503 41259
rect 14197 41225 14231 41259
rect 2329 41157 2363 41191
rect 41705 41157 41739 41191
rect 43453 41157 43487 41191
rect 1777 41089 1811 41123
rect 2421 41089 2455 41123
rect 3065 41089 3099 41123
rect 3525 41089 3559 41123
rect 5457 41089 5491 41123
rect 6561 41089 6595 41123
rect 9045 41089 9079 41123
rect 10701 41089 10735 41123
rect 11897 41089 11931 41123
rect 14105 41089 14139 41123
rect 32505 41089 32539 41123
rect 32597 41089 32631 41123
rect 32781 41089 32815 41123
rect 33425 41089 33459 41123
rect 43361 41089 43395 41123
rect 4721 41021 4755 41055
rect 9597 41021 9631 41055
rect 41337 41021 41371 41055
rect 41889 41021 41923 41055
rect 42717 41021 42751 41055
rect 10885 40953 10919 40987
rect 13369 40885 13403 40919
rect 32965 40885 32999 40919
rect 33609 40885 33643 40919
rect 44189 40885 44223 40919
rect 2881 40681 2915 40715
rect 13461 40681 13495 40715
rect 32321 40681 32355 40715
rect 37289 40613 37323 40647
rect 40785 40613 40819 40647
rect 12173 40545 12207 40579
rect 27445 40545 27479 40579
rect 43269 40545 43303 40579
rect 44005 40545 44039 40579
rect 44189 40545 44223 40579
rect 2053 40477 2087 40511
rect 3893 40477 3927 40511
rect 4629 40477 4663 40511
rect 6929 40477 6963 40511
rect 9321 40477 9355 40511
rect 11989 40477 12023 40511
rect 27629 40477 27663 40511
rect 31125 40477 31159 40511
rect 32137 40477 32171 40511
rect 34161 40477 34195 40511
rect 35081 40477 35115 40511
rect 37013 40477 37047 40511
rect 39313 40477 39347 40511
rect 40049 40477 40083 40511
rect 40509 40477 40543 40511
rect 7481 40409 7515 40443
rect 10149 40409 10183 40443
rect 33894 40409 33928 40443
rect 37289 40409 37323 40443
rect 39068 40409 39102 40443
rect 40785 40409 40819 40443
rect 4077 40341 4111 40375
rect 5917 40341 5951 40375
rect 27813 40341 27847 40375
rect 30941 40341 30975 40375
rect 32781 40341 32815 40375
rect 35265 40341 35299 40375
rect 37105 40341 37139 40375
rect 37933 40341 37967 40375
rect 39865 40341 39899 40375
rect 40601 40341 40635 40375
rect 28365 40137 28399 40171
rect 31125 40137 31159 40171
rect 33517 40137 33551 40171
rect 38669 40137 38703 40171
rect 2145 40069 2179 40103
rect 29837 40069 29871 40103
rect 30053 40069 30087 40103
rect 32137 40069 32171 40103
rect 32353 40069 32387 40103
rect 33333 40069 33367 40103
rect 35642 40069 35676 40103
rect 39497 40069 39531 40103
rect 40754 40069 40788 40103
rect 1961 40001 1995 40035
rect 4721 40001 4755 40035
rect 11989 40001 12023 40035
rect 18972 40001 19006 40035
rect 20545 40001 20579 40035
rect 24308 40001 24342 40035
rect 27241 40001 27275 40035
rect 30665 40001 30699 40035
rect 37545 40001 37579 40035
rect 2789 39933 2823 39967
rect 4905 39933 4939 39967
rect 12173 39933 12207 39967
rect 18705 39933 18739 39967
rect 24041 39933 24075 39967
rect 26985 39933 27019 39967
rect 35909 39933 35943 39967
rect 37289 39933 37323 39967
rect 40509 39933 40543 39967
rect 31033 39865 31067 39899
rect 32505 39865 32539 39899
rect 32965 39865 32999 39899
rect 39129 39865 39163 39899
rect 39681 39865 39715 39899
rect 20085 39797 20119 39831
rect 20729 39797 20763 39831
rect 25421 39797 25455 39831
rect 30021 39797 30055 39831
rect 30205 39797 30239 39831
rect 32321 39797 32355 39831
rect 33333 39797 33367 39831
rect 34529 39797 34563 39831
rect 39497 39797 39531 39831
rect 41889 39797 41923 39831
rect 43821 39797 43855 39831
rect 2881 39593 2915 39627
rect 3801 39593 3835 39627
rect 19257 39593 19291 39627
rect 24593 39593 24627 39627
rect 27077 39593 27111 39627
rect 28917 39593 28951 39627
rect 32137 39593 32171 39627
rect 34161 39593 34195 39627
rect 35081 39593 35115 39627
rect 35265 39593 35299 39627
rect 37381 39593 37415 39627
rect 38945 39593 38979 39627
rect 39129 39593 39163 39627
rect 39865 39593 39899 39627
rect 40877 39593 40911 39627
rect 32689 39525 32723 39559
rect 40969 39525 41003 39559
rect 20453 39457 20487 39491
rect 25973 39457 26007 39491
rect 26433 39457 26467 39491
rect 26801 39457 26835 39491
rect 30757 39457 30791 39491
rect 37289 39457 37323 39491
rect 37473 39457 37507 39491
rect 40785 39457 40819 39491
rect 42717 39457 42751 39491
rect 44189 39457 44223 39491
rect 2973 39389 3007 39423
rect 4813 39389 4847 39423
rect 5641 39389 5675 39423
rect 19441 39389 19475 39423
rect 19533 39389 19567 39423
rect 24409 39389 24443 39423
rect 24685 39389 24719 39423
rect 25513 39389 25547 39423
rect 25605 39389 25639 39423
rect 25789 39389 25823 39423
rect 26893 39389 26927 39423
rect 27537 39389 27571 39423
rect 30297 39389 30331 39423
rect 31024 39389 31058 39423
rect 32873 39389 32907 39423
rect 33793 39389 33827 39423
rect 33977 39389 34011 39423
rect 34713 39389 34747 39423
rect 37565 39389 37599 39423
rect 40049 39389 40083 39423
rect 40325 39389 40359 39423
rect 41061 39389 41095 39423
rect 41705 39389 41739 39423
rect 20720 39321 20754 39355
rect 24501 39321 24535 39355
rect 27804 39321 27838 39355
rect 30113 39321 30147 39355
rect 39113 39321 39147 39355
rect 39313 39321 39347 39355
rect 40233 39321 40267 39355
rect 44005 39321 44039 39355
rect 19901 39253 19935 39287
rect 21833 39253 21867 39287
rect 29929 39253 29963 39287
rect 32965 39253 32999 39287
rect 33057 39253 33091 39287
rect 33241 39253 33275 39287
rect 35081 39253 35115 39287
rect 41521 39253 41555 39287
rect 20361 39049 20395 39083
rect 24685 39049 24719 39083
rect 26341 39049 26375 39083
rect 27905 39049 27939 39083
rect 30849 39049 30883 39083
rect 31309 39049 31343 39083
rect 43453 39049 43487 39083
rect 26985 38981 27019 39015
rect 32873 38981 32907 39015
rect 39773 38981 39807 39015
rect 16865 38913 16899 38947
rect 16957 38913 16991 38947
rect 17141 38913 17175 38947
rect 19073 38913 19107 38947
rect 19349 38913 19383 38947
rect 19533 38913 19567 38947
rect 20177 38913 20211 38947
rect 22192 38913 22226 38947
rect 24409 38913 24443 38947
rect 25145 38913 25179 38947
rect 25329 38913 25363 38947
rect 25513 38913 25547 38947
rect 25973 38913 26007 38947
rect 27169 38913 27203 38947
rect 28089 38913 28123 38947
rect 29469 38913 29503 38947
rect 29736 38913 29770 38947
rect 31309 38913 31343 38947
rect 31493 38913 31527 38947
rect 33149 38913 33183 38947
rect 33333 38913 33367 38947
rect 34069 38913 34103 38947
rect 36737 38913 36771 38947
rect 37473 38913 37507 38947
rect 37657 38913 37691 38947
rect 37749 38913 37783 38947
rect 38853 38913 38887 38947
rect 38945 38913 38979 38947
rect 39589 38913 39623 38947
rect 39865 38913 39899 38947
rect 39957 38913 39991 38947
rect 43361 38913 43395 38947
rect 19993 38845 20027 38879
rect 21925 38845 21959 38879
rect 24685 38845 24719 38879
rect 26065 38845 26099 38879
rect 27445 38845 27479 38879
rect 39129 38845 39163 38879
rect 40785 38845 40819 38879
rect 41061 38845 41095 38879
rect 23305 38777 23339 38811
rect 27353 38777 27387 38811
rect 40141 38777 40175 38811
rect 16865 38709 16899 38743
rect 19165 38709 19199 38743
rect 24501 38709 24535 38743
rect 25973 38709 26007 38743
rect 33057 38709 33091 38743
rect 33517 38709 33551 38743
rect 34253 38709 34287 38743
rect 36553 38709 36587 38743
rect 37289 38709 37323 38743
rect 39037 38709 39071 38743
rect 44189 38709 44223 38743
rect 19349 38505 19383 38539
rect 22201 38505 22235 38539
rect 29929 38505 29963 38539
rect 34989 38437 35023 38471
rect 19717 38369 19751 38403
rect 21649 38369 21683 38403
rect 33333 38369 33367 38403
rect 36093 38369 36127 38403
rect 38485 38369 38519 38403
rect 38577 38369 38611 38403
rect 40509 38369 40543 38403
rect 42717 38369 42751 38403
rect 44189 38369 44223 38403
rect 16313 38301 16347 38335
rect 16580 38301 16614 38335
rect 19533 38301 19567 38335
rect 19809 38301 19843 38335
rect 22109 38301 22143 38335
rect 22293 38301 22327 38335
rect 22845 38301 22879 38335
rect 25605 38301 25639 38335
rect 25881 38301 25915 38335
rect 26525 38301 26559 38335
rect 30113 38301 30147 38335
rect 33609 38301 33643 38335
rect 34713 38301 34747 38335
rect 34989 38301 35023 38335
rect 36360 38301 36394 38335
rect 38209 38301 38243 38335
rect 39865 38301 39899 38335
rect 40049 38301 40083 38335
rect 21382 38233 21416 38267
rect 38694 38233 38728 38267
rect 40776 38233 40810 38267
rect 44005 38233 44039 38267
rect 17693 38165 17727 38199
rect 20269 38165 20303 38199
rect 23029 38165 23063 38199
rect 25421 38165 25455 38199
rect 25789 38165 25823 38199
rect 26617 38165 26651 38199
rect 34805 38165 34839 38199
rect 37473 38165 37507 38199
rect 38853 38165 38887 38199
rect 39957 38165 39991 38199
rect 41889 38165 41923 38199
rect 17325 37961 17359 37995
rect 18429 37961 18463 37995
rect 20545 37961 20579 37995
rect 21281 37961 21315 37995
rect 33425 37961 33459 37995
rect 34253 37961 34287 37995
rect 37289 37961 37323 37995
rect 38485 37961 38519 37995
rect 41153 37961 41187 37995
rect 42717 37961 42751 37995
rect 43637 37961 43671 37995
rect 37457 37893 37491 37927
rect 37657 37893 37691 37927
rect 39598 37893 39632 37927
rect 17049 37825 17083 37859
rect 18613 37825 18647 37859
rect 18797 37825 18831 37859
rect 18889 37825 18923 37859
rect 19533 37825 19567 37859
rect 20177 37825 20211 37859
rect 21005 37825 21039 37859
rect 22937 37825 22971 37859
rect 23204 37825 23238 37859
rect 25053 37825 25087 37859
rect 25605 37825 25639 37859
rect 27353 37825 27387 37859
rect 28089 37825 28123 37859
rect 31493 37825 31527 37859
rect 32137 37825 32171 37859
rect 32229 37825 32263 37859
rect 32413 37825 32447 37859
rect 33517 37825 33551 37859
rect 33609 37825 33643 37859
rect 33793 37825 33827 37859
rect 35366 37825 35400 37859
rect 39865 37825 39899 37859
rect 41061 37825 41095 37859
rect 41245 37825 41279 37859
rect 41705 37825 41739 37859
rect 41889 37825 41923 37859
rect 42441 37825 42475 37859
rect 43545 37825 43579 37859
rect 17325 37757 17359 37791
rect 19349 37757 19383 37791
rect 20269 37757 20303 37791
rect 21281 37757 21315 37791
rect 24777 37757 24811 37791
rect 25881 37757 25915 37791
rect 27629 37757 27663 37791
rect 35633 37757 35667 37791
rect 42533 37757 42567 37791
rect 42717 37757 42751 37791
rect 19717 37689 19751 37723
rect 24317 37689 24351 37723
rect 27445 37689 27479 37723
rect 2145 37621 2179 37655
rect 17141 37621 17175 37655
rect 20177 37621 20211 37655
rect 21097 37621 21131 37655
rect 24869 37621 24903 37655
rect 24961 37621 24995 37655
rect 27353 37621 27387 37655
rect 28181 37621 28215 37655
rect 31309 37621 31343 37655
rect 32597 37621 32631 37655
rect 33241 37621 33275 37655
rect 37473 37621 37507 37655
rect 41889 37621 41923 37655
rect 18521 37417 18555 37451
rect 23397 37417 23431 37451
rect 25881 37417 25915 37451
rect 32505 37417 32539 37451
rect 32689 37417 32723 37451
rect 33517 37417 33551 37451
rect 34897 37417 34931 37451
rect 37289 37417 37323 37451
rect 41705 37417 41739 37451
rect 23765 37349 23799 37383
rect 19533 37281 19567 37315
rect 23489 37281 23523 37315
rect 23581 37281 23615 37315
rect 24961 37281 24995 37315
rect 25973 37281 26007 37315
rect 28365 37281 28399 37315
rect 28641 37281 28675 37315
rect 33057 37281 33091 37315
rect 33885 37281 33919 37315
rect 34989 37281 35023 37315
rect 41613 37281 41647 37315
rect 1409 37213 1443 37247
rect 3249 37213 3283 37247
rect 18337 37213 18371 37247
rect 19257 37213 19291 37247
rect 21005 37213 21039 37247
rect 23857 37213 23891 37247
rect 24777 37213 24811 37247
rect 25053 37213 25087 37247
rect 26157 37213 26191 37247
rect 27440 37213 27474 37247
rect 27629 37213 27663 37247
rect 27812 37213 27846 37247
rect 27905 37213 27939 37247
rect 28733 37213 28767 37247
rect 30665 37213 30699 37247
rect 30932 37213 30966 37247
rect 33701 37213 33735 37247
rect 34713 37213 34747 37247
rect 34805 37213 34839 37247
rect 37289 37213 37323 37247
rect 39313 37213 39347 37247
rect 41429 37213 41463 37247
rect 42441 37213 42475 37247
rect 3065 37145 3099 37179
rect 18153 37145 18187 37179
rect 25881 37145 25915 37179
rect 27537 37145 27571 37179
rect 32689 37145 32723 37179
rect 37013 37145 37047 37179
rect 37197 37145 37231 37179
rect 41889 37145 41923 37179
rect 42686 37145 42720 37179
rect 21097 37077 21131 37111
rect 25421 37077 25455 37111
rect 26341 37077 26375 37111
rect 27261 37077 27295 37111
rect 32045 37077 32079 37111
rect 39129 37077 39163 37111
rect 41245 37077 41279 37111
rect 43821 37077 43855 37111
rect 2697 36873 2731 36907
rect 18705 36873 18739 36907
rect 24317 36873 24351 36907
rect 25421 36873 25455 36907
rect 33241 36873 33275 36907
rect 34989 36873 35023 36907
rect 41337 36873 41371 36907
rect 41613 36873 41647 36907
rect 41705 36873 41739 36907
rect 42441 36873 42475 36907
rect 43269 36873 43303 36907
rect 17601 36805 17635 36839
rect 18613 36805 18647 36839
rect 18981 36805 19015 36839
rect 34253 36805 34287 36839
rect 37381 36805 37415 36839
rect 37565 36805 37599 36839
rect 42593 36805 42627 36839
rect 42809 36805 42843 36839
rect 2789 36737 2823 36771
rect 16865 36737 16899 36771
rect 17141 36737 17175 36771
rect 17877 36737 17911 36771
rect 19625 36737 19659 36771
rect 20453 36737 20487 36771
rect 20637 36737 20671 36771
rect 20729 36737 20763 36771
rect 21005 36737 21039 36771
rect 22109 36737 22143 36771
rect 22201 36737 22235 36771
rect 22293 36737 22327 36771
rect 22477 36737 22511 36771
rect 24225 36737 24259 36771
rect 25053 36737 25087 36771
rect 26341 36737 26375 36771
rect 26433 36737 26467 36771
rect 27716 36737 27750 36771
rect 27813 36737 27847 36771
rect 27905 36737 27939 36771
rect 28088 36737 28122 36771
rect 28181 36737 28215 36771
rect 28641 36737 28675 36771
rect 28825 36737 28859 36771
rect 28917 36737 28951 36771
rect 29193 36737 29227 36771
rect 30961 36737 30995 36771
rect 31217 36737 31251 36771
rect 32321 36737 32355 36771
rect 33333 36737 33367 36771
rect 34897 36737 34931 36771
rect 35173 36737 35207 36771
rect 38669 36737 38703 36771
rect 38936 36737 38970 36771
rect 41521 36737 41555 36771
rect 41889 36737 41923 36771
rect 43545 36737 43579 36771
rect 16773 36669 16807 36703
rect 17601 36669 17635 36703
rect 20913 36669 20947 36703
rect 24961 36669 24995 36703
rect 26157 36669 26191 36703
rect 28733 36669 28767 36703
rect 32137 36669 32171 36703
rect 32597 36669 32631 36703
rect 43269 36669 43303 36703
rect 17049 36601 17083 36635
rect 17785 36601 17819 36635
rect 18797 36601 18831 36635
rect 33885 36601 33919 36635
rect 35357 36601 35391 36635
rect 43453 36601 43487 36635
rect 16681 36533 16715 36567
rect 18889 36533 18923 36567
rect 19533 36533 19567 36567
rect 20821 36533 20855 36567
rect 21833 36533 21867 36567
rect 26249 36533 26283 36567
rect 27537 36533 27571 36567
rect 29101 36533 29135 36567
rect 29837 36533 29871 36567
rect 32505 36533 32539 36567
rect 34253 36533 34287 36567
rect 34437 36533 34471 36567
rect 40049 36533 40083 36567
rect 42625 36533 42659 36567
rect 44189 36533 44223 36567
rect 18613 36329 18647 36363
rect 21649 36329 21683 36363
rect 22109 36329 22143 36363
rect 26249 36329 26283 36363
rect 31125 36329 31159 36363
rect 33977 36329 34011 36363
rect 34805 36329 34839 36363
rect 39129 36329 39163 36363
rect 40233 36329 40267 36363
rect 20085 36261 20119 36295
rect 20177 36261 20211 36295
rect 33793 36261 33827 36295
rect 38025 36261 38059 36295
rect 39313 36261 39347 36295
rect 18705 36193 18739 36227
rect 33333 36193 33367 36227
rect 36185 36193 36219 36227
rect 36645 36193 36679 36227
rect 38669 36193 38703 36227
rect 41061 36193 41095 36227
rect 42717 36193 42751 36227
rect 44189 36193 44223 36227
rect 15945 36125 15979 36159
rect 16212 36125 16246 36159
rect 17785 36125 17819 36159
rect 18429 36125 18463 36159
rect 18521 36125 18555 36159
rect 19809 36125 19843 36159
rect 19993 36125 20027 36159
rect 20269 36125 20303 36159
rect 21005 36125 21039 36159
rect 21098 36125 21132 36159
rect 21470 36125 21504 36159
rect 22247 36125 22281 36159
rect 22385 36125 22419 36159
rect 22660 36125 22694 36159
rect 22753 36125 22787 36159
rect 23489 36125 23523 36159
rect 25697 36125 25731 36159
rect 26157 36125 26191 36159
rect 26341 36125 26375 36159
rect 27169 36125 27203 36159
rect 27332 36125 27366 36159
rect 27448 36122 27482 36156
rect 27557 36125 27591 36159
rect 28273 36125 28307 36159
rect 30941 36125 30975 36159
rect 31309 36125 31343 36159
rect 31401 36125 31435 36159
rect 38761 36125 38795 36159
rect 39129 36125 39163 36159
rect 40049 36125 40083 36159
rect 40233 36125 40267 36159
rect 40877 36125 40911 36159
rect 41521 36125 41555 36159
rect 41705 36125 41739 36159
rect 21281 36057 21315 36091
rect 21373 36057 21407 36091
rect 22477 36057 22511 36091
rect 33149 36057 33183 36091
rect 34161 36057 34195 36091
rect 35918 36057 35952 36091
rect 36890 36057 36924 36091
rect 44005 36057 44039 36091
rect 17325 35989 17359 36023
rect 17877 35989 17911 36023
rect 23673 35989 23707 36023
rect 25605 35989 25639 36023
rect 27813 35989 27847 36023
rect 28365 35989 28399 36023
rect 33961 35989 33995 36023
rect 39865 35989 39899 36023
rect 40693 35989 40727 36023
rect 41613 35989 41647 36023
rect 19073 35785 19107 35819
rect 31493 35785 31527 35819
rect 39313 35785 39347 35819
rect 40693 35785 40727 35819
rect 41889 35785 41923 35819
rect 43361 35785 43395 35819
rect 22017 35717 22051 35751
rect 22201 35717 22235 35751
rect 23866 35717 23900 35751
rect 33425 35717 33459 35751
rect 36737 35717 36771 35751
rect 37289 35717 37323 35751
rect 39497 35717 39531 35751
rect 40325 35717 40359 35751
rect 18705 35649 18739 35683
rect 20361 35649 20395 35683
rect 24133 35649 24167 35683
rect 26985 35649 27019 35683
rect 27169 35649 27203 35683
rect 27813 35649 27847 35683
rect 31401 35649 31435 35683
rect 32597 35649 32631 35683
rect 33701 35649 33735 35683
rect 34345 35649 34379 35683
rect 35265 35649 35299 35683
rect 36461 35649 36495 35683
rect 36553 35649 36587 35683
rect 37565 35649 37599 35683
rect 38577 35649 38611 35683
rect 38853 35649 38887 35683
rect 40509 35649 40543 35683
rect 40785 35649 40819 35683
rect 41613 35649 41647 35683
rect 41705 35649 41739 35683
rect 43269 35649 43303 35683
rect 18613 35581 18647 35615
rect 20269 35581 20303 35615
rect 20729 35581 20763 35615
rect 33517 35581 33551 35615
rect 34437 35581 34471 35615
rect 37289 35581 37323 35615
rect 32781 35513 32815 35547
rect 33885 35513 33919 35547
rect 35449 35513 35483 35547
rect 36737 35513 36771 35547
rect 39865 35513 39899 35547
rect 22753 35445 22787 35479
rect 27077 35445 27111 35479
rect 27905 35445 27939 35479
rect 33425 35445 33459 35479
rect 34437 35445 34471 35479
rect 34713 35445 34747 35479
rect 37473 35445 37507 35479
rect 39497 35445 39531 35479
rect 44097 35445 44131 35479
rect 22201 35241 22235 35275
rect 22937 35241 22971 35275
rect 23121 35241 23155 35275
rect 23673 35241 23707 35275
rect 27813 35241 27847 35275
rect 28733 35241 28767 35275
rect 34069 35241 34103 35275
rect 36001 35241 36035 35275
rect 41889 35241 41923 35275
rect 27997 35173 28031 35207
rect 29561 35173 29595 35207
rect 33517 35173 33551 35207
rect 35357 35173 35391 35207
rect 38485 35173 38519 35207
rect 39037 35173 39071 35207
rect 26801 35105 26835 35139
rect 27721 35105 27755 35139
rect 30941 35105 30975 35139
rect 32321 35105 32355 35139
rect 40509 35105 40543 35139
rect 42717 35105 42751 35139
rect 44189 35105 44223 35139
rect 19993 35037 20027 35071
rect 22109 35037 22143 35071
rect 24777 35037 24811 35071
rect 25605 35037 25639 35071
rect 25973 35037 26007 35071
rect 26525 35037 26559 35071
rect 26709 35037 26743 35071
rect 27813 35037 27847 35071
rect 32505 35037 32539 35071
rect 32597 35037 32631 35071
rect 33977 35037 34011 35071
rect 34161 35037 34195 35071
rect 40776 35037 40810 35071
rect 17233 34969 17267 35003
rect 17417 34969 17451 35003
rect 22753 34969 22787 35003
rect 23765 34969 23799 35003
rect 27537 34969 27571 35003
rect 28549 34969 28583 35003
rect 28765 34969 28799 35003
rect 30674 34969 30708 35003
rect 33333 34969 33367 35003
rect 35173 34969 35207 35003
rect 35909 34969 35943 35003
rect 38761 34969 38795 35003
rect 38853 34969 38887 35003
rect 44005 34969 44039 35003
rect 17601 34901 17635 34935
rect 19809 34901 19843 34935
rect 22963 34901 22997 34935
rect 24961 34901 24995 34935
rect 28917 34901 28951 34935
rect 32321 34901 32355 34935
rect 38669 34901 38703 34935
rect 16129 34697 16163 34731
rect 18061 34697 18095 34731
rect 19901 34697 19935 34731
rect 22845 34697 22879 34731
rect 23857 34697 23891 34731
rect 26065 34697 26099 34731
rect 29193 34697 29227 34731
rect 29653 34697 29687 34731
rect 30757 34697 30791 34731
rect 32889 34697 32923 34731
rect 38761 34697 38795 34731
rect 41245 34697 41279 34731
rect 43637 34697 43671 34731
rect 16926 34629 16960 34663
rect 21097 34629 21131 34663
rect 21281 34629 21315 34663
rect 22201 34629 22235 34663
rect 23121 34629 23155 34663
rect 24952 34629 24986 34663
rect 28917 34629 28951 34663
rect 32689 34629 32723 34663
rect 15945 34561 15979 34595
rect 18521 34561 18555 34595
rect 18705 34561 18739 34595
rect 18889 34561 18923 34595
rect 19533 34561 19567 34595
rect 19717 34561 19751 34595
rect 23029 34561 23063 34595
rect 23213 34561 23247 34595
rect 23397 34561 23431 34595
rect 23857 34561 23891 34595
rect 24041 34561 24075 34595
rect 24685 34561 24719 34595
rect 27353 34561 27387 34595
rect 27629 34561 27663 34595
rect 28641 34561 28675 34595
rect 28825 34561 28859 34595
rect 29009 34561 29043 34595
rect 29653 34561 29687 34595
rect 29837 34561 29871 34595
rect 30481 34561 30515 34595
rect 30573 34561 30607 34595
rect 37381 34561 37415 34595
rect 38669 34561 38703 34595
rect 38945 34561 38979 34595
rect 39957 34561 39991 34595
rect 40141 34561 40175 34595
rect 41521 34561 41555 34595
rect 43545 34561 43579 34595
rect 16681 34493 16715 34527
rect 22385 34493 22419 34527
rect 37657 34493 37691 34527
rect 39865 34493 39899 34527
rect 41245 34493 41279 34527
rect 41429 34425 41463 34459
rect 20913 34357 20947 34391
rect 32873 34357 32907 34391
rect 33057 34357 33091 34391
rect 39129 34357 39163 34391
rect 40325 34357 40359 34391
rect 42901 34357 42935 34391
rect 16773 34153 16807 34187
rect 19809 34153 19843 34187
rect 22937 34153 22971 34187
rect 24869 34153 24903 34187
rect 26065 34153 26099 34187
rect 27629 34153 27663 34187
rect 28365 34153 28399 34187
rect 29745 34153 29779 34187
rect 32413 34153 32447 34187
rect 36645 34153 36679 34187
rect 38761 34153 38795 34187
rect 21005 34085 21039 34119
rect 31953 34085 31987 34119
rect 33517 34085 33551 34119
rect 15393 34017 15427 34051
rect 17509 34017 17543 34051
rect 20453 34017 20487 34051
rect 21465 34017 21499 34051
rect 26525 34017 26559 34051
rect 30573 34017 30607 34051
rect 32781 34017 32815 34051
rect 35357 34017 35391 34051
rect 37381 34017 37415 34051
rect 39957 34017 39991 34051
rect 42349 34017 42383 34051
rect 44097 34017 44131 34051
rect 17785 33949 17819 33983
rect 19993 33949 20027 33983
rect 20177 33949 20211 33983
rect 20295 33949 20329 33983
rect 21557 33949 21591 33983
rect 22201 33949 22235 33983
rect 22385 33949 22419 33983
rect 22845 33949 22879 33983
rect 25053 33949 25087 33983
rect 25145 33949 25179 33983
rect 25697 33949 25731 33983
rect 25881 33949 25915 33983
rect 26709 33949 26743 33983
rect 26893 33949 26927 33983
rect 27169 33949 27203 33983
rect 27629 33949 27663 33983
rect 27813 33949 27847 33983
rect 28273 33949 28307 33983
rect 29561 33949 29595 33983
rect 32597 33949 32631 33983
rect 33701 33949 33735 33983
rect 34713 33949 34747 33983
rect 34897 33949 34931 33983
rect 35541 33949 35575 33983
rect 35633 33949 35667 33983
rect 36093 33949 36127 33983
rect 37105 33949 37139 33983
rect 37197 33949 37231 33983
rect 38393 33949 38427 33983
rect 40224 33949 40258 33983
rect 15660 33881 15694 33915
rect 20085 33881 20119 33915
rect 21005 33881 21039 33915
rect 21741 33881 21775 33915
rect 26801 33881 26835 33915
rect 27031 33881 27065 33915
rect 30840 33881 30874 33915
rect 33793 33881 33827 33915
rect 36461 33881 36495 33915
rect 38761 33881 38795 33915
rect 42533 33881 42567 33915
rect 22293 33813 22327 33847
rect 33885 33813 33919 33847
rect 34069 33813 34103 33847
rect 34805 33813 34839 33847
rect 35357 33813 35391 33847
rect 36277 33813 36311 33847
rect 36369 33813 36403 33847
rect 37381 33813 37415 33847
rect 38945 33813 38979 33847
rect 41337 33813 41371 33847
rect 18797 33609 18831 33643
rect 38409 33609 38443 33643
rect 38577 33609 38611 33643
rect 39773 33609 39807 33643
rect 43545 33609 43579 33643
rect 18429 33541 18463 33575
rect 19502 33541 19536 33575
rect 21189 33541 21223 33575
rect 23581 33541 23615 33575
rect 24501 33541 24535 33575
rect 24685 33541 24719 33575
rect 29653 33541 29687 33575
rect 31493 33541 31527 33575
rect 34253 33541 34287 33575
rect 36461 33541 36495 33575
rect 37749 33541 37783 33575
rect 38209 33541 38243 33575
rect 39865 33541 39899 33575
rect 15945 33473 15979 33507
rect 16129 33473 16163 33507
rect 16957 33473 16991 33507
rect 18245 33473 18279 33507
rect 18521 33473 18555 33507
rect 18613 33473 18647 33507
rect 21097 33473 21131 33507
rect 21281 33473 21315 33507
rect 22845 33473 22879 33507
rect 22937 33473 22971 33507
rect 23673 33473 23707 33507
rect 25973 33473 26007 33507
rect 26985 33473 27019 33507
rect 27169 33473 27203 33507
rect 27905 33473 27939 33507
rect 28089 33473 28123 33507
rect 29469 33473 29503 33507
rect 31401 33473 31435 33507
rect 31585 33473 31619 33507
rect 32137 33473 32171 33507
rect 32404 33473 32438 33507
rect 33977 33473 34011 33507
rect 35633 33473 35667 33507
rect 37289 33473 37323 33507
rect 37381 33473 37415 33507
rect 37565 33473 37599 33507
rect 39497 33473 39531 33507
rect 39957 33473 39991 33507
rect 42993 33473 43027 33507
rect 43453 33473 43487 33507
rect 17233 33405 17267 33439
rect 19257 33405 19291 33439
rect 22661 33405 22695 33439
rect 22753 33405 22787 33439
rect 27997 33405 28031 33439
rect 28181 33405 28215 33439
rect 34253 33405 34287 33439
rect 35357 33405 35391 33439
rect 36093 33405 36127 33439
rect 20637 33337 20671 33371
rect 25789 33337 25823 33371
rect 33517 33337 33551 33371
rect 34069 33337 34103 33371
rect 16037 33269 16071 33303
rect 22477 33269 22511 33303
rect 27077 33269 27111 33303
rect 27721 33269 27755 33303
rect 36461 33269 36495 33303
rect 36645 33269 36679 33303
rect 38393 33269 38427 33303
rect 42901 33269 42935 33303
rect 16221 33065 16255 33099
rect 19441 33065 19475 33099
rect 23857 33065 23891 33099
rect 26065 33065 26099 33099
rect 32137 33065 32171 33099
rect 32689 33065 32723 33099
rect 35265 33065 35299 33099
rect 35541 33065 35575 33099
rect 36461 33065 36495 33099
rect 36645 33065 36679 33099
rect 27261 32997 27295 33031
rect 34161 32997 34195 33031
rect 37289 32997 37323 33031
rect 15669 32929 15703 32963
rect 17877 32929 17911 32963
rect 32045 32929 32079 32963
rect 32229 32929 32263 32963
rect 38669 32929 38703 32963
rect 42533 32929 42567 32963
rect 44097 32929 44131 32963
rect 15761 32861 15795 32895
rect 16497 32861 16531 32895
rect 16589 32861 16623 32895
rect 16681 32861 16715 32895
rect 16865 32861 16899 32895
rect 18061 32861 18095 32895
rect 19257 32861 19291 32895
rect 19441 32861 19475 32895
rect 22477 32861 22511 32895
rect 24685 32861 24719 32895
rect 26801 32861 26835 32895
rect 27077 32861 27111 32895
rect 27721 32861 27755 32895
rect 27905 32861 27939 32895
rect 27997 32861 28031 32895
rect 28089 32861 28123 32895
rect 31953 32861 31987 32895
rect 32689 32861 32723 32895
rect 32873 32861 32907 32895
rect 33977 32861 34011 32895
rect 35449 32861 35483 32895
rect 35817 32861 35851 32895
rect 35909 32861 35943 32895
rect 39129 32861 39163 32895
rect 42349 32861 42383 32895
rect 18245 32793 18279 32827
rect 22744 32793 22778 32827
rect 24952 32793 24986 32827
rect 36613 32793 36647 32827
rect 36829 32793 36863 32827
rect 38402 32793 38436 32827
rect 26893 32725 26927 32759
rect 28365 32725 28399 32759
rect 39313 32725 39347 32759
rect 22845 32521 22879 32555
rect 24961 32521 24995 32555
rect 27353 32521 27387 32555
rect 28641 32521 28675 32555
rect 33425 32521 33459 32555
rect 35449 32521 35483 32555
rect 36185 32521 36219 32555
rect 37381 32521 37415 32555
rect 38853 32521 38887 32555
rect 17877 32453 17911 32487
rect 23673 32453 23707 32487
rect 24409 32453 24443 32487
rect 29754 32453 29788 32487
rect 34560 32453 34594 32487
rect 35265 32453 35299 32487
rect 15577 32385 15611 32419
rect 15945 32385 15979 32419
rect 16129 32385 16163 32419
rect 16865 32385 16899 32419
rect 18245 32385 18279 32419
rect 18981 32385 19015 32419
rect 19165 32385 19199 32419
rect 19257 32385 19291 32419
rect 19349 32385 19383 32419
rect 21097 32385 21131 32419
rect 21281 32385 21315 32419
rect 22201 32385 22235 32419
rect 22385 32385 22419 32419
rect 22477 32385 22511 32419
rect 22569 32385 22603 32419
rect 23489 32385 23523 32419
rect 23765 32385 23799 32419
rect 25237 32385 25271 32419
rect 25326 32391 25360 32425
rect 25421 32388 25455 32422
rect 25605 32385 25639 32419
rect 26249 32385 26283 32419
rect 27169 32385 27203 32419
rect 27445 32385 27479 32419
rect 27905 32385 27939 32419
rect 28089 32385 28123 32419
rect 30665 32385 30699 32419
rect 35541 32385 35575 32419
rect 36001 32385 36035 32419
rect 37289 32385 37323 32419
rect 37473 32385 37507 32419
rect 39966 32385 40000 32419
rect 40233 32385 40267 32419
rect 43637 32385 43671 32419
rect 15761 32317 15795 32351
rect 15853 32317 15887 32351
rect 17049 32317 17083 32351
rect 17969 32317 18003 32351
rect 18337 32317 18371 32351
rect 23305 32317 23339 32351
rect 27997 32317 28031 32351
rect 30021 32317 30055 32351
rect 34805 32317 34839 32351
rect 16681 32249 16715 32283
rect 18521 32249 18555 32283
rect 24225 32249 24259 32283
rect 26985 32249 27019 32283
rect 30481 32249 30515 32283
rect 15393 32181 15427 32215
rect 19625 32181 19659 32215
rect 21189 32181 21223 32215
rect 26433 32181 26467 32215
rect 35265 32181 35299 32215
rect 18521 31977 18555 32011
rect 22661 31977 22695 32011
rect 23305 31977 23339 32011
rect 24685 31977 24719 32011
rect 25881 31977 25915 32011
rect 28641 31977 28675 32011
rect 36185 31977 36219 32011
rect 15485 31909 15519 31943
rect 18337 31909 18371 31943
rect 29837 31909 29871 31943
rect 16129 31841 16163 31875
rect 16313 31841 16347 31875
rect 27261 31841 27295 31875
rect 14105 31773 14139 31807
rect 16221 31773 16255 31807
rect 16405 31773 16439 31807
rect 17049 31773 17083 31807
rect 17325 31773 17359 31807
rect 17601 31773 17635 31807
rect 17785 31773 17819 31807
rect 20637 31773 20671 31807
rect 21189 31773 21223 31807
rect 21373 31773 21407 31807
rect 22201 31773 22235 31807
rect 22477 31773 22511 31807
rect 24593 31773 24627 31807
rect 24777 31773 24811 31807
rect 27517 31773 27551 31807
rect 29653 31773 29687 31807
rect 31421 31773 31455 31807
rect 31677 31773 31711 31807
rect 34805 31773 34839 31807
rect 35072 31773 35106 31807
rect 36829 31773 36863 31807
rect 14372 31705 14406 31739
rect 18705 31705 18739 31739
rect 20370 31705 20404 31739
rect 22293 31705 22327 31739
rect 23284 31705 23318 31739
rect 23489 31705 23523 31739
rect 25973 31705 26007 31739
rect 15945 31637 15979 31671
rect 17601 31637 17635 31671
rect 18505 31637 18539 31671
rect 19257 31637 19291 31671
rect 23121 31637 23155 31671
rect 30297 31637 30331 31671
rect 36645 31637 36679 31671
rect 16037 31433 16071 31467
rect 23397 31433 23431 31467
rect 27235 31433 27269 31467
rect 31585 31433 31619 31467
rect 32137 31433 32171 31467
rect 24593 31365 24627 31399
rect 27445 31365 27479 31399
rect 31217 31365 31251 31399
rect 31417 31365 31451 31399
rect 35173 31365 35207 31399
rect 14188 31297 14222 31331
rect 15853 31297 15887 31331
rect 16129 31297 16163 31331
rect 16681 31297 16715 31331
rect 16957 31297 16991 31331
rect 19901 31297 19935 31331
rect 20168 31297 20202 31331
rect 22284 31297 22318 31331
rect 25605 31297 25639 31331
rect 26341 31297 26375 31331
rect 28273 31297 28307 31331
rect 30205 31297 30239 31331
rect 32321 31297 32355 31331
rect 13921 31229 13955 31263
rect 18981 31229 19015 31263
rect 19257 31229 19291 31263
rect 22017 31229 22051 31263
rect 29929 31229 29963 31263
rect 15853 31161 15887 31195
rect 24777 31161 24811 31195
rect 27077 31161 27111 31195
rect 34989 31161 35023 31195
rect 15301 31093 15335 31127
rect 21281 31093 21315 31127
rect 25329 31093 25363 31127
rect 26157 31093 26191 31127
rect 27261 31093 27295 31127
rect 28089 31093 28123 31127
rect 31401 31093 31435 31127
rect 15485 30889 15519 30923
rect 16681 30889 16715 30923
rect 17693 30889 17727 30923
rect 20269 30889 20303 30923
rect 22385 30889 22419 30923
rect 23765 30889 23799 30923
rect 25513 30889 25547 30923
rect 28273 30889 28307 30923
rect 28457 30889 28491 30923
rect 31125 30889 31159 30923
rect 37381 30889 37415 30923
rect 15853 30821 15887 30855
rect 26617 30821 26651 30855
rect 15761 30753 15795 30787
rect 17969 30753 18003 30787
rect 18153 30753 18187 30787
rect 24593 30753 24627 30787
rect 24777 30753 24811 30787
rect 27537 30753 27571 30787
rect 1777 30685 1811 30719
rect 15669 30685 15703 30719
rect 15945 30685 15979 30719
rect 16129 30685 16163 30719
rect 16773 30685 16807 30719
rect 17877 30685 17911 30719
rect 18061 30685 18095 30719
rect 19257 30685 19291 30719
rect 20545 30685 20579 30719
rect 20637 30685 20671 30719
rect 20729 30685 20763 30719
rect 20913 30685 20947 30719
rect 22569 30685 22603 30719
rect 24501 30685 24535 30719
rect 24685 30685 24719 30719
rect 25789 30685 25823 30719
rect 27445 30685 27479 30719
rect 30665 30685 30699 30719
rect 30941 30685 30975 30719
rect 31585 30685 31619 30719
rect 31764 30685 31798 30719
rect 31864 30682 31898 30716
rect 31953 30685 31987 30719
rect 32781 30685 32815 30719
rect 36001 30685 36035 30719
rect 36268 30685 36302 30719
rect 23673 30617 23707 30651
rect 26433 30617 26467 30651
rect 28089 30617 28123 30651
rect 30757 30617 30791 30651
rect 32229 30617 32263 30651
rect 33026 30617 33060 30651
rect 43729 30617 43763 30651
rect 44097 30617 44131 30651
rect 19349 30549 19383 30583
rect 24961 30549 24995 30583
rect 27077 30549 27111 30583
rect 28299 30549 28333 30583
rect 34161 30549 34195 30583
rect 26341 30345 26375 30379
rect 30481 30345 30515 30379
rect 18153 30277 18187 30311
rect 22477 30277 22511 30311
rect 25973 30277 26007 30311
rect 26189 30277 26223 30311
rect 28080 30277 28114 30311
rect 31585 30277 31619 30311
rect 33026 30277 33060 30311
rect 36185 30277 36219 30311
rect 1777 30209 1811 30243
rect 17049 30209 17083 30243
rect 17141 30209 17175 30243
rect 17325 30209 17359 30243
rect 18056 30209 18090 30243
rect 18245 30209 18279 30243
rect 18428 30209 18462 30243
rect 18521 30209 18555 30243
rect 22293 30209 22327 30243
rect 24317 30209 24351 30243
rect 24501 30209 24535 30243
rect 25145 30209 25179 30243
rect 27169 30209 27203 30243
rect 30021 30209 30055 30243
rect 30481 30209 30515 30243
rect 30941 30209 30975 30243
rect 31125 30209 31159 30243
rect 31217 30209 31251 30243
rect 31355 30209 31389 30243
rect 32137 30209 32171 30243
rect 32321 30209 32355 30243
rect 34897 30209 34931 30243
rect 37473 30209 37507 30243
rect 43361 30209 43395 30243
rect 1961 30141 1995 30175
rect 2789 30141 2823 30175
rect 24225 30141 24259 30175
rect 24409 30141 24443 30175
rect 27813 30141 27847 30175
rect 32781 30141 32815 30175
rect 34621 30141 34655 30175
rect 17325 30073 17359 30107
rect 17877 30073 17911 30107
rect 25329 30073 25363 30107
rect 27077 30073 27111 30107
rect 32229 30073 32263 30107
rect 36369 30073 36403 30107
rect 24685 30005 24719 30039
rect 26157 30005 26191 30039
rect 29193 30005 29227 30039
rect 30159 30005 30193 30039
rect 30297 30005 30331 30039
rect 34161 30005 34195 30039
rect 37289 30005 37323 30039
rect 43453 30005 43487 30039
rect 44189 30005 44223 30039
rect 2237 29801 2271 29835
rect 15853 29801 15887 29835
rect 16773 29801 16807 29835
rect 18153 29801 18187 29835
rect 19257 29801 19291 29835
rect 20637 29801 20671 29835
rect 28273 29801 28307 29835
rect 28825 29801 28859 29835
rect 30665 29801 30699 29835
rect 34069 29733 34103 29767
rect 17693 29665 17727 29699
rect 30757 29665 30791 29699
rect 31493 29665 31527 29699
rect 42717 29665 42751 29699
rect 44005 29665 44039 29699
rect 44189 29665 44223 29699
rect 2329 29597 2363 29631
rect 14473 29597 14507 29631
rect 15761 29597 15795 29631
rect 15945 29597 15979 29631
rect 16589 29597 16623 29631
rect 17601 29597 17635 29631
rect 17877 29597 17911 29631
rect 17969 29597 18003 29631
rect 19441 29597 19475 29631
rect 19809 29597 19843 29631
rect 20453 29597 20487 29631
rect 25697 29597 25731 29631
rect 25964 29597 25998 29631
rect 27905 29597 27939 29631
rect 28733 29597 28767 29631
rect 28917 29597 28951 29631
rect 30481 29597 30515 29631
rect 30573 29597 30607 29631
rect 31217 29597 31251 29631
rect 32781 29597 32815 29631
rect 34897 29597 34931 29631
rect 36665 29597 36699 29631
rect 36921 29597 36955 29631
rect 16405 29529 16439 29563
rect 19533 29529 19567 29563
rect 19625 29529 19659 29563
rect 28089 29529 28123 29563
rect 33333 29529 33367 29563
rect 34069 29529 34103 29563
rect 34989 29529 35023 29563
rect 14289 29461 14323 29495
rect 27077 29461 27111 29495
rect 32689 29461 32723 29495
rect 33517 29461 33551 29495
rect 33609 29461 33643 29495
rect 35541 29461 35575 29495
rect 17877 29257 17911 29291
rect 18889 29257 18923 29291
rect 29561 29257 29595 29291
rect 30573 29257 30607 29291
rect 31585 29257 31619 29291
rect 24593 29189 24627 29223
rect 25237 29189 25271 29223
rect 25437 29189 25471 29223
rect 36001 29189 36035 29223
rect 13645 29121 13679 29155
rect 13912 29121 13946 29155
rect 17049 29121 17083 29155
rect 18061 29121 18095 29155
rect 18153 29121 18187 29155
rect 18429 29121 18463 29155
rect 18889 29121 18923 29155
rect 19073 29121 19107 29155
rect 20269 29121 20303 29155
rect 22089 29121 22123 29155
rect 28825 29121 28859 29155
rect 29469 29121 29503 29155
rect 29653 29121 29687 29155
rect 31125 29121 31159 29155
rect 31217 29121 31251 29155
rect 32321 29121 32355 29155
rect 32505 29121 32539 29155
rect 33517 29121 33551 29155
rect 33885 29121 33919 29155
rect 33977 29121 34011 29155
rect 35817 29121 35851 29155
rect 36461 29121 36495 29155
rect 36645 29121 36679 29155
rect 17325 29053 17359 29087
rect 21833 29053 21867 29087
rect 30113 29053 30147 29087
rect 31309 29053 31343 29087
rect 31401 29053 31435 29087
rect 15025 28985 15059 29019
rect 16865 28985 16899 29019
rect 18337 28985 18371 29019
rect 20085 28985 20119 29019
rect 24225 28985 24259 29019
rect 24777 28985 24811 29019
rect 25605 28985 25639 29019
rect 28733 28985 28767 29019
rect 30389 28985 30423 29019
rect 34161 28985 34195 29019
rect 17233 28917 17267 28951
rect 23213 28917 23247 28951
rect 24593 28917 24627 28951
rect 25421 28917 25455 28951
rect 32137 28917 32171 28951
rect 33609 28917 33643 28951
rect 35633 28917 35667 28951
rect 36553 28917 36587 28951
rect 21281 28713 21315 28747
rect 21925 28713 21959 28747
rect 27721 28713 27755 28747
rect 27905 28713 27939 28747
rect 34989 28713 35023 28747
rect 35725 28713 35759 28747
rect 35909 28713 35943 28747
rect 15669 28645 15703 28679
rect 17693 28645 17727 28679
rect 25789 28645 25823 28679
rect 16497 28577 16531 28611
rect 17601 28577 17635 28611
rect 17969 28577 18003 28611
rect 18521 28577 18555 28611
rect 18705 28577 18739 28611
rect 24409 28577 24443 28611
rect 26157 28577 26191 28611
rect 30941 28577 30975 28611
rect 31309 28577 31343 28611
rect 33609 28577 33643 28611
rect 14289 28509 14323 28543
rect 16589 28509 16623 28543
rect 17509 28509 17543 28543
rect 17785 28509 17819 28543
rect 18429 28509 18463 28543
rect 19901 28509 19935 28543
rect 22293 28509 22327 28543
rect 22845 28509 22879 28543
rect 23029 28509 23063 28543
rect 23121 28509 23155 28543
rect 23213 28509 23247 28543
rect 24685 28509 24719 28543
rect 26801 28509 26835 28543
rect 27077 28509 27111 28543
rect 28733 28509 28767 28543
rect 30205 28509 30239 28543
rect 30481 28509 30515 28543
rect 32045 28509 32079 28543
rect 32229 28509 32263 28543
rect 32321 28509 32355 28543
rect 33333 28509 33367 28543
rect 34989 28509 35023 28543
rect 35081 28509 35115 28543
rect 36461 28509 36495 28543
rect 43453 28509 43487 28543
rect 14556 28441 14590 28475
rect 16773 28441 16807 28475
rect 20168 28441 20202 28475
rect 26893 28441 26927 28475
rect 27889 28441 27923 28475
rect 28089 28441 28123 28475
rect 30021 28441 30055 28475
rect 31426 28441 31460 28475
rect 35541 28441 35575 28475
rect 35757 28441 35791 28475
rect 36728 28441 36762 28475
rect 16129 28373 16163 28407
rect 18705 28373 18739 28407
rect 21741 28373 21775 28407
rect 21925 28373 21959 28407
rect 23489 28373 23523 28407
rect 25697 28373 25731 28407
rect 27261 28373 27295 28407
rect 28549 28373 28583 28407
rect 30389 28373 30423 28407
rect 31217 28373 31251 28407
rect 31585 28373 31619 28407
rect 34713 28373 34747 28407
rect 37841 28373 37875 28407
rect 43545 28373 43579 28407
rect 14841 28169 14875 28203
rect 16037 28169 16071 28203
rect 21189 28169 21223 28203
rect 22201 28169 22235 28203
rect 24501 28169 24535 28203
rect 25789 28169 25823 28203
rect 27353 28169 27387 28203
rect 27537 28169 27571 28203
rect 29193 28169 29227 28203
rect 30573 28169 30607 28203
rect 33793 28169 33827 28203
rect 36737 28169 36771 28203
rect 17509 28101 17543 28135
rect 22569 28101 22603 28135
rect 26065 28101 26099 28135
rect 30205 28101 30239 28135
rect 30405 28101 30439 28135
rect 15025 28033 15059 28067
rect 16129 28033 16163 28067
rect 17325 28033 17359 28067
rect 17601 28033 17635 28067
rect 18061 28033 18095 28067
rect 19533 28033 19567 28067
rect 20821 28033 20855 28067
rect 21281 28033 21315 28067
rect 22385 28033 22419 28067
rect 22661 28033 22695 28067
rect 23121 28033 23155 28067
rect 23388 28033 23422 28067
rect 25145 28033 25179 28067
rect 26433 28033 26467 28067
rect 28365 28033 28399 28067
rect 28549 28033 28583 28067
rect 29561 28033 29595 28067
rect 31309 28033 31343 28067
rect 31585 28033 31619 28067
rect 32413 28033 32447 28067
rect 32680 28033 32714 28067
rect 34437 28033 34471 28067
rect 34621 28033 34655 28067
rect 36093 28033 36127 28067
rect 36277 28033 36311 28067
rect 36369 28033 36403 28067
rect 36461 28033 36495 28067
rect 37473 28033 37507 28067
rect 15209 27965 15243 27999
rect 18337 27965 18371 27999
rect 25948 27965 25982 27999
rect 26157 27965 26191 27999
rect 27905 27965 27939 27999
rect 28733 27965 28767 27999
rect 29469 27965 29503 27999
rect 34253 27965 34287 27999
rect 31033 27897 31067 27931
rect 17141 27829 17175 27863
rect 19441 27829 19475 27863
rect 21005 27829 21039 27863
rect 25329 27829 25363 27863
rect 27537 27829 27571 27863
rect 29561 27829 29595 27863
rect 30389 27829 30423 27863
rect 31493 27829 31527 27863
rect 37381 27829 37415 27863
rect 43821 27829 43855 27863
rect 16313 27625 16347 27659
rect 17233 27625 17267 27659
rect 17601 27625 17635 27659
rect 21097 27625 21131 27659
rect 22477 27625 22511 27659
rect 22661 27625 22695 27659
rect 23397 27625 23431 27659
rect 31033 27625 31067 27659
rect 32689 27625 32723 27659
rect 36185 27625 36219 27659
rect 16681 27557 16715 27591
rect 18245 27557 18279 27591
rect 20729 27557 20763 27591
rect 21833 27557 21867 27591
rect 27077 27557 27111 27591
rect 31585 27557 31619 27591
rect 31861 27557 31895 27591
rect 18061 27489 18095 27523
rect 21189 27489 21223 27523
rect 25697 27489 25731 27523
rect 29561 27489 29595 27523
rect 29837 27489 29871 27523
rect 42717 27489 42751 27523
rect 44005 27489 44039 27523
rect 44189 27489 44223 27523
rect 16497 27421 16531 27455
rect 16773 27421 16807 27455
rect 17417 27421 17451 27455
rect 17601 27421 17635 27455
rect 18337 27421 18371 27455
rect 20913 27421 20947 27455
rect 21649 27421 21683 27455
rect 23305 27421 23339 27455
rect 23489 27421 23523 27455
rect 25053 27421 25087 27455
rect 27629 27421 27663 27455
rect 27896 27421 27930 27455
rect 30849 27421 30883 27455
rect 31861 27421 31895 27455
rect 32045 27421 32079 27455
rect 32505 27421 32539 27455
rect 34713 27421 34747 27455
rect 34897 27421 34931 27455
rect 36093 27421 36127 27455
rect 36277 27421 36311 27455
rect 22845 27353 22879 27387
rect 25942 27353 25976 27387
rect 18337 27285 18371 27319
rect 22645 27285 22679 27319
rect 25145 27285 25179 27319
rect 29009 27285 29043 27319
rect 34805 27285 34839 27319
rect 16129 27081 16163 27115
rect 28641 27081 28675 27115
rect 29009 27081 29043 27115
rect 17279 27013 17313 27047
rect 17417 27013 17451 27047
rect 17509 27013 17543 27047
rect 18337 27013 18371 27047
rect 23121 27013 23155 27047
rect 27813 27013 27847 27047
rect 34897 27013 34931 27047
rect 36470 27013 36504 27047
rect 14749 26945 14783 26979
rect 15016 26945 15050 26979
rect 17601 26945 17635 26979
rect 18429 26945 18463 26979
rect 22937 26945 22971 26979
rect 23213 26945 23247 26979
rect 28733 26945 28767 26979
rect 28825 26945 28859 26979
rect 33609 26945 33643 26979
rect 33793 26945 33827 26979
rect 34253 26945 34287 26979
rect 34437 26945 34471 26979
rect 34529 26945 34563 26979
rect 34621 26945 34655 26979
rect 17141 26877 17175 26911
rect 27997 26877 28031 26911
rect 33333 26877 33367 26911
rect 36737 26877 36771 26911
rect 28457 26809 28491 26843
rect 33425 26809 33459 26843
rect 17785 26741 17819 26775
rect 23029 26741 23063 26775
rect 35357 26741 35391 26775
rect 15485 26537 15519 26571
rect 16681 26537 16715 26571
rect 17601 26537 17635 26571
rect 28641 26537 28675 26571
rect 32229 26537 32263 26571
rect 32965 26537 32999 26571
rect 35081 26537 35115 26571
rect 23857 26469 23891 26503
rect 31033 26469 31067 26503
rect 35817 26469 35851 26503
rect 18061 26401 18095 26435
rect 19533 26401 19567 26435
rect 23305 26401 23339 26435
rect 24777 26401 24811 26435
rect 25053 26401 25087 26435
rect 33701 26401 33735 26435
rect 34713 26401 34747 26435
rect 42073 26401 42107 26435
rect 15393 26333 15427 26367
rect 15577 26333 15611 26367
rect 16773 26333 16807 26367
rect 17417 26333 17451 26367
rect 18245 26333 18279 26367
rect 18337 26333 18371 26367
rect 19257 26333 19291 26367
rect 21005 26333 21039 26367
rect 21373 26333 21407 26367
rect 22089 26333 22123 26367
rect 22201 26333 22235 26367
rect 22293 26333 22327 26367
rect 22477 26333 22511 26367
rect 23489 26333 23523 26367
rect 24685 26333 24719 26367
rect 25513 26333 25547 26367
rect 25697 26333 25731 26367
rect 25881 26333 25915 26367
rect 26525 26333 26559 26367
rect 28549 26333 28583 26367
rect 31217 26333 31251 26367
rect 31309 26333 31343 26367
rect 32137 26333 32171 26367
rect 32321 26333 32355 26367
rect 33609 26333 33643 26367
rect 33885 26333 33919 26367
rect 37197 26333 37231 26367
rect 41613 26333 41647 26367
rect 43913 26333 43947 26367
rect 17233 26265 17267 26299
rect 21097 26265 21131 26299
rect 21189 26265 21223 26299
rect 21833 26265 21867 26299
rect 31033 26265 31067 26299
rect 32781 26265 32815 26299
rect 35081 26265 35115 26299
rect 36930 26265 36964 26299
rect 41797 26265 41831 26299
rect 18061 26197 18095 26231
rect 20821 26197 20855 26231
rect 23397 26197 23431 26231
rect 26341 26197 26375 26231
rect 32991 26197 33025 26231
rect 33149 26197 33183 26231
rect 34069 26197 34103 26231
rect 35265 26197 35299 26231
rect 31125 25993 31159 26027
rect 33517 25993 33551 26027
rect 34713 25993 34747 26027
rect 35173 25993 35207 26027
rect 36001 25993 36035 26027
rect 42441 25993 42475 26027
rect 3341 25925 3375 25959
rect 24041 25925 24075 25959
rect 24501 25925 24535 25959
rect 25320 25925 25354 25959
rect 27261 25925 27295 25959
rect 33425 25925 33459 25959
rect 34345 25925 34379 25959
rect 5181 25857 5215 25891
rect 15853 25857 15887 25891
rect 15945 25857 15979 25891
rect 16129 25857 16163 25891
rect 17049 25857 17083 25891
rect 17877 25857 17911 25891
rect 18144 25857 18178 25891
rect 19717 25857 19751 25891
rect 19984 25857 20018 25891
rect 21925 25857 21959 25891
rect 22192 25857 22226 25891
rect 25053 25857 25087 25891
rect 26985 25857 27019 25891
rect 28549 25857 28583 25891
rect 28733 25857 28767 25891
rect 28825 25857 28859 25891
rect 28917 25857 28951 25891
rect 30665 25857 30699 25891
rect 31184 25857 31218 25891
rect 32321 25857 32355 25891
rect 33333 25857 33367 25891
rect 33793 25857 33827 25891
rect 34253 25857 34287 25891
rect 34529 25857 34563 25891
rect 35357 25857 35391 25891
rect 35817 25857 35851 25891
rect 37545 25857 37579 25891
rect 39221 25857 39255 25891
rect 42625 25857 42659 25891
rect 4997 25789 5031 25823
rect 16773 25789 16807 25823
rect 16957 25789 16991 25823
rect 23949 25789 23983 25823
rect 27261 25789 27295 25823
rect 32505 25789 32539 25823
rect 37289 25789 37323 25823
rect 16865 25721 16899 25755
rect 19257 25721 19291 25755
rect 23305 25721 23339 25755
rect 24501 25721 24535 25755
rect 26433 25721 26467 25755
rect 15853 25653 15887 25687
rect 21097 25653 21131 25687
rect 23765 25653 23799 25687
rect 27077 25653 27111 25687
rect 29193 25653 29227 25687
rect 30757 25653 30791 25687
rect 31309 25653 31343 25687
rect 32137 25653 32171 25687
rect 39405 25653 39439 25687
rect 43821 25653 43855 25687
rect 3893 25449 3927 25483
rect 16957 25449 16991 25483
rect 17969 25449 18003 25483
rect 18245 25449 18279 25483
rect 21281 25449 21315 25483
rect 22109 25449 22143 25483
rect 26295 25449 26329 25483
rect 27629 25449 27663 25483
rect 29653 25449 29687 25483
rect 29745 25449 29779 25483
rect 30573 25449 30607 25483
rect 38945 25449 38979 25483
rect 25237 25381 25271 25415
rect 30757 25381 30791 25415
rect 32781 25381 32815 25415
rect 15577 25313 15611 25347
rect 18153 25313 18187 25347
rect 19993 25313 20027 25347
rect 21097 25313 21131 25347
rect 23581 25313 23615 25347
rect 24777 25313 24811 25347
rect 26525 25313 26559 25347
rect 28733 25313 28767 25347
rect 29745 25313 29779 25347
rect 31309 25313 31343 25347
rect 31401 25313 31435 25347
rect 41337 25313 41371 25347
rect 41889 25313 41923 25347
rect 44097 25313 44131 25347
rect 3985 25245 4019 25279
rect 15844 25245 15878 25279
rect 17877 25245 17911 25279
rect 18245 25245 18279 25279
rect 20177 25245 20211 25279
rect 21005 25245 21039 25279
rect 22109 25245 22143 25279
rect 22293 25245 22327 25279
rect 23305 25245 23339 25279
rect 24685 25245 24719 25279
rect 24961 25245 24995 25279
rect 25053 25245 25087 25279
rect 26985 25245 27019 25279
rect 27169 25245 27203 25279
rect 27445 25245 27479 25279
rect 28457 25245 28491 25279
rect 28641 25245 28675 25279
rect 28825 25245 28859 25279
rect 29009 25245 29043 25279
rect 29561 25245 29595 25279
rect 31493 25245 31527 25279
rect 31585 25245 31619 25279
rect 33894 25245 33928 25279
rect 34161 25245 34195 25279
rect 39129 25245 39163 25279
rect 39313 25245 39347 25279
rect 42349 25245 42383 25279
rect 29929 25177 29963 25211
rect 30389 25177 30423 25211
rect 41705 25177 41739 25211
rect 42533 25177 42567 25211
rect 20361 25109 20395 25143
rect 28273 25109 28307 25143
rect 30589 25109 30623 25143
rect 31769 25109 31803 25143
rect 20177 24905 20211 24939
rect 39681 24905 39715 24939
rect 32137 24837 32171 24871
rect 20361 24769 20395 24803
rect 23029 24769 23063 24803
rect 23305 24769 23339 24803
rect 24685 24769 24719 24803
rect 24777 24769 24811 24803
rect 25329 24769 25363 24803
rect 25605 24769 25639 24803
rect 25697 24769 25731 24803
rect 29101 24769 29135 24803
rect 29561 24769 29595 24803
rect 30849 24769 30883 24803
rect 31033 24769 31067 24803
rect 31217 24769 31251 24803
rect 31401 24769 31435 24803
rect 32321 24769 32355 24803
rect 32413 24769 32447 24803
rect 32873 24769 32907 24803
rect 38301 24769 38335 24803
rect 38568 24769 38602 24803
rect 40397 24769 40431 24803
rect 42441 24769 42475 24803
rect 43269 24769 43303 24803
rect 43913 24769 43947 24803
rect 44005 24769 44039 24803
rect 22845 24701 22879 24735
rect 23121 24701 23155 24735
rect 23213 24701 23247 24735
rect 25421 24701 25455 24735
rect 29837 24701 29871 24735
rect 31125 24701 31159 24735
rect 40141 24701 40175 24735
rect 42533 24701 42567 24735
rect 25881 24633 25915 24667
rect 27813 24633 27847 24667
rect 31585 24565 31619 24599
rect 32137 24565 32171 24599
rect 32965 24565 32999 24599
rect 41521 24565 41555 24599
rect 43361 24565 43395 24599
rect 26157 24361 26191 24395
rect 26985 24361 27019 24395
rect 27905 24361 27939 24395
rect 28825 24361 28859 24395
rect 30205 24361 30239 24395
rect 31309 24361 31343 24395
rect 32045 24361 32079 24395
rect 32137 24361 32171 24395
rect 41061 24361 41095 24395
rect 41797 24361 41831 24395
rect 30297 24293 30331 24327
rect 15577 24225 15611 24259
rect 17969 24225 18003 24259
rect 18245 24225 18279 24259
rect 20177 24225 20211 24259
rect 20453 24225 20487 24259
rect 25237 24225 25271 24259
rect 32045 24225 32079 24259
rect 40693 24225 40727 24259
rect 42717 24225 42751 24259
rect 44005 24225 44039 24259
rect 44189 24225 44223 24259
rect 18337 24157 18371 24191
rect 23765 24157 23799 24191
rect 24961 24157 24995 24191
rect 26065 24157 26099 24191
rect 26249 24157 26283 24191
rect 26709 24157 26743 24191
rect 27445 24157 27479 24191
rect 27537 24157 27571 24191
rect 27721 24157 27755 24191
rect 28641 24157 28675 24191
rect 30389 24157 30423 24191
rect 31033 24157 31067 24191
rect 31125 24157 31159 24191
rect 31401 24157 31435 24191
rect 32229 24157 32263 24191
rect 35909 24157 35943 24191
rect 37841 24157 37875 24191
rect 38025 24157 38059 24191
rect 40877 24157 40911 24191
rect 41705 24157 41739 24191
rect 15844 24089 15878 24123
rect 23489 24089 23523 24123
rect 23673 24089 23707 24123
rect 26985 24089 27019 24123
rect 28457 24089 28491 24123
rect 30113 24089 30147 24123
rect 31861 24089 31895 24123
rect 36154 24089 36188 24123
rect 38209 24089 38243 24123
rect 16957 24021 16991 24055
rect 23587 24021 23621 24055
rect 26801 24021 26835 24055
rect 30849 24021 30883 24055
rect 17969 23817 18003 23851
rect 25053 23817 25087 23851
rect 31585 23817 31619 23851
rect 37657 23817 37691 23851
rect 38485 23817 38519 23851
rect 41061 23817 41095 23851
rect 18337 23749 18371 23783
rect 18475 23749 18509 23783
rect 22385 23749 22419 23783
rect 23918 23749 23952 23783
rect 27629 23749 27663 23783
rect 28549 23749 28583 23783
rect 32229 23749 32263 23783
rect 2145 23681 2179 23715
rect 15945 23681 15979 23715
rect 16129 23681 16163 23715
rect 17233 23681 17267 23715
rect 18153 23681 18187 23715
rect 18245 23681 18279 23715
rect 19073 23681 19107 23715
rect 19165 23681 19199 23715
rect 19349 23681 19383 23715
rect 20177 23681 20211 23715
rect 20361 23681 20395 23715
rect 20821 23681 20855 23715
rect 23673 23681 23707 23715
rect 27813 23681 27847 23715
rect 27997 23681 28031 23715
rect 29193 23681 29227 23715
rect 30389 23681 30423 23715
rect 30573 23681 30607 23715
rect 31125 23681 31159 23715
rect 31217 23681 31251 23715
rect 31401 23681 31435 23715
rect 32137 23681 32171 23715
rect 32321 23681 32355 23715
rect 33609 23681 33643 23715
rect 34069 23681 34103 23715
rect 34325 23681 34359 23715
rect 35909 23681 35943 23715
rect 37289 23681 37323 23715
rect 37473 23681 37507 23715
rect 38669 23681 38703 23715
rect 40877 23681 40911 23715
rect 41521 23681 41555 23715
rect 41705 23681 41739 23715
rect 41797 23681 41831 23715
rect 42625 23681 42659 23715
rect 43269 23681 43303 23715
rect 17049 23613 17083 23647
rect 18613 23613 18647 23647
rect 19993 23613 20027 23647
rect 28733 23613 28767 23647
rect 30481 23613 30515 23647
rect 33333 23613 33367 23647
rect 36185 23613 36219 23647
rect 38761 23613 38795 23647
rect 38853 23613 38887 23647
rect 2053 23545 2087 23579
rect 22201 23545 22235 23579
rect 31309 23545 31343 23579
rect 33517 23545 33551 23579
rect 35449 23545 35483 23579
rect 2789 23477 2823 23511
rect 16037 23477 16071 23511
rect 19349 23477 19383 23511
rect 21005 23477 21039 23511
rect 29193 23477 29227 23511
rect 33425 23477 33459 23511
rect 42441 23477 42475 23511
rect 43177 23477 43211 23511
rect 43913 23477 43947 23511
rect 16773 23273 16807 23307
rect 23581 23273 23615 23307
rect 23673 23273 23707 23307
rect 25973 23273 26007 23307
rect 26341 23273 26375 23307
rect 26985 23273 27019 23307
rect 33609 23273 33643 23307
rect 36553 23273 36587 23307
rect 41337 23273 41371 23307
rect 31125 23205 31159 23239
rect 1409 23137 1443 23171
rect 3249 23137 3283 23171
rect 17417 23137 17451 23171
rect 17693 23137 17727 23171
rect 23489 23137 23523 23171
rect 26249 23137 26283 23171
rect 28365 23137 28399 23171
rect 37105 23137 37139 23171
rect 39957 23137 39991 23171
rect 42717 23137 42751 23171
rect 44189 23137 44223 23171
rect 15393 23069 15427 23103
rect 19441 23069 19475 23103
rect 19625 23069 19659 23103
rect 19743 23069 19777 23103
rect 19901 23069 19935 23103
rect 21005 23069 21039 23103
rect 21272 23069 21306 23103
rect 23765 23069 23799 23103
rect 24409 23069 24443 23103
rect 26341 23069 26375 23103
rect 26893 23069 26927 23103
rect 28089 23069 28123 23103
rect 30205 23069 30239 23103
rect 30849 23069 30883 23103
rect 31033 23069 31067 23103
rect 33609 23069 33643 23103
rect 33885 23069 33919 23103
rect 36369 23069 36403 23103
rect 36553 23069 36587 23103
rect 37197 23069 37231 23103
rect 38669 23069 38703 23103
rect 38853 23069 38887 23103
rect 39129 23069 39163 23103
rect 3065 23001 3099 23035
rect 15660 23001 15694 23035
rect 19533 23001 19567 23035
rect 30021 23001 30055 23035
rect 30389 23001 30423 23035
rect 39313 23001 39347 23035
rect 40202 23001 40236 23035
rect 44005 23001 44039 23035
rect 19257 22933 19291 22967
rect 22385 22933 22419 22967
rect 24593 22933 24627 22967
rect 33793 22933 33827 22967
rect 37565 22933 37599 22967
rect 39405 22729 39439 22763
rect 42809 22729 42843 22763
rect 43453 22729 43487 22763
rect 16941 22661 16975 22695
rect 17141 22661 17175 22695
rect 22661 22661 22695 22695
rect 25513 22661 25547 22695
rect 28825 22661 28859 22695
rect 29929 22661 29963 22695
rect 33517 22661 33551 22695
rect 34161 22661 34195 22695
rect 39037 22661 39071 22695
rect 6377 22593 6411 22627
rect 15761 22593 15795 22627
rect 15853 22593 15887 22627
rect 15945 22593 15979 22627
rect 16129 22593 16163 22627
rect 17601 22593 17635 22627
rect 17785 22593 17819 22627
rect 18705 22593 18739 22627
rect 18972 22593 19006 22627
rect 20729 22593 20763 22627
rect 20913 22593 20947 22627
rect 22477 22593 22511 22627
rect 23489 22593 23523 22627
rect 25881 22593 25915 22627
rect 26157 22593 26191 22627
rect 27813 22593 27847 22627
rect 28917 22593 28951 22627
rect 29193 22593 29227 22627
rect 29837 22593 29871 22627
rect 30573 22593 30607 22627
rect 30849 22593 30883 22627
rect 32413 22593 32447 22627
rect 32597 22593 32631 22627
rect 34345 22593 34379 22627
rect 34529 22593 34563 22627
rect 34621 22593 34655 22627
rect 35725 22593 35759 22627
rect 36553 22593 36587 22627
rect 36737 22593 36771 22627
rect 38209 22593 38243 22627
rect 38945 22593 38979 22627
rect 39221 22593 39255 22627
rect 42625 22593 42659 22627
rect 43361 22593 43395 22627
rect 1961 22525 1995 22559
rect 2145 22525 2179 22559
rect 2973 22525 3007 22559
rect 6561 22525 6595 22559
rect 15485 22525 15519 22559
rect 25697 22525 25731 22559
rect 27537 22525 27571 22559
rect 29377 22525 29411 22559
rect 35817 22525 35851 22559
rect 36645 22525 36679 22559
rect 38301 22525 38335 22559
rect 38393 22525 38427 22559
rect 42441 22525 42475 22559
rect 23305 22457 23339 22491
rect 31125 22457 31159 22491
rect 33149 22457 33183 22491
rect 36093 22457 36127 22491
rect 16773 22389 16807 22423
rect 16957 22389 16991 22423
rect 17785 22389 17819 22423
rect 17969 22389 18003 22423
rect 20085 22389 20119 22423
rect 21097 22389 21131 22423
rect 30665 22389 30699 22423
rect 32413 22389 32447 22423
rect 33517 22389 33551 22423
rect 33701 22389 33735 22423
rect 38025 22389 38059 22423
rect 2053 22185 2087 22219
rect 33977 22185 34011 22219
rect 41797 22185 41831 22219
rect 25881 22117 25915 22151
rect 26893 22117 26927 22151
rect 30297 22117 30331 22151
rect 30481 22117 30515 22151
rect 33793 22117 33827 22151
rect 38025 22117 38059 22151
rect 2881 22049 2915 22083
rect 6469 22049 6503 22083
rect 19349 22049 19383 22083
rect 25973 22049 26007 22083
rect 26801 22049 26835 22083
rect 27629 22049 27663 22083
rect 30021 22049 30055 22083
rect 31953 22049 31987 22083
rect 42349 22049 42383 22083
rect 42533 22049 42567 22083
rect 42809 22049 42843 22083
rect 2973 21981 3007 22015
rect 6285 21981 6319 22015
rect 16037 21981 16071 22015
rect 17509 21981 17543 22015
rect 17785 21981 17819 22015
rect 19257 21981 19291 22015
rect 19441 21981 19475 22015
rect 20085 21981 20119 22015
rect 20269 21981 20303 22015
rect 20913 21981 20947 22015
rect 21557 21981 21591 22015
rect 25789 21981 25823 22015
rect 26709 21981 26743 22015
rect 26985 21981 27019 22015
rect 27905 21981 27939 22015
rect 32505 21981 32539 22015
rect 32781 21981 32815 22015
rect 34713 21981 34747 22015
rect 35633 21981 35667 22015
rect 35817 21981 35851 22015
rect 36001 21981 36035 22015
rect 37657 21981 37691 22015
rect 38853 21981 38887 22015
rect 39129 21981 39163 22015
rect 40417 21981 40451 22015
rect 15761 21913 15795 21947
rect 21802 21913 21836 21947
rect 26157 21913 26191 21947
rect 31769 21913 31803 21947
rect 32597 21913 32631 21947
rect 34161 21913 34195 21947
rect 35909 21913 35943 21947
rect 38945 21913 38979 21947
rect 40662 21913 40696 21947
rect 15859 21845 15893 21879
rect 15945 21845 15979 21879
rect 20177 21845 20211 21879
rect 21097 21845 21131 21879
rect 22937 21845 22971 21879
rect 26065 21845 26099 21879
rect 27169 21845 27203 21879
rect 31309 21845 31343 21879
rect 31677 21845 31711 21879
rect 32682 21845 32716 21879
rect 33961 21845 33995 21879
rect 34897 21845 34931 21879
rect 36185 21845 36219 21879
rect 38117 21845 38151 21879
rect 39313 21845 39347 21879
rect 8033 21641 8067 21675
rect 19809 21641 19843 21675
rect 25697 21641 25731 21675
rect 27261 21641 27295 21675
rect 33701 21641 33735 21675
rect 38209 21641 38243 21675
rect 40141 21641 40175 21675
rect 6745 21573 6779 21607
rect 18153 21573 18187 21607
rect 19257 21573 19291 21607
rect 19901 21573 19935 21607
rect 29469 21573 29503 21607
rect 34814 21573 34848 21607
rect 38761 21573 38795 21607
rect 5733 21505 5767 21539
rect 15016 21505 15050 21539
rect 17877 21505 17911 21539
rect 18061 21505 18095 21539
rect 18245 21505 18279 21539
rect 18363 21505 18397 21539
rect 18521 21505 18555 21539
rect 18981 21505 19015 21539
rect 19073 21505 19107 21539
rect 20913 21505 20947 21539
rect 21097 21505 21131 21539
rect 22017 21505 22051 21539
rect 22733 21505 22767 21539
rect 24584 21505 24618 21539
rect 27445 21505 27479 21539
rect 27721 21505 27755 21539
rect 28549 21505 28583 21539
rect 30573 21505 30607 21539
rect 31033 21505 31067 21539
rect 36369 21505 36403 21539
rect 38117 21505 38151 21539
rect 38301 21505 38335 21539
rect 39957 21505 39991 21539
rect 42441 21505 42475 21539
rect 5457 21437 5491 21471
rect 14749 21437 14783 21471
rect 20729 21437 20763 21471
rect 22477 21437 22511 21471
rect 24317 21437 24351 21471
rect 27537 21437 27571 21471
rect 28641 21437 28675 21471
rect 28917 21437 28951 21471
rect 30849 21437 30883 21471
rect 35081 21437 35115 21471
rect 36277 21437 36311 21471
rect 39221 21437 39255 21471
rect 19257 21369 19291 21403
rect 36737 21369 36771 21403
rect 39037 21369 39071 21403
rect 16129 21301 16163 21335
rect 21833 21301 21867 21335
rect 23857 21301 23891 21335
rect 27721 21301 27755 21335
rect 29561 21301 29595 21335
rect 30711 21301 30745 21335
rect 30941 21301 30975 21335
rect 42533 21301 42567 21335
rect 43637 21301 43671 21335
rect 5549 21097 5583 21131
rect 23305 21097 23339 21131
rect 24593 21097 24627 21131
rect 26065 21097 26099 21131
rect 26249 21097 26283 21131
rect 27905 21097 27939 21131
rect 28641 21097 28675 21131
rect 30205 21097 30239 21131
rect 31953 21097 31987 21131
rect 33057 21097 33091 21131
rect 38945 21097 38979 21131
rect 22845 21029 22879 21063
rect 23765 21029 23799 21063
rect 27169 21029 27203 21063
rect 35909 21029 35943 21063
rect 6837 20961 6871 20995
rect 17509 20961 17543 20995
rect 17785 20961 17819 20995
rect 19625 20961 19659 20995
rect 21465 20961 21499 20995
rect 23397 20961 23431 20995
rect 25973 20961 26007 20995
rect 29837 20961 29871 20995
rect 31401 20961 31435 20995
rect 33793 20961 33827 20995
rect 35449 20961 35483 20995
rect 40417 20961 40451 20995
rect 42349 20961 42383 20995
rect 44097 20961 44131 20995
rect 1777 20893 1811 20927
rect 5365 20893 5399 20927
rect 6101 20893 6135 20927
rect 11345 20893 11379 20927
rect 14565 20893 14599 20927
rect 14749 20893 14783 20927
rect 15393 20893 15427 20927
rect 15485 20893 15519 20927
rect 15853 20893 15887 20927
rect 16681 20893 16715 20927
rect 21732 20893 21766 20927
rect 23581 20893 23615 20927
rect 24409 20893 24443 20927
rect 25881 20893 25915 20927
rect 26893 20893 26927 20927
rect 27169 20893 27203 20927
rect 28457 20893 28491 20927
rect 28641 20893 28675 20927
rect 30021 20893 30055 20927
rect 30297 20893 30331 20927
rect 30941 20893 30975 20927
rect 31033 20893 31067 20927
rect 31309 20893 31343 20927
rect 32045 20893 32079 20927
rect 32873 20893 32907 20927
rect 33149 20893 33183 20927
rect 33609 20893 33643 20927
rect 34069 20893 34103 20927
rect 35541 20893 35575 20927
rect 38761 20893 38795 20927
rect 40601 20893 40635 20927
rect 14657 20825 14691 20859
rect 15577 20825 15611 20859
rect 15695 20825 15729 20859
rect 16865 20825 16899 20859
rect 19892 20825 19926 20859
rect 23305 20825 23339 20859
rect 27813 20825 27847 20859
rect 32689 20825 32723 20859
rect 42533 20825 42567 20859
rect 11529 20757 11563 20791
rect 15209 20757 15243 20791
rect 17049 20757 17083 20791
rect 21005 20757 21039 20791
rect 30757 20757 30791 20791
rect 33977 20757 34011 20791
rect 40785 20757 40819 20791
rect 15945 20553 15979 20587
rect 18521 20553 18555 20587
rect 19717 20553 19751 20587
rect 41061 20553 41095 20587
rect 43085 20553 43119 20587
rect 17601 20485 17635 20519
rect 19441 20485 19475 20519
rect 29386 20485 29420 20519
rect 31401 20485 31435 20519
rect 32229 20485 32263 20519
rect 1685 20417 1719 20451
rect 12357 20417 12391 20451
rect 14013 20417 14047 20451
rect 14280 20417 14314 20451
rect 16037 20417 16071 20451
rect 17325 20417 17359 20451
rect 17417 20417 17451 20451
rect 18337 20417 18371 20451
rect 19165 20417 19199 20451
rect 19349 20417 19383 20451
rect 19533 20417 19567 20451
rect 20453 20417 20487 20451
rect 23029 20417 23063 20451
rect 25309 20417 25343 20451
rect 29653 20417 29687 20451
rect 30389 20417 30423 20451
rect 31217 20417 31251 20451
rect 31309 20417 31343 20451
rect 31585 20417 31619 20451
rect 32137 20417 32171 20451
rect 32321 20417 32355 20451
rect 33885 20417 33919 20451
rect 34152 20417 34186 20451
rect 37841 20417 37875 20451
rect 38108 20417 38142 20451
rect 39681 20417 39715 20451
rect 39937 20417 39971 20451
rect 42993 20417 43027 20451
rect 1869 20349 1903 20383
rect 2789 20349 2823 20383
rect 12633 20349 12667 20383
rect 18153 20349 18187 20383
rect 20729 20349 20763 20383
rect 21833 20349 21867 20383
rect 25053 20349 25087 20383
rect 30481 20349 30515 20383
rect 22201 20281 22235 20315
rect 23397 20281 23431 20315
rect 26433 20281 26467 20315
rect 35265 20281 35299 20315
rect 15393 20213 15427 20247
rect 22293 20213 22327 20247
rect 23489 20213 23523 20247
rect 31033 20213 31067 20247
rect 39221 20213 39255 20247
rect 43637 20213 43671 20247
rect 2053 20009 2087 20043
rect 15025 20009 15059 20043
rect 15209 20009 15243 20043
rect 17233 20009 17267 20043
rect 18337 20009 18371 20043
rect 18521 20009 18555 20043
rect 20085 20009 20119 20043
rect 22293 20009 22327 20043
rect 27445 20009 27479 20043
rect 31217 20009 31251 20043
rect 20269 19941 20303 19975
rect 15853 19873 15887 19907
rect 26065 19873 26099 19907
rect 32505 19873 32539 19907
rect 32965 19873 32999 19907
rect 35449 19873 35483 19907
rect 39313 19873 39347 19907
rect 40417 19873 40451 19907
rect 42073 19873 42107 19907
rect 43085 19873 43119 19907
rect 2145 19805 2179 19839
rect 12265 19805 12299 19839
rect 16129 19805 16163 19839
rect 17141 19805 17175 19839
rect 17417 19805 17451 19839
rect 19901 19805 19935 19839
rect 19993 19805 20027 19839
rect 20729 19805 20763 19839
rect 20913 19805 20947 19839
rect 21557 19805 21591 19839
rect 22845 19805 22879 19839
rect 31033 19805 31067 19839
rect 32597 19805 32631 19839
rect 35705 19805 35739 19839
rect 39129 19805 39163 19839
rect 40141 19805 40175 19839
rect 41889 19805 41923 19839
rect 12909 19737 12943 19771
rect 15193 19737 15227 19771
rect 15393 19737 15427 19771
rect 18153 19737 18187 19771
rect 18358 19737 18392 19771
rect 22201 19737 22235 19771
rect 26332 19737 26366 19771
rect 30849 19737 30883 19771
rect 17601 19669 17635 19703
rect 20821 19669 20855 19703
rect 21465 19669 21499 19703
rect 23029 19669 23063 19703
rect 36829 19669 36863 19703
rect 38945 19669 38979 19703
rect 41521 19465 41555 19499
rect 12725 19397 12759 19431
rect 15302 19397 15336 19431
rect 15511 19397 15545 19431
rect 18429 19397 18463 19431
rect 22201 19397 22235 19431
rect 23734 19397 23768 19431
rect 30472 19397 30506 19431
rect 33578 19397 33612 19431
rect 12173 19329 12207 19363
rect 13277 19329 13311 19363
rect 13553 19329 13587 19363
rect 15025 19329 15059 19363
rect 15209 19329 15243 19363
rect 15393 19329 15427 19363
rect 18705 19329 18739 19363
rect 19533 19329 19567 19363
rect 19625 19329 19659 19363
rect 19809 19329 19843 19363
rect 19901 19329 19935 19363
rect 20361 19329 20395 19363
rect 20637 19329 20671 19363
rect 23489 19329 23523 19363
rect 27169 19329 27203 19363
rect 27353 19329 27387 19363
rect 33333 19329 33367 19363
rect 38945 19329 38979 19363
rect 41337 19329 41371 19363
rect 42901 19329 42935 19363
rect 42993 19329 43027 19363
rect 15669 19261 15703 19295
rect 20821 19261 20855 19295
rect 26985 19261 27019 19295
rect 30205 19261 30239 19295
rect 20453 19193 20487 19227
rect 21833 19193 21867 19227
rect 19349 19125 19383 19159
rect 22201 19125 22235 19159
rect 22385 19125 22419 19159
rect 24869 19125 24903 19159
rect 31585 19125 31619 19159
rect 34713 19125 34747 19159
rect 38761 19125 38795 19159
rect 43821 19125 43855 19159
rect 17141 18921 17175 18955
rect 18521 18921 18555 18955
rect 25835 18921 25869 18955
rect 25973 18853 26007 18887
rect 15485 18785 15519 18819
rect 17325 18785 17359 18819
rect 21649 18785 21683 18819
rect 21925 18785 21959 18819
rect 34805 18785 34839 18819
rect 35265 18785 35299 18819
rect 42717 18785 42751 18819
rect 44189 18785 44223 18819
rect 2053 18717 2087 18751
rect 12725 18717 12759 18751
rect 15218 18717 15252 18751
rect 15945 18717 15979 18751
rect 16129 18717 16163 18751
rect 17141 18717 17175 18751
rect 17417 18717 17451 18751
rect 18337 18717 18371 18751
rect 18613 18717 18647 18751
rect 23029 18717 23063 18751
rect 25697 18717 25731 18751
rect 26157 18717 26191 18751
rect 26801 18717 26835 18751
rect 26985 18717 27019 18751
rect 28365 18717 28399 18751
rect 31217 18717 31251 18751
rect 31473 18717 31507 18751
rect 34897 18717 34931 18751
rect 36829 18717 36863 18751
rect 36921 18717 36955 18751
rect 37473 18717 37507 18751
rect 37657 18717 37691 18751
rect 38301 18717 38335 18751
rect 12173 18649 12207 18683
rect 28549 18649 28583 18683
rect 29929 18649 29963 18683
rect 30113 18649 30147 18683
rect 44005 18649 44039 18683
rect 14105 18581 14139 18615
rect 16037 18581 16071 18615
rect 17601 18581 17635 18615
rect 18061 18581 18095 18615
rect 23213 18581 23247 18615
rect 26157 18581 26191 18615
rect 27813 18581 27847 18615
rect 32597 18581 32631 18615
rect 36645 18581 36679 18615
rect 37565 18581 37599 18615
rect 38393 18581 38427 18615
rect 43453 18377 43487 18411
rect 16833 18309 16867 18343
rect 17049 18309 17083 18343
rect 18521 18309 18555 18343
rect 25136 18309 25170 18343
rect 27537 18309 27571 18343
rect 28632 18309 28666 18343
rect 34897 18309 34931 18343
rect 38393 18309 38427 18343
rect 2053 18241 2087 18275
rect 13829 18241 13863 18275
rect 14013 18241 14047 18275
rect 14657 18241 14691 18275
rect 14749 18241 14783 18275
rect 16129 18241 16163 18275
rect 17785 18241 17819 18275
rect 17969 18241 18003 18275
rect 18705 18241 18739 18275
rect 19625 18241 19659 18275
rect 20269 18241 20303 18275
rect 20453 18241 20487 18275
rect 21097 18241 21131 18275
rect 22109 18241 22143 18275
rect 23029 18241 23063 18275
rect 23285 18241 23319 18275
rect 24869 18241 24903 18275
rect 27169 18241 27203 18275
rect 30205 18241 30239 18275
rect 32965 18241 32999 18275
rect 33057 18241 33091 18275
rect 33149 18241 33183 18275
rect 34529 18241 34563 18275
rect 34677 18241 34711 18275
rect 34805 18241 34839 18275
rect 34994 18241 35028 18275
rect 36001 18241 36035 18275
rect 37289 18241 37323 18275
rect 37473 18241 37507 18275
rect 43361 18241 43395 18275
rect 2237 18173 2271 18207
rect 2973 18173 3007 18207
rect 15853 18173 15887 18207
rect 18061 18173 18095 18207
rect 18889 18173 18923 18207
rect 19349 18173 19383 18207
rect 19533 18173 19567 18207
rect 20913 18173 20947 18207
rect 21833 18173 21867 18207
rect 26985 18173 27019 18207
rect 28365 18173 28399 18207
rect 30481 18173 30515 18207
rect 33333 18173 33367 18207
rect 35909 18173 35943 18207
rect 38209 18173 38243 18207
rect 39957 18173 39991 18207
rect 14013 18105 14047 18139
rect 20453 18105 20487 18139
rect 26249 18105 26283 18139
rect 14473 18037 14507 18071
rect 16681 18037 16715 18071
rect 16874 18037 16908 18071
rect 17601 18037 17635 18071
rect 19441 18037 19475 18071
rect 21281 18037 21315 18071
rect 21925 18037 21959 18071
rect 22293 18037 22327 18071
rect 24409 18037 24443 18071
rect 27445 18037 27479 18071
rect 29745 18037 29779 18071
rect 30297 18037 30331 18071
rect 30389 18037 30423 18071
rect 35173 18037 35207 18071
rect 36277 18037 36311 18071
rect 37473 18037 37507 18071
rect 2881 17833 2915 17867
rect 17601 17833 17635 17867
rect 22201 17833 22235 17867
rect 26249 17833 26283 17867
rect 26801 17833 26835 17867
rect 27905 17833 27939 17867
rect 30941 17833 30975 17867
rect 36185 17833 36219 17867
rect 25881 17765 25915 17799
rect 32229 17765 32263 17799
rect 15485 17697 15519 17731
rect 26249 17697 26283 17731
rect 26893 17697 26927 17731
rect 29561 17697 29595 17731
rect 32781 17697 32815 17731
rect 32965 17697 32999 17731
rect 34805 17697 34839 17731
rect 36921 17697 36955 17731
rect 37381 17697 37415 17731
rect 42349 17697 42383 17731
rect 42533 17697 42567 17731
rect 43085 17697 43119 17731
rect 1869 17629 1903 17663
rect 2973 17629 3007 17663
rect 15945 17629 15979 17663
rect 16221 17629 16255 17663
rect 17601 17629 17635 17663
rect 17693 17629 17727 17663
rect 19257 17629 19291 17663
rect 19533 17629 19567 17663
rect 19717 17629 19751 17663
rect 20821 17629 20855 17663
rect 26065 17629 26099 17663
rect 26801 17629 26835 17663
rect 28549 17629 28583 17663
rect 28733 17629 28767 17663
rect 32045 17629 32079 17663
rect 33241 17629 33275 17663
rect 34897 17629 34931 17663
rect 35265 17629 35299 17663
rect 35725 17629 35759 17663
rect 35817 17629 35851 17663
rect 36001 17629 36035 17663
rect 37013 17629 37047 17663
rect 15218 17561 15252 17595
rect 21066 17561 21100 17595
rect 26341 17561 26375 17595
rect 28089 17561 28123 17595
rect 29806 17561 29840 17595
rect 33149 17561 33183 17595
rect 35173 17561 35207 17595
rect 14105 17493 14139 17527
rect 17969 17493 18003 17527
rect 19349 17493 19383 17527
rect 27169 17493 27203 17527
rect 27721 17493 27755 17527
rect 27889 17493 27923 17527
rect 28733 17493 28767 17527
rect 15301 17289 15335 17323
rect 24869 17289 24903 17323
rect 29929 17289 29963 17323
rect 30573 17289 30607 17323
rect 14749 17221 14783 17255
rect 17049 17221 17083 17255
rect 23756 17221 23790 17255
rect 25329 17221 25363 17255
rect 25513 17221 25547 17255
rect 35817 17221 35851 17255
rect 1777 17153 1811 17187
rect 14657 17153 14691 17187
rect 14841 17153 14875 17187
rect 15577 17153 15611 17187
rect 15669 17153 15703 17187
rect 15761 17153 15795 17187
rect 15945 17153 15979 17187
rect 16865 17153 16899 17187
rect 16957 17153 16991 17187
rect 17233 17153 17267 17187
rect 17693 17153 17727 17187
rect 17785 17153 17819 17187
rect 19441 17153 19475 17187
rect 19625 17153 19659 17187
rect 20453 17153 20487 17187
rect 21833 17153 21867 17187
rect 22017 17153 22051 17187
rect 26065 17153 26099 17187
rect 27169 17153 27203 17187
rect 28816 17153 28850 17187
rect 30481 17153 30515 17187
rect 32873 17153 32907 17187
rect 33057 17153 33091 17187
rect 37289 17153 37323 17187
rect 37473 17153 37507 17187
rect 43361 17153 43395 17187
rect 1961 17085 1995 17119
rect 2789 17085 2823 17119
rect 18153 17085 18187 17119
rect 19349 17085 19383 17119
rect 20269 17085 20303 17119
rect 23489 17085 23523 17119
rect 27077 17085 27111 17119
rect 28549 17085 28583 17119
rect 36277 17085 36311 17119
rect 16681 17017 16715 17051
rect 19809 17017 19843 17051
rect 26249 17017 26283 17051
rect 27537 17017 27571 17051
rect 36093 17017 36127 17051
rect 17969 16949 18003 16983
rect 20637 16949 20671 16983
rect 22017 16949 22051 16983
rect 32965 16949 32999 16983
rect 37657 16949 37691 16983
rect 43453 16949 43487 16983
rect 44189 16949 44223 16983
rect 2329 16745 2363 16779
rect 15761 16745 15795 16779
rect 23121 16745 23155 16779
rect 20821 16677 20855 16711
rect 22753 16677 22787 16711
rect 32413 16677 32447 16711
rect 37105 16677 37139 16711
rect 15301 16609 15335 16643
rect 15393 16609 15427 16643
rect 15485 16609 15519 16643
rect 17325 16609 17359 16643
rect 19533 16609 19567 16643
rect 21465 16609 21499 16643
rect 24869 16609 24903 16643
rect 31033 16609 31067 16643
rect 33793 16609 33827 16643
rect 33885 16609 33919 16643
rect 34069 16609 34103 16643
rect 34989 16609 35023 16643
rect 37657 16609 37691 16643
rect 44005 16609 44039 16643
rect 44189 16609 44223 16643
rect 1777 16541 1811 16575
rect 2421 16541 2455 16575
rect 13461 16541 13495 16575
rect 15577 16541 15611 16575
rect 16221 16541 16255 16575
rect 16405 16541 16439 16575
rect 16497 16541 16531 16575
rect 16589 16541 16623 16575
rect 19257 16541 19291 16575
rect 21649 16541 21683 16575
rect 24409 16541 24443 16575
rect 24685 16541 24719 16575
rect 31289 16541 31323 16575
rect 36737 16541 36771 16575
rect 37933 16541 37967 16575
rect 42349 16541 42383 16575
rect 16865 16473 16899 16507
rect 17570 16473 17604 16507
rect 20545 16473 20579 16507
rect 23121 16473 23155 16507
rect 35817 16473 35851 16507
rect 13277 16405 13311 16439
rect 18705 16405 18739 16439
rect 21005 16405 21039 16439
rect 23305 16405 23339 16439
rect 24501 16405 24535 16439
rect 33425 16405 33459 16439
rect 37197 16405 37231 16439
rect 17877 16201 17911 16235
rect 22293 16201 22327 16235
rect 23489 16201 23523 16235
rect 33241 16201 33275 16235
rect 33885 16201 33919 16235
rect 19533 16133 19567 16167
rect 23305 16133 23339 16167
rect 28816 16133 28850 16167
rect 32873 16133 32907 16167
rect 33057 16133 33091 16167
rect 1685 16065 1719 16099
rect 12909 16065 12943 16099
rect 15761 16065 15795 16099
rect 15945 16065 15979 16099
rect 16911 16065 16945 16099
rect 17049 16065 17083 16099
rect 17141 16068 17175 16102
rect 17325 16065 17359 16099
rect 17877 16065 17911 16099
rect 18153 16065 18187 16099
rect 20269 16065 20303 16099
rect 20453 16065 20487 16099
rect 21833 16065 21867 16099
rect 22109 16065 22143 16099
rect 24205 16065 24239 16099
rect 26985 16065 27019 16099
rect 27169 16065 27203 16099
rect 27813 16065 27847 16099
rect 28549 16065 28583 16099
rect 33701 16065 33735 16099
rect 33885 16065 33919 16099
rect 36553 16065 36587 16099
rect 36737 16065 36771 16099
rect 37749 16065 37783 16099
rect 38117 16065 38151 16099
rect 43361 16065 43395 16099
rect 1869 15997 1903 16031
rect 2789 15997 2823 16031
rect 13093 15997 13127 16031
rect 14749 15997 14783 16031
rect 15669 15997 15703 16031
rect 15853 15997 15887 16031
rect 20177 15997 20211 16031
rect 20637 15997 20671 16031
rect 23949 15997 23983 16031
rect 19349 15929 19383 15963
rect 22937 15929 22971 15963
rect 25329 15929 25363 15963
rect 37565 15929 37599 15963
rect 16129 15861 16163 15895
rect 16681 15861 16715 15895
rect 21925 15861 21959 15895
rect 23305 15861 23339 15895
rect 27169 15861 27203 15895
rect 27629 15861 27663 15895
rect 29929 15861 29963 15895
rect 36737 15861 36771 15895
rect 37933 15861 37967 15895
rect 42717 15861 42751 15895
rect 43453 15861 43487 15895
rect 44189 15861 44223 15895
rect 2237 15657 2271 15691
rect 13185 15657 13219 15691
rect 15301 15657 15335 15691
rect 17233 15657 17267 15691
rect 19717 15657 19751 15691
rect 20545 15657 20579 15691
rect 21189 15657 21223 15691
rect 22201 15657 22235 15691
rect 22569 15657 22603 15691
rect 26525 15657 26559 15691
rect 23121 15589 23155 15623
rect 36093 15589 36127 15623
rect 16681 15521 16715 15555
rect 21097 15521 21131 15555
rect 23305 15521 23339 15555
rect 37657 15521 37691 15555
rect 42625 15521 42659 15555
rect 44189 15521 44223 15555
rect 2329 15453 2363 15487
rect 13277 15453 13311 15487
rect 16425 15453 16459 15487
rect 17325 15453 17359 15487
rect 20361 15453 20395 15487
rect 20545 15453 20579 15487
rect 21373 15453 21407 15487
rect 22201 15453 22235 15487
rect 22293 15453 22327 15487
rect 23029 15453 23063 15487
rect 24409 15453 24443 15487
rect 27905 15453 27939 15487
rect 29653 15453 29687 15487
rect 30941 15453 30975 15487
rect 31208 15453 31242 15487
rect 32781 15453 32815 15487
rect 32965 15453 32999 15487
rect 33609 15453 33643 15487
rect 33793 15453 33827 15487
rect 36093 15453 36127 15487
rect 36277 15453 36311 15487
rect 36369 15453 36403 15487
rect 37933 15453 37967 15487
rect 38945 15453 38979 15487
rect 19809 15385 19843 15419
rect 21557 15385 21591 15419
rect 24654 15385 24688 15419
rect 27638 15385 27672 15419
rect 37013 15385 37047 15419
rect 37197 15385 37231 15419
rect 44005 15385 44039 15419
rect 23305 15317 23339 15351
rect 25789 15317 25823 15351
rect 29745 15317 29779 15351
rect 32321 15317 32355 15351
rect 33149 15317 33183 15351
rect 33701 15317 33735 15351
rect 36829 15317 36863 15351
rect 39037 15317 39071 15351
rect 17509 15113 17543 15147
rect 17677 15113 17711 15147
rect 25513 15113 25547 15147
rect 30573 15113 30607 15147
rect 35357 15113 35391 15147
rect 39497 15113 39531 15147
rect 43453 15113 43487 15147
rect 17877 15045 17911 15079
rect 23305 15045 23339 15079
rect 23949 15045 23983 15079
rect 25421 15045 25455 15079
rect 30757 15045 30791 15079
rect 36579 15045 36613 15079
rect 39129 15045 39163 15079
rect 13369 14977 13403 15011
rect 18521 14977 18555 15011
rect 19533 14977 19567 15011
rect 20821 14977 20855 15011
rect 21005 14977 21039 15011
rect 21833 14977 21867 15011
rect 23121 14977 23155 15011
rect 26249 14977 26283 15011
rect 26433 14977 26467 15011
rect 27169 14977 27203 15011
rect 28089 14977 28123 15011
rect 29000 14977 29034 15011
rect 32229 14977 32263 15011
rect 32413 14977 32447 15011
rect 32689 14977 32723 15011
rect 33609 14977 33643 15011
rect 33885 14977 33919 15011
rect 35265 14977 35299 15011
rect 36277 14977 36311 15011
rect 36369 14977 36403 15011
rect 36461 14977 36495 15011
rect 36737 14977 36771 15011
rect 38853 14977 38887 15011
rect 38946 14977 38980 15011
rect 39221 14977 39255 15011
rect 39318 14977 39352 15011
rect 43361 14977 43395 15011
rect 18705 14909 18739 14943
rect 19257 14909 19291 14943
rect 22109 14909 22143 14943
rect 27077 14909 27111 14943
rect 28733 14909 28767 14943
rect 34253 14909 34287 14943
rect 35541 14909 35575 14943
rect 37565 14909 37599 14943
rect 37841 14909 37875 14943
rect 24133 14841 24167 14875
rect 28273 14841 28307 14875
rect 31125 14841 31159 14875
rect 13461 14773 13495 14807
rect 17693 14773 17727 14807
rect 18337 14773 18371 14807
rect 19349 14773 19383 14807
rect 19717 14773 19751 14807
rect 20913 14773 20947 14807
rect 26341 14773 26375 14807
rect 27537 14773 27571 14807
rect 30113 14773 30147 14807
rect 30757 14773 30791 14807
rect 32413 14773 32447 14807
rect 34897 14773 34931 14807
rect 36093 14773 36127 14807
rect 18245 14569 18279 14603
rect 21833 14569 21867 14603
rect 22845 14569 22879 14603
rect 25973 14569 26007 14603
rect 27077 14569 27111 14603
rect 27445 14569 27479 14603
rect 30021 14569 30055 14603
rect 30205 14569 30239 14603
rect 36185 14569 36219 14603
rect 21005 14501 21039 14535
rect 26157 14501 26191 14535
rect 38025 14501 38059 14535
rect 38577 14501 38611 14535
rect 14289 14433 14323 14467
rect 25789 14433 25823 14467
rect 29929 14433 29963 14467
rect 31217 14433 31251 14467
rect 31677 14433 31711 14467
rect 32597 14433 32631 14467
rect 35541 14433 35575 14467
rect 36737 14433 36771 14467
rect 37381 14433 37415 14467
rect 37749 14433 37783 14467
rect 37841 14433 37875 14467
rect 42349 14433 42383 14467
rect 44097 14433 44131 14467
rect 2145 14365 2179 14399
rect 3065 14365 3099 14399
rect 14105 14365 14139 14399
rect 17877 14365 17911 14399
rect 18061 14365 18095 14399
rect 18337 14365 18371 14399
rect 19625 14365 19659 14399
rect 19881 14365 19915 14399
rect 22569 14365 22603 14399
rect 22661 14365 22695 14399
rect 23673 14365 23707 14399
rect 25973 14365 26007 14399
rect 26985 14365 27019 14399
rect 30021 14365 30055 14399
rect 31309 14365 31343 14399
rect 32689 14365 32723 14399
rect 33977 14365 34011 14399
rect 34161 14365 34195 14399
rect 35357 14365 35391 14399
rect 36645 14365 36679 14399
rect 38477 14365 38511 14399
rect 38669 14365 38703 14399
rect 15945 14297 15979 14331
rect 21817 14297 21851 14331
rect 22017 14297 22051 14331
rect 23489 14297 23523 14331
rect 25697 14297 25731 14331
rect 29745 14297 29779 14331
rect 34069 14297 34103 14331
rect 35449 14297 35483 14331
rect 42533 14297 42567 14331
rect 2973 14229 3007 14263
rect 21649 14229 21683 14263
rect 23305 14229 23339 14263
rect 33517 14229 33551 14263
rect 34989 14229 35023 14263
rect 36553 14229 36587 14263
rect 14013 14025 14047 14059
rect 20361 14025 20395 14059
rect 21189 14025 21223 14059
rect 23581 14025 23615 14059
rect 26157 14025 26191 14059
rect 29653 14025 29687 14059
rect 30113 14025 30147 14059
rect 32321 14025 32355 14059
rect 34345 14025 34379 14059
rect 34437 14025 34471 14059
rect 37457 14025 37491 14059
rect 2237 13957 2271 13991
rect 20177 13957 20211 13991
rect 20821 13957 20855 13991
rect 27721 13957 27755 13991
rect 37657 13957 37691 13991
rect 38853 13957 38887 13991
rect 2053 13889 2087 13923
rect 13829 13889 13863 13923
rect 16681 13889 16715 13923
rect 16948 13889 16982 13923
rect 19809 13889 19843 13923
rect 21005 13889 21039 13923
rect 21281 13889 21315 13923
rect 22201 13889 22235 13923
rect 22457 13889 22491 13923
rect 26341 13889 26375 13923
rect 28273 13889 28307 13923
rect 28540 13889 28574 13923
rect 31226 13889 31260 13923
rect 32229 13889 32263 13923
rect 32413 13889 32447 13923
rect 35725 13889 35759 13923
rect 38209 13889 38243 13923
rect 39129 13889 39163 13923
rect 39589 13889 39623 13923
rect 39773 13889 39807 13923
rect 43637 13889 43671 13923
rect 2789 13821 2823 13855
rect 19073 13821 19107 13855
rect 19349 13821 19383 13855
rect 31493 13821 31527 13855
rect 34529 13821 34563 13855
rect 36001 13821 36035 13855
rect 38853 13821 38887 13855
rect 18061 13753 18095 13787
rect 27537 13753 27571 13787
rect 39037 13753 39071 13787
rect 20177 13685 20211 13719
rect 33977 13685 34011 13719
rect 37289 13685 37323 13719
rect 37473 13685 37507 13719
rect 38301 13685 38335 13719
rect 39681 13685 39715 13719
rect 42809 13685 42843 13719
rect 43545 13685 43579 13719
rect 16865 13481 16899 13515
rect 18061 13481 18095 13515
rect 18521 13481 18555 13515
rect 21373 13481 21407 13515
rect 25789 13481 25823 13515
rect 36737 13481 36771 13515
rect 38945 13481 38979 13515
rect 17325 13413 17359 13447
rect 18429 13345 18463 13379
rect 21833 13345 21867 13379
rect 23029 13345 23063 13379
rect 36553 13345 36587 13379
rect 42349 13345 42383 13379
rect 44097 13345 44131 13379
rect 1777 13277 1811 13311
rect 16681 13277 16715 13311
rect 18245 13277 18279 13311
rect 19717 13277 19751 13311
rect 19993 13277 20027 13311
rect 21097 13277 21131 13311
rect 22017 13277 22051 13311
rect 22109 13277 22143 13311
rect 22753 13277 22787 13311
rect 24409 13277 24443 13311
rect 32505 13277 32539 13311
rect 36829 13277 36863 13311
rect 37473 13277 37507 13311
rect 37657 13277 37691 13311
rect 37749 13277 37783 13311
rect 37841 13277 37875 13311
rect 17509 13209 17543 13243
rect 18521 13209 18555 13243
rect 21373 13209 21407 13243
rect 21833 13209 21867 13243
rect 24676 13209 24710 13243
rect 38577 13209 38611 13243
rect 38761 13209 38795 13243
rect 42533 13209 42567 13243
rect 21189 13141 21223 13175
rect 32689 13141 32723 13175
rect 36277 13141 36311 13175
rect 38117 13141 38151 13175
rect 18337 12937 18371 12971
rect 19533 12937 19567 12971
rect 21281 12937 21315 12971
rect 23857 12937 23891 12971
rect 25789 12937 25823 12971
rect 27169 12937 27203 12971
rect 36093 12937 36127 12971
rect 39129 12937 39163 12971
rect 18705 12869 18739 12903
rect 20913 12869 20947 12903
rect 21129 12869 21163 12903
rect 21833 12869 21867 12903
rect 27261 12869 27295 12903
rect 31033 12869 31067 12903
rect 31217 12869 31251 12903
rect 41705 12869 41739 12903
rect 43545 12869 43579 12903
rect 1685 12801 1719 12835
rect 9229 12801 9263 12835
rect 18521 12801 18555 12835
rect 19717 12801 19751 12835
rect 19901 12801 19935 12835
rect 22017 12801 22051 12835
rect 22201 12801 22235 12835
rect 22293 12801 22327 12835
rect 22937 12801 22971 12835
rect 23673 12801 23707 12835
rect 24665 12801 24699 12835
rect 27813 12801 27847 12835
rect 27997 12801 28031 12835
rect 28181 12801 28215 12835
rect 28641 12801 28675 12835
rect 29837 12801 29871 12835
rect 33250 12801 33284 12835
rect 33517 12801 33551 12835
rect 35633 12801 35667 12835
rect 38301 12801 38335 12835
rect 39037 12801 39071 12835
rect 39221 12801 39255 12835
rect 43637 12801 43671 12835
rect 1869 12733 1903 12767
rect 2789 12733 2823 12767
rect 24409 12733 24443 12767
rect 35725 12733 35759 12767
rect 38577 12733 38611 12767
rect 41337 12733 41371 12767
rect 41889 12733 41923 12767
rect 42809 12733 42843 12767
rect 9321 12597 9355 12631
rect 21097 12597 21131 12631
rect 22753 12597 22787 12631
rect 28825 12597 28859 12631
rect 30481 12597 30515 12631
rect 32137 12597 32171 12631
rect 35449 12597 35483 12631
rect 2237 12393 2271 12427
rect 18429 12393 18463 12427
rect 21557 12393 21591 12427
rect 23857 12393 23891 12427
rect 19901 12257 19935 12291
rect 20177 12257 20211 12291
rect 24593 12257 24627 12291
rect 32229 12257 32263 12291
rect 32321 12257 32355 12291
rect 35357 12257 35391 12291
rect 36461 12257 36495 12291
rect 37841 12257 37875 12291
rect 38025 12257 38059 12291
rect 42717 12257 42751 12291
rect 2329 12189 2363 12223
rect 18153 12189 18187 12223
rect 22670 12189 22704 12223
rect 22937 12189 22971 12223
rect 23673 12189 23707 12223
rect 24777 12189 24811 12223
rect 25421 12189 25455 12223
rect 27261 12189 27295 12223
rect 27528 12189 27562 12223
rect 29653 12189 29687 12223
rect 33333 12189 33367 12223
rect 33977 12189 34011 12223
rect 35173 12189 35207 12223
rect 38577 12189 38611 12223
rect 38761 12189 38795 12223
rect 44189 12189 44223 12223
rect 18429 12121 18463 12155
rect 25688 12121 25722 12155
rect 29920 12121 29954 12155
rect 37749 12121 37783 12155
rect 44005 12121 44039 12155
rect 18245 12053 18279 12087
rect 24961 12053 24995 12087
rect 26801 12053 26835 12087
rect 31033 12053 31067 12087
rect 31769 12053 31803 12087
rect 32137 12053 32171 12087
rect 33149 12053 33183 12087
rect 33793 12053 33827 12087
rect 34713 12053 34747 12087
rect 35081 12053 35115 12087
rect 35909 12053 35943 12087
rect 36277 12053 36311 12087
rect 36369 12053 36403 12087
rect 37381 12053 37415 12087
rect 38669 12053 38703 12087
rect 24593 11849 24627 11883
rect 25697 11849 25731 11883
rect 29837 11849 29871 11883
rect 30849 11849 30883 11883
rect 31217 11849 31251 11883
rect 32137 11849 32171 11883
rect 34345 11849 34379 11883
rect 35541 11849 35575 11883
rect 35725 11849 35759 11883
rect 37289 11849 37323 11883
rect 43453 11849 43487 11883
rect 20269 11781 20303 11815
rect 28724 11781 28758 11815
rect 33250 11781 33284 11815
rect 34805 11781 34839 11815
rect 37381 11781 37415 11815
rect 37565 11781 37599 11815
rect 38025 11781 38059 11815
rect 17224 11713 17258 11747
rect 20637 11713 20671 11747
rect 23765 11713 23799 11747
rect 24409 11713 24443 11747
rect 25053 11713 25087 11747
rect 25881 11713 25915 11747
rect 28457 11713 28491 11747
rect 33517 11713 33551 11747
rect 34713 11713 34747 11747
rect 35722 11713 35756 11747
rect 37291 11713 37325 11747
rect 38209 11713 38243 11747
rect 38301 11713 38335 11747
rect 43361 11713 43395 11747
rect 44189 11713 44223 11747
rect 16957 11645 16991 11679
rect 18797 11645 18831 11679
rect 19073 11645 19107 11679
rect 31309 11645 31343 11679
rect 31401 11645 31435 11679
rect 34989 11645 35023 11679
rect 36185 11645 36219 11679
rect 18337 11577 18371 11611
rect 38025 11577 38059 11611
rect 20085 11509 20119 11543
rect 20269 11509 20303 11543
rect 23949 11509 23983 11543
rect 25237 11509 25271 11543
rect 36093 11509 36127 11543
rect 18521 11305 18555 11339
rect 18705 11305 18739 11339
rect 21649 11305 21683 11339
rect 23673 11305 23707 11339
rect 24777 11305 24811 11339
rect 27169 11305 27203 11339
rect 27353 11305 27387 11339
rect 31861 11305 31895 11339
rect 35265 11305 35299 11339
rect 26709 11237 26743 11271
rect 32045 11237 32079 11271
rect 32781 11237 32815 11271
rect 17601 11169 17635 11203
rect 20269 11169 20303 11203
rect 23305 11169 23339 11203
rect 27537 11169 27571 11203
rect 36369 11169 36403 11203
rect 43729 11169 43763 11203
rect 2053 11101 2087 11135
rect 17785 11101 17819 11135
rect 17877 11101 17911 11135
rect 19625 11101 19659 11135
rect 23489 11101 23523 11135
rect 24409 11101 24443 11135
rect 24593 11101 24627 11135
rect 25329 11101 25363 11135
rect 25585 11101 25619 11135
rect 27353 11101 27387 11135
rect 28273 11101 28307 11135
rect 30205 11101 30239 11135
rect 34161 11101 34195 11135
rect 35449 11101 35483 11135
rect 35725 11101 35759 11135
rect 35909 11101 35943 11135
rect 44189 11101 44223 11135
rect 18337 11033 18371 11067
rect 20514 11033 20548 11067
rect 27629 11033 27663 11067
rect 28089 11033 28123 11067
rect 32321 11033 32355 11067
rect 33894 11033 33928 11067
rect 36553 11033 36587 11067
rect 36737 11033 36771 11067
rect 44005 11033 44039 11067
rect 17601 10965 17635 10999
rect 18537 10965 18571 10999
rect 19809 10965 19843 10999
rect 28457 10965 28491 10999
rect 30849 10965 30883 10999
rect 17693 10761 17727 10795
rect 20453 10761 20487 10795
rect 23673 10761 23707 10795
rect 26433 10761 26467 10795
rect 28365 10761 28399 10795
rect 30205 10761 30239 10795
rect 43453 10761 43487 10795
rect 17509 10693 17543 10727
rect 29070 10693 29104 10727
rect 2605 10625 2639 10659
rect 17785 10625 17819 10659
rect 18337 10625 18371 10659
rect 18521 10625 18555 10659
rect 20637 10625 20671 10659
rect 20729 10625 20763 10659
rect 23489 10625 23523 10659
rect 24225 10625 24259 10659
rect 24317 10625 24351 10659
rect 25309 10625 25343 10659
rect 28181 10625 28215 10659
rect 28825 10625 28859 10659
rect 43361 10625 43395 10659
rect 44189 10625 44223 10659
rect 18705 10557 18739 10591
rect 20821 10557 20855 10591
rect 20913 10557 20947 10591
rect 23305 10557 23339 10591
rect 25053 10557 25087 10591
rect 17509 10489 17543 10523
rect 1961 10421 1995 10455
rect 2513 10421 2547 10455
rect 24501 10421 24535 10455
rect 18705 10217 18739 10251
rect 22293 10217 22327 10251
rect 22937 10217 22971 10251
rect 23121 10217 23155 10251
rect 31677 10217 31711 10251
rect 20821 10149 20855 10183
rect 21925 10149 21959 10183
rect 22477 10149 22511 10183
rect 1409 10081 1443 10115
rect 3249 10081 3283 10115
rect 17325 10081 17359 10115
rect 19625 10081 19659 10115
rect 24409 10081 24443 10115
rect 30297 10081 30331 10115
rect 3985 10013 4019 10047
rect 19809 10013 19843 10047
rect 19901 10013 19935 10047
rect 24593 10013 24627 10047
rect 25237 10013 25271 10047
rect 27445 10013 27479 10047
rect 30564 10013 30598 10047
rect 3065 9945 3099 9979
rect 3893 9945 3927 9979
rect 17592 9945 17626 9979
rect 20545 9945 20579 9979
rect 23305 9945 23339 9979
rect 25504 9945 25538 9979
rect 27690 9945 27724 9979
rect 19625 9877 19659 9911
rect 21005 9877 21039 9911
rect 22293 9877 22327 9911
rect 23105 9877 23139 9911
rect 24777 9877 24811 9911
rect 26617 9877 26651 9911
rect 17693 9673 17727 9707
rect 24961 9673 24995 9707
rect 25605 9673 25639 9707
rect 17601 9537 17635 9571
rect 17785 9537 17819 9571
rect 18429 9537 18463 9571
rect 18521 9537 18555 9571
rect 19349 9537 19383 9571
rect 19616 9537 19650 9571
rect 22385 9537 22419 9571
rect 23673 9537 23707 9571
rect 24777 9537 24811 9571
rect 25421 9537 25455 9571
rect 42809 9537 42843 9571
rect 1961 9469 1995 9503
rect 2145 9469 2179 9503
rect 2789 9469 2823 9503
rect 18245 9469 18279 9503
rect 22661 9469 22695 9503
rect 18337 9401 18371 9435
rect 20729 9401 20763 9435
rect 23857 9333 23891 9367
rect 42901 9333 42935 9367
rect 1961 9129 1995 9163
rect 2513 9129 2547 9163
rect 19625 9129 19659 9163
rect 22753 9129 22787 9163
rect 42533 8993 42567 9027
rect 2605 8925 2639 8959
rect 19625 8925 19659 8959
rect 19901 8925 19935 8959
rect 20913 8925 20947 8959
rect 22937 8925 22971 8959
rect 23213 8925 23247 8959
rect 42349 8925 42383 8959
rect 19809 8857 19843 8891
rect 21180 8857 21214 8891
rect 23121 8857 23155 8891
rect 44189 8857 44223 8891
rect 22293 8789 22327 8823
rect 21189 8585 21223 8619
rect 22753 8585 22787 8619
rect 2145 8517 2179 8551
rect 23866 8517 23900 8551
rect 1961 8449 1995 8483
rect 21005 8449 21039 8483
rect 24133 8449 24167 8483
rect 43637 8449 43671 8483
rect 2881 8381 2915 8415
rect 44189 7837 44223 7871
rect 44005 7701 44039 7735
rect 3433 7361 3467 7395
rect 43545 7361 43579 7395
rect 3525 7157 3559 7191
rect 4077 7157 4111 7191
rect 43637 7157 43671 7191
rect 3801 6817 3835 6851
rect 4721 6817 4755 6851
rect 42717 6817 42751 6851
rect 44005 6817 44039 6851
rect 1777 6749 1811 6783
rect 44189 6749 44223 6783
rect 3985 6681 4019 6715
rect 1685 6273 1719 6307
rect 43821 6273 43855 6307
rect 1869 6205 1903 6239
rect 2789 6205 2823 6239
rect 2145 5865 2179 5899
rect 42717 5729 42751 5763
rect 1593 5661 1627 5695
rect 2237 5661 2271 5695
rect 2973 5661 3007 5695
rect 3801 5661 3835 5695
rect 4445 5661 4479 5695
rect 44189 5661 44223 5695
rect 44005 5593 44039 5627
rect 2881 5525 2915 5559
rect 2145 5253 2179 5287
rect 1961 5185 1995 5219
rect 4445 5185 4479 5219
rect 42809 5185 42843 5219
rect 2789 5117 2823 5151
rect 4353 4981 4387 5015
rect 4905 4981 4939 5015
rect 42901 4981 42935 5015
rect 43637 4981 43671 5015
rect 1961 4641 1995 4675
rect 4077 4641 4111 4675
rect 4261 4641 4295 4675
rect 4813 4641 4847 4675
rect 38025 4641 38059 4675
rect 42349 4641 42383 4675
rect 42533 4641 42567 4675
rect 44097 4641 44131 4675
rect 2605 4573 2639 4607
rect 3249 4573 3283 4607
rect 6377 4573 6411 4607
rect 37381 4573 37415 4607
rect 37565 4505 37599 4539
rect 3157 4437 3191 4471
rect 2053 4097 2087 4131
rect 4353 4097 4387 4131
rect 5365 4097 5399 4131
rect 11805 4097 11839 4131
rect 21005 4097 21039 4131
rect 36553 4097 36587 4131
rect 37933 4097 37967 4131
rect 41705 4097 41739 4131
rect 43361 4097 43395 4131
rect 2789 4029 2823 4063
rect 4169 4029 4203 4063
rect 38853 4029 38887 4063
rect 39037 4029 39071 4063
rect 40693 4029 40727 4063
rect 36645 3961 36679 3995
rect 1961 3893 1995 3927
rect 5457 3893 5491 3927
rect 6377 3893 6411 3927
rect 7389 3893 7423 3927
rect 9321 3893 9355 3927
rect 11897 3893 11931 3927
rect 12449 3893 12483 3927
rect 15577 3893 15611 3927
rect 20913 3893 20947 3927
rect 24225 3893 24259 3927
rect 37289 3893 37323 3927
rect 41797 3893 41831 3927
rect 42441 3893 42475 3927
rect 43453 3893 43487 3927
rect 44005 3893 44039 3927
rect 38301 3689 38335 3723
rect 38853 3689 38887 3723
rect 44097 3689 44131 3723
rect 3249 3553 3283 3587
rect 5365 3553 5399 3587
rect 5549 3553 5583 3587
rect 5825 3553 5859 3587
rect 9229 3553 9263 3587
rect 9413 3553 9447 3587
rect 9689 3553 9723 3587
rect 15485 3553 15519 3587
rect 16129 3553 16163 3587
rect 20821 3553 20855 3587
rect 21281 3553 21315 3587
rect 35817 3553 35851 3587
rect 36093 3553 36127 3587
rect 41705 3553 41739 3587
rect 41889 3553 41923 3587
rect 42533 3553 42567 3587
rect 1409 3485 1443 3519
rect 4537 3485 4571 3519
rect 8309 3485 8343 3519
rect 12265 3485 12299 3519
rect 12909 3485 12943 3519
rect 17785 3485 17819 3519
rect 18705 3485 18739 3519
rect 19441 3485 19475 3519
rect 20177 3485 20211 3519
rect 20637 3485 20671 3519
rect 22937 3485 22971 3519
rect 23673 3485 23707 3519
rect 24777 3485 24811 3519
rect 25237 3485 25271 3519
rect 29009 3485 29043 3519
rect 29745 3485 29779 3519
rect 35633 3485 35667 3519
rect 38209 3485 38243 3519
rect 40049 3485 40083 3519
rect 40877 3485 40911 3519
rect 44005 3485 44039 3519
rect 3065 3417 3099 3451
rect 15669 3417 15703 3451
rect 4445 3349 4479 3383
rect 8217 3349 8251 3383
rect 12173 3349 12207 3383
rect 19349 3349 19383 3383
rect 23765 3349 23799 3383
rect 24685 3349 24719 3383
rect 29653 3349 29687 3383
rect 40785 3349 40819 3383
rect 2237 3145 2271 3179
rect 15761 3145 15795 3179
rect 36645 3145 36679 3179
rect 2973 3077 3007 3111
rect 3709 3077 3743 3111
rect 7481 3077 7515 3111
rect 13185 3077 13219 3111
rect 18981 3077 19015 3111
rect 24593 3077 24627 3111
rect 29377 3077 29411 3111
rect 2329 3009 2363 3043
rect 3065 3009 3099 3043
rect 3525 3009 3559 3043
rect 6377 3009 6411 3043
rect 7297 3009 7331 3043
rect 13369 3009 13403 3043
rect 15853 3009 15887 3043
rect 16957 3009 16991 3043
rect 18797 3009 18831 3043
rect 22109 3009 22143 3043
rect 24409 3009 24443 3043
rect 29193 3009 29227 3043
rect 35725 3009 35759 3043
rect 36553 3009 36587 3043
rect 39589 3009 39623 3043
rect 40049 3009 40083 3043
rect 42993 3009 43027 3043
rect 43821 3009 43855 3043
rect 3985 2941 4019 2975
rect 7757 2941 7791 2975
rect 11621 2941 11655 2975
rect 19349 2941 19383 2975
rect 22293 2941 22327 2975
rect 23213 2941 23247 2975
rect 25145 2941 25179 2975
rect 29653 2941 29687 2975
rect 39129 2941 39163 2975
rect 39405 2941 39439 2975
rect 40233 2941 40267 2975
rect 41245 2941 41279 2975
rect 42901 2873 42935 2907
rect 1501 2805 1535 2839
rect 6469 2805 6503 2839
rect 17049 2805 17083 2839
rect 22937 2601 22971 2635
rect 42993 2601 43027 2635
rect 1409 2465 1443 2499
rect 1593 2465 1627 2499
rect 2789 2465 2823 2499
rect 3801 2465 3835 2499
rect 3985 2465 4019 2499
rect 4721 2465 4755 2499
rect 6377 2465 6411 2499
rect 6561 2465 6595 2499
rect 6929 2465 6963 2499
rect 11713 2465 11747 2499
rect 11897 2465 11931 2499
rect 12265 2465 12299 2499
rect 16865 2465 16899 2499
rect 17049 2465 17083 2499
rect 17417 2465 17451 2499
rect 24409 2465 24443 2499
rect 24869 2465 24903 2499
rect 37289 2465 37323 2499
rect 37473 2465 37507 2499
rect 38669 2465 38703 2499
rect 41337 2465 41371 2499
rect 41705 2465 41739 2499
rect 23029 2397 23063 2431
rect 41889 2397 41923 2431
rect 24593 2329 24627 2363
<< metal1 >>
rect 23842 44072 23848 44124
rect 23900 44112 23906 44124
rect 24854 44112 24860 44124
rect 23900 44084 24860 44112
rect 23900 44072 23906 44084
rect 24854 44072 24860 44084
rect 24912 44072 24918 44124
rect 1104 43546 44896 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 44896 43546
rect 1104 43472 44896 43494
rect 6886 43404 16574 43432
rect 6886 43364 6914 43404
rect 3344 43336 6914 43364
rect 13173 43367 13231 43373
rect 3344 43308 3372 43336
rect 13173 43333 13185 43367
rect 13219 43364 13231 43367
rect 14277 43367 14335 43373
rect 14277 43364 14289 43367
rect 13219 43336 14289 43364
rect 13219 43333 13231 43336
rect 13173 43327 13231 43333
rect 14277 43333 14289 43336
rect 14323 43333 14335 43367
rect 14277 43327 14335 43333
rect 1854 43296 1860 43308
rect 1815 43268 1860 43296
rect 1854 43256 1860 43268
rect 1912 43256 1918 43308
rect 2869 43299 2927 43305
rect 2869 43265 2881 43299
rect 2915 43296 2927 43299
rect 3326 43296 3332 43308
rect 2915 43268 3332 43296
rect 2915 43265 2927 43268
rect 2869 43259 2927 43265
rect 3326 43256 3332 43268
rect 3384 43256 3390 43308
rect 7742 43256 7748 43308
rect 7800 43296 7806 43308
rect 7837 43299 7895 43305
rect 7837 43296 7849 43299
rect 7800 43268 7849 43296
rect 7800 43256 7806 43268
rect 7837 43265 7849 43268
rect 7883 43265 7895 43299
rect 12526 43296 12532 43308
rect 12487 43268 12532 43296
rect 7837 43259 7895 43265
rect 12526 43256 12532 43268
rect 12584 43256 12590 43308
rect 13078 43296 13084 43308
rect 13039 43268 13084 43296
rect 13078 43256 13084 43268
rect 13136 43256 13142 43308
rect 2133 43231 2191 43237
rect 2133 43197 2145 43231
rect 2179 43228 2191 43231
rect 3602 43228 3608 43240
rect 2179 43200 3608 43228
rect 2179 43197 2191 43200
rect 2133 43191 2191 43197
rect 3602 43188 3608 43200
rect 3660 43188 3666 43240
rect 3786 43228 3792 43240
rect 3747 43200 3792 43228
rect 3786 43188 3792 43200
rect 3844 43188 3850 43240
rect 3970 43228 3976 43240
rect 3931 43200 3976 43228
rect 3970 43188 3976 43200
rect 4028 43188 4034 43240
rect 4249 43231 4307 43237
rect 4249 43197 4261 43231
rect 4295 43197 4307 43231
rect 14090 43228 14096 43240
rect 14051 43200 14096 43228
rect 4249 43191 4307 43197
rect 2038 43120 2044 43172
rect 2096 43160 2102 43172
rect 4264 43160 4292 43191
rect 14090 43188 14096 43200
rect 14148 43188 14154 43240
rect 14553 43231 14611 43237
rect 14553 43197 14565 43231
rect 14599 43197 14611 43231
rect 14553 43191 14611 43197
rect 2096 43132 4292 43160
rect 2096 43120 2102 43132
rect 13538 43120 13544 43172
rect 13596 43160 13602 43172
rect 14568 43160 14596 43191
rect 13596 43132 14596 43160
rect 16546 43160 16574 43404
rect 23474 43324 23480 43376
rect 23532 43364 23538 43376
rect 24581 43367 24639 43373
rect 24581 43364 24593 43367
rect 23532 43336 24593 43364
rect 23532 43324 23538 43336
rect 24581 43333 24593 43336
rect 24627 43333 24639 43367
rect 24581 43327 24639 43333
rect 25774 43324 25780 43376
rect 25832 43364 25838 43376
rect 27525 43367 27583 43373
rect 27525 43364 27537 43367
rect 25832 43336 27537 43364
rect 25832 43324 25838 43336
rect 27525 43333 27537 43336
rect 27571 43333 27583 43367
rect 27525 43327 27583 43333
rect 23477 43231 23535 43237
rect 23477 43197 23489 43231
rect 23523 43228 23535 43231
rect 24397 43231 24455 43237
rect 24397 43228 24409 43231
rect 23523 43200 24409 43228
rect 23523 43197 23535 43200
rect 23477 43191 23535 43197
rect 24397 43197 24409 43200
rect 24443 43197 24455 43231
rect 24854 43228 24860 43240
rect 24815 43200 24860 43228
rect 24397 43191 24455 43197
rect 24854 43188 24860 43200
rect 24912 43188 24918 43240
rect 32309 43231 32367 43237
rect 32309 43197 32321 43231
rect 32355 43197 32367 43231
rect 32309 43191 32367 43197
rect 32493 43231 32551 43237
rect 32493 43197 32505 43231
rect 32539 43228 32551 43231
rect 33318 43228 33324 43240
rect 32539 43200 33324 43228
rect 32539 43197 32551 43200
rect 32493 43191 32551 43197
rect 32324 43160 32352 43191
rect 33318 43188 33324 43200
rect 33376 43188 33382 43240
rect 33502 43228 33508 43240
rect 33463 43200 33508 43228
rect 33502 43188 33508 43200
rect 33560 43188 33566 43240
rect 33134 43160 33140 43172
rect 16546 43132 30604 43160
rect 32324 43132 33140 43160
rect 13596 43120 13602 43132
rect 2774 43092 2780 43104
rect 2735 43064 2780 43092
rect 2774 43052 2780 43064
rect 2832 43052 2838 43104
rect 6546 43092 6552 43104
rect 6507 43064 6552 43092
rect 6546 43052 6552 43064
rect 6604 43052 6610 43104
rect 8018 43092 8024 43104
rect 7979 43064 8024 43092
rect 8018 43052 8024 43064
rect 8076 43052 8082 43104
rect 10965 43095 11023 43101
rect 10965 43061 10977 43095
rect 11011 43092 11023 43095
rect 11514 43092 11520 43104
rect 11011 43064 11520 43092
rect 11011 43061 11023 43064
rect 10965 43055 11023 43061
rect 11514 43052 11520 43064
rect 11572 43052 11578 43104
rect 11606 43052 11612 43104
rect 11664 43092 11670 43104
rect 11701 43095 11759 43101
rect 11701 43092 11713 43095
rect 11664 43064 11713 43092
rect 11664 43052 11670 43064
rect 11701 43061 11713 43064
rect 11747 43061 11759 43095
rect 12434 43092 12440 43104
rect 12395 43064 12440 43092
rect 11701 43055 11759 43061
rect 12434 43052 12440 43064
rect 12492 43052 12498 43104
rect 20806 43092 20812 43104
rect 20767 43064 20812 43092
rect 20806 43052 20812 43064
rect 20864 43052 20870 43104
rect 22646 43092 22652 43104
rect 22607 43064 22652 43092
rect 22646 43052 22652 43064
rect 22704 43052 22710 43104
rect 27154 43052 27160 43104
rect 27212 43092 27218 43104
rect 27433 43095 27491 43101
rect 27433 43092 27445 43095
rect 27212 43064 27445 43092
rect 27212 43052 27218 43064
rect 27433 43061 27445 43064
rect 27479 43061 27491 43095
rect 27433 43055 27491 43061
rect 27798 43052 27804 43104
rect 27856 43092 27862 43104
rect 28077 43095 28135 43101
rect 28077 43092 28089 43095
rect 27856 43064 28089 43092
rect 27856 43052 27862 43064
rect 28077 43061 28089 43064
rect 28123 43061 28135 43095
rect 30466 43092 30472 43104
rect 30427 43064 30472 43092
rect 28077 43055 28135 43061
rect 30466 43052 30472 43064
rect 30524 43052 30530 43104
rect 30576 43092 30604 43132
rect 33134 43120 33140 43132
rect 33192 43120 33198 43172
rect 34514 43092 34520 43104
rect 30576 43064 34520 43092
rect 34514 43052 34520 43064
rect 34572 43052 34578 43104
rect 40034 43092 40040 43104
rect 39995 43064 40040 43092
rect 40034 43052 40040 43064
rect 40092 43052 40098 43104
rect 42886 43092 42892 43104
rect 42847 43064 42892 43092
rect 42886 43052 42892 43064
rect 42944 43052 42950 43104
rect 43809 43095 43867 43101
rect 43809 43061 43821 43095
rect 43855 43092 43867 43095
rect 44174 43092 44180 43104
rect 43855 43064 44180 43092
rect 43855 43061 43867 43064
rect 43809 43055 43867 43061
rect 44174 43052 44180 43064
rect 44232 43052 44238 43104
rect 1104 43002 44896 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 44896 43002
rect 1104 42928 44896 42950
rect 13078 42848 13084 42900
rect 13136 42888 13142 42900
rect 22554 42888 22560 42900
rect 13136 42860 22560 42888
rect 13136 42848 13142 42860
rect 22554 42848 22560 42860
rect 22612 42848 22618 42900
rect 24486 42780 24492 42832
rect 24544 42780 24550 42832
rect 40034 42780 40040 42832
rect 40092 42780 40098 42832
rect 2777 42755 2835 42761
rect 2777 42721 2789 42755
rect 2823 42752 2835 42755
rect 2866 42752 2872 42764
rect 2823 42724 2872 42752
rect 2823 42721 2835 42724
rect 2777 42715 2835 42721
rect 2866 42712 2872 42724
rect 2924 42712 2930 42764
rect 4341 42755 4399 42761
rect 4341 42721 4353 42755
rect 4387 42752 4399 42755
rect 6641 42755 6699 42761
rect 6641 42752 6653 42755
rect 4387 42724 6653 42752
rect 4387 42721 4399 42724
rect 4341 42715 4399 42721
rect 6641 42721 6653 42724
rect 6687 42721 6699 42755
rect 10318 42752 10324 42764
rect 10279 42724 10324 42752
rect 6641 42715 6699 42721
rect 10318 42712 10324 42724
rect 10376 42712 10382 42764
rect 11606 42752 11612 42764
rect 11567 42724 11612 42752
rect 11606 42712 11612 42724
rect 11664 42712 11670 42764
rect 12250 42712 12256 42764
rect 12308 42752 12314 42764
rect 12437 42755 12495 42761
rect 12437 42752 12449 42755
rect 12308 42724 12449 42752
rect 12308 42712 12314 42724
rect 12437 42721 12449 42724
rect 12483 42721 12495 42755
rect 14826 42752 14832 42764
rect 14787 42724 14832 42752
rect 12437 42715 12495 42721
rect 14826 42712 14832 42724
rect 14884 42712 14890 42764
rect 20806 42752 20812 42764
rect 20767 42724 20812 42752
rect 20806 42712 20812 42724
rect 20864 42712 20870 42764
rect 21266 42752 21272 42764
rect 21227 42724 21272 42752
rect 21266 42712 21272 42724
rect 21324 42712 21330 42764
rect 24504 42752 24532 42780
rect 24857 42755 24915 42761
rect 24857 42752 24869 42755
rect 24504 42724 24869 42752
rect 24857 42721 24869 42724
rect 24903 42721 24915 42755
rect 24857 42715 24915 42721
rect 27062 42712 27068 42764
rect 27120 42752 27126 42764
rect 27157 42755 27215 42761
rect 27157 42752 27169 42755
rect 27120 42724 27169 42752
rect 27120 42712 27126 42724
rect 27157 42721 27169 42724
rect 27203 42721 27215 42755
rect 30466 42752 30472 42764
rect 30427 42724 30472 42752
rect 27157 42715 27215 42721
rect 30466 42712 30472 42724
rect 30524 42712 30530 42764
rect 30926 42752 30932 42764
rect 30887 42724 30932 42752
rect 30926 42712 30932 42724
rect 30984 42712 30990 42764
rect 33134 42752 33140 42764
rect 33095 42724 33140 42752
rect 33134 42712 33140 42724
rect 33192 42712 33198 42764
rect 37366 42752 37372 42764
rect 37327 42724 37372 42752
rect 37366 42712 37372 42724
rect 37424 42712 37430 42764
rect 39945 42755 40003 42761
rect 39945 42721 39957 42755
rect 39991 42752 40003 42755
rect 40052 42752 40080 42780
rect 41782 42752 41788 42764
rect 39991 42724 40080 42752
rect 41743 42724 41788 42752
rect 39991 42721 40003 42724
rect 39945 42715 40003 42721
rect 41782 42712 41788 42724
rect 41840 42712 41846 42764
rect 42337 42755 42395 42761
rect 42337 42721 42349 42755
rect 42383 42752 42395 42755
rect 42886 42752 42892 42764
rect 42383 42724 42892 42752
rect 42383 42721 42395 42724
rect 42337 42715 42395 42721
rect 42886 42712 42892 42724
rect 42944 42712 42950 42764
rect 43806 42752 43812 42764
rect 43767 42724 43812 42752
rect 43806 42712 43812 42724
rect 43864 42712 43870 42764
rect 3234 42644 3240 42696
rect 3292 42684 3298 42696
rect 3292 42656 3337 42684
rect 3292 42644 3298 42656
rect 4614 42644 4620 42696
rect 4672 42684 4678 42696
rect 4801 42687 4859 42693
rect 4801 42684 4813 42687
rect 4672 42656 4813 42684
rect 4672 42644 4678 42656
rect 4801 42653 4813 42656
rect 4847 42653 4859 42687
rect 7098 42684 7104 42696
rect 7059 42656 7104 42684
rect 4801 42647 4859 42653
rect 7098 42644 7104 42656
rect 7156 42644 7162 42696
rect 9306 42684 9312 42696
rect 9267 42656 9312 42684
rect 9306 42644 9312 42656
rect 9364 42644 9370 42696
rect 14366 42684 14372 42696
rect 14327 42656 14372 42684
rect 14366 42644 14372 42656
rect 14424 42644 14430 42696
rect 15746 42644 15752 42696
rect 15804 42684 15810 42696
rect 16669 42687 16727 42693
rect 16669 42684 16681 42687
rect 15804 42656 16681 42684
rect 15804 42644 15810 42656
rect 16669 42653 16681 42656
rect 16715 42653 16727 42687
rect 16669 42647 16727 42653
rect 23845 42687 23903 42693
rect 23845 42653 23857 42687
rect 23891 42684 23903 42687
rect 24397 42687 24455 42693
rect 24397 42684 24409 42687
rect 23891 42656 24409 42684
rect 23891 42653 23903 42656
rect 23845 42647 23903 42653
rect 24397 42653 24409 42656
rect 24443 42653 24455 42687
rect 24397 42647 24455 42653
rect 26418 42644 26424 42696
rect 26476 42684 26482 42696
rect 26697 42687 26755 42693
rect 26697 42684 26709 42687
rect 26476 42656 26709 42684
rect 26476 42644 26482 42656
rect 26697 42653 26709 42656
rect 26743 42653 26755 42687
rect 33962 42684 33968 42696
rect 33923 42656 33968 42684
rect 26697 42647 26755 42653
rect 33962 42644 33968 42656
rect 34020 42644 34026 42696
rect 35434 42684 35440 42696
rect 35395 42656 35440 42684
rect 35434 42644 35440 42656
rect 35492 42644 35498 42696
rect 36265 42687 36323 42693
rect 36265 42653 36277 42687
rect 36311 42684 36323 42687
rect 36725 42687 36783 42693
rect 36725 42684 36737 42687
rect 36311 42656 36737 42684
rect 36311 42653 36323 42656
rect 36265 42647 36323 42653
rect 36725 42653 36737 42656
rect 36771 42653 36783 42687
rect 36725 42647 36783 42653
rect 3053 42619 3111 42625
rect 3053 42585 3065 42619
rect 3099 42585 3111 42619
rect 6454 42616 6460 42628
rect 6415 42588 6460 42616
rect 3053 42579 3111 42585
rect 3068 42548 3096 42579
rect 6454 42576 6460 42588
rect 6512 42576 6518 42628
rect 9493 42619 9551 42625
rect 9493 42585 9505 42619
rect 9539 42616 9551 42619
rect 10042 42616 10048 42628
rect 9539 42588 10048 42616
rect 9539 42585 9551 42588
rect 9493 42579 9551 42585
rect 10042 42576 10048 42588
rect 10100 42576 10106 42628
rect 11790 42616 11796 42628
rect 11751 42588 11796 42616
rect 11790 42576 11796 42588
rect 11848 42576 11854 42628
rect 14550 42616 14556 42628
rect 14511 42588 14556 42616
rect 14550 42576 14556 42588
rect 14608 42576 14614 42628
rect 20990 42616 20996 42628
rect 20951 42588 20996 42616
rect 20990 42576 20996 42588
rect 21048 42576 21054 42628
rect 24578 42616 24584 42628
rect 24539 42588 24584 42616
rect 24578 42576 24584 42588
rect 24636 42576 24642 42628
rect 26881 42619 26939 42625
rect 26881 42585 26893 42619
rect 26927 42616 26939 42619
rect 27062 42616 27068 42628
rect 26927 42588 27068 42616
rect 26927 42585 26939 42588
rect 26881 42579 26939 42585
rect 27062 42576 27068 42588
rect 27120 42576 27126 42628
rect 30650 42616 30656 42628
rect 30611 42588 30656 42616
rect 30650 42576 30656 42588
rect 30708 42576 30714 42628
rect 36909 42619 36967 42625
rect 36909 42585 36921 42619
rect 36955 42616 36967 42619
rect 37826 42616 37832 42628
rect 36955 42588 37832 42616
rect 36955 42585 36967 42588
rect 36909 42579 36967 42585
rect 37826 42576 37832 42588
rect 37884 42576 37890 42628
rect 39942 42576 39948 42628
rect 40000 42616 40006 42628
rect 40129 42619 40187 42625
rect 40129 42616 40141 42619
rect 40000 42588 40141 42616
rect 40000 42576 40006 42588
rect 40129 42585 40141 42588
rect 40175 42585 40187 42619
rect 40129 42579 40187 42585
rect 42521 42619 42579 42625
rect 42521 42585 42533 42619
rect 42567 42616 42579 42619
rect 42702 42616 42708 42628
rect 42567 42588 42708 42616
rect 42567 42585 42579 42588
rect 42521 42579 42579 42585
rect 42702 42576 42708 42588
rect 42760 42576 42766 42628
rect 3142 42548 3148 42560
rect 3068 42520 3148 42548
rect 3142 42508 3148 42520
rect 3200 42508 3206 42560
rect 12526 42508 12532 42560
rect 12584 42548 12590 42560
rect 33410 42548 33416 42560
rect 12584 42520 33416 42548
rect 12584 42508 12590 42520
rect 33410 42508 33416 42520
rect 33468 42508 33474 42560
rect 1104 42458 44896 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 44896 42458
rect 1104 42384 44896 42406
rect 2590 42304 2596 42356
rect 2648 42344 2654 42356
rect 10873 42347 10931 42353
rect 2648 42316 6914 42344
rect 2648 42304 2654 42316
rect 2041 42279 2099 42285
rect 2041 42245 2053 42279
rect 2087 42276 2099 42279
rect 2774 42276 2780 42288
rect 2087 42248 2780 42276
rect 2087 42245 2099 42248
rect 2041 42239 2099 42245
rect 2774 42236 2780 42248
rect 2832 42236 2838 42288
rect 5445 42279 5503 42285
rect 5445 42245 5457 42279
rect 5491 42276 5503 42279
rect 6549 42279 6607 42285
rect 6549 42276 6561 42279
rect 5491 42248 6561 42276
rect 5491 42245 5503 42248
rect 5445 42239 5503 42245
rect 6549 42245 6561 42248
rect 6595 42245 6607 42279
rect 6886 42276 6914 42316
rect 10873 42313 10885 42347
rect 10919 42344 10931 42347
rect 11790 42344 11796 42356
rect 10919 42316 11796 42344
rect 10919 42313 10931 42316
rect 10873 42307 10931 42313
rect 11790 42304 11796 42316
rect 11848 42304 11854 42356
rect 20901 42347 20959 42353
rect 20901 42313 20913 42347
rect 20947 42344 20959 42347
rect 20990 42344 20996 42356
rect 20947 42316 20996 42344
rect 20947 42313 20959 42316
rect 20901 42307 20959 42313
rect 20990 42304 20996 42316
rect 21048 42304 21054 42356
rect 27062 42344 27068 42356
rect 27023 42316 27068 42344
rect 27062 42304 27068 42316
rect 27120 42304 27126 42356
rect 30650 42344 30656 42356
rect 30611 42316 30656 42344
rect 30650 42304 30656 42316
rect 30708 42304 30714 42356
rect 33318 42344 33324 42356
rect 33279 42316 33324 42344
rect 33318 42304 33324 42316
rect 33376 42304 33382 42356
rect 34146 42304 34152 42356
rect 34204 42344 34210 42356
rect 34882 42344 34888 42356
rect 34204 42316 34888 42344
rect 34204 42304 34210 42316
rect 34882 42304 34888 42316
rect 34940 42304 34946 42356
rect 38654 42344 38660 42356
rect 35866 42316 38660 42344
rect 12161 42279 12219 42285
rect 6886 42248 7788 42276
rect 6549 42239 6607 42245
rect 4709 42211 4767 42217
rect 4709 42177 4721 42211
rect 4755 42208 4767 42211
rect 4982 42208 4988 42220
rect 4755 42180 4988 42208
rect 4755 42177 4767 42180
rect 4709 42171 4767 42177
rect 4982 42168 4988 42180
rect 5040 42168 5046 42220
rect 5537 42211 5595 42217
rect 5537 42177 5549 42211
rect 5583 42177 5595 42211
rect 5537 42171 5595 42177
rect 1854 42140 1860 42152
rect 1815 42112 1860 42140
rect 1854 42100 1860 42112
rect 1912 42100 1918 42152
rect 2866 42140 2872 42152
rect 2827 42112 2872 42140
rect 2866 42100 2872 42112
rect 2924 42100 2930 42152
rect 5552 42072 5580 42171
rect 6365 42143 6423 42149
rect 6365 42109 6377 42143
rect 6411 42140 6423 42143
rect 7098 42140 7104 42152
rect 6411 42112 7104 42140
rect 6411 42109 6423 42112
rect 6365 42103 6423 42109
rect 7098 42100 7104 42112
rect 7156 42100 7162 42152
rect 7760 42149 7788 42248
rect 12161 42245 12173 42279
rect 12207 42276 12219 42279
rect 12434 42276 12440 42288
rect 12207 42248 12440 42276
rect 12207 42245 12219 42248
rect 12161 42239 12219 42245
rect 12434 42236 12440 42248
rect 12492 42236 12498 42288
rect 15746 42276 15752 42288
rect 14292 42248 15752 42276
rect 9306 42168 9312 42220
rect 9364 42208 9370 42220
rect 9861 42211 9919 42217
rect 9861 42208 9873 42211
rect 9364 42180 9873 42208
rect 9364 42168 9370 42180
rect 9861 42177 9873 42180
rect 9907 42177 9919 42211
rect 9861 42171 9919 42177
rect 10781 42211 10839 42217
rect 10781 42177 10793 42211
rect 10827 42177 10839 42211
rect 10781 42171 10839 42177
rect 7745 42143 7803 42149
rect 7745 42109 7757 42143
rect 7791 42109 7803 42143
rect 7745 42103 7803 42109
rect 7466 42072 7472 42084
rect 5552 42044 7472 42072
rect 7466 42032 7472 42044
rect 7524 42032 7530 42084
rect 10796 42072 10824 42171
rect 11514 42168 11520 42220
rect 11572 42208 11578 42220
rect 14292 42217 14320 42248
rect 15746 42236 15752 42248
rect 15804 42236 15810 42288
rect 16117 42279 16175 42285
rect 16117 42245 16129 42279
rect 16163 42276 16175 42279
rect 35866 42276 35894 42316
rect 38654 42304 38660 42316
rect 38712 42304 38718 42356
rect 42702 42344 42708 42356
rect 42663 42316 42708 42344
rect 42702 42304 42708 42316
rect 42760 42304 42766 42356
rect 16163 42248 35894 42276
rect 37461 42279 37519 42285
rect 16163 42245 16175 42248
rect 16117 42239 16175 42245
rect 37461 42245 37473 42279
rect 37507 42276 37519 42279
rect 38289 42279 38347 42285
rect 38289 42276 38301 42279
rect 37507 42248 38301 42276
rect 37507 42245 37519 42248
rect 37461 42239 37519 42245
rect 38289 42245 38301 42248
rect 38335 42245 38347 42279
rect 38289 42239 38347 42245
rect 39945 42279 40003 42285
rect 39945 42245 39957 42279
rect 39991 42276 40003 42279
rect 42610 42276 42616 42288
rect 39991 42248 42616 42276
rect 39991 42245 40003 42248
rect 39945 42239 40003 42245
rect 42610 42236 42616 42248
rect 42668 42236 42674 42288
rect 11977 42211 12035 42217
rect 11977 42208 11989 42211
rect 11572 42180 11989 42208
rect 11572 42168 11578 42180
rect 11977 42177 11989 42180
rect 12023 42177 12035 42211
rect 11977 42171 12035 42177
rect 14277 42211 14335 42217
rect 14277 42177 14289 42211
rect 14323 42177 14335 42211
rect 20806 42208 20812 42220
rect 20767 42180 20812 42208
rect 14277 42171 14335 42177
rect 20806 42168 20812 42180
rect 20864 42168 20870 42220
rect 22646 42208 22652 42220
rect 22607 42180 22652 42208
rect 22646 42168 22652 42180
rect 22704 42168 22710 42220
rect 26418 42208 26424 42220
rect 26379 42180 26424 42208
rect 26418 42168 26424 42180
rect 26476 42168 26482 42220
rect 27157 42211 27215 42217
rect 27157 42177 27169 42211
rect 27203 42177 27215 42211
rect 27798 42208 27804 42220
rect 27759 42180 27804 42208
rect 27157 42171 27215 42177
rect 12894 42140 12900 42152
rect 12855 42112 12900 42140
rect 12894 42100 12900 42112
rect 12952 42100 12958 42152
rect 14458 42140 14464 42152
rect 14419 42112 14464 42140
rect 14458 42100 14464 42112
rect 14516 42100 14522 42152
rect 22830 42140 22836 42152
rect 22791 42112 22836 42140
rect 22830 42100 22836 42112
rect 22888 42100 22894 42152
rect 23198 42140 23204 42152
rect 23159 42112 23204 42140
rect 23198 42100 23204 42112
rect 23256 42100 23262 42152
rect 27172 42140 27200 42171
rect 27798 42168 27804 42180
rect 27856 42168 27862 42220
rect 30558 42208 30564 42220
rect 30519 42180 30564 42208
rect 30558 42168 30564 42180
rect 30616 42168 30622 42220
rect 33410 42208 33416 42220
rect 33371 42180 33416 42208
rect 33410 42168 33416 42180
rect 33468 42168 33474 42220
rect 33962 42208 33968 42220
rect 33923 42180 33968 42208
rect 33962 42168 33968 42180
rect 34020 42168 34026 42220
rect 36446 42208 36452 42220
rect 36407 42180 36452 42208
rect 36446 42168 36452 42180
rect 36504 42208 36510 42220
rect 37369 42211 37427 42217
rect 37369 42208 37381 42211
rect 36504 42180 37381 42208
rect 36504 42168 36510 42180
rect 37369 42177 37381 42180
rect 37415 42177 37427 42211
rect 42794 42208 42800 42220
rect 42755 42180 42800 42208
rect 37369 42171 37427 42177
rect 42794 42168 42800 42180
rect 42852 42168 42858 42220
rect 43441 42211 43499 42217
rect 43441 42208 43453 42211
rect 42904 42180 43453 42208
rect 27985 42143 28043 42149
rect 27172 42112 27844 42140
rect 13998 42072 14004 42084
rect 10796 42044 14004 42072
rect 13998 42032 14004 42044
rect 14056 42032 14062 42084
rect 20806 42032 20812 42084
rect 20864 42072 20870 42084
rect 27062 42072 27068 42084
rect 20864 42044 27068 42072
rect 20864 42032 20870 42044
rect 27062 42032 27068 42044
rect 27120 42032 27126 42084
rect 4801 42007 4859 42013
rect 4801 41973 4813 42007
rect 4847 42004 4859 42007
rect 6362 42004 6368 42016
rect 4847 41976 6368 42004
rect 4847 41973 4859 41976
rect 4801 41967 4859 41973
rect 6362 41964 6368 41976
rect 6420 41964 6426 42016
rect 27816 42004 27844 42112
rect 27985 42109 27997 42143
rect 28031 42140 28043 42143
rect 28074 42140 28080 42152
rect 28031 42112 28080 42140
rect 28031 42109 28043 42112
rect 27985 42103 28043 42109
rect 28074 42100 28080 42112
rect 28132 42100 28138 42152
rect 28350 42140 28356 42152
rect 28311 42112 28356 42140
rect 28350 42100 28356 42112
rect 28408 42100 28414 42152
rect 34149 42143 34207 42149
rect 34149 42109 34161 42143
rect 34195 42140 34207 42143
rect 34790 42140 34796 42152
rect 34195 42112 34796 42140
rect 34195 42109 34207 42112
rect 34149 42103 34207 42109
rect 34790 42100 34796 42112
rect 34848 42100 34854 42152
rect 34882 42100 34888 42152
rect 34940 42140 34946 42152
rect 38105 42143 38163 42149
rect 34940 42112 34985 42140
rect 35268 42112 38056 42140
rect 34940 42100 34946 42112
rect 35268 42004 35296 42112
rect 35342 42032 35348 42084
rect 35400 42072 35406 42084
rect 38028 42072 38056 42112
rect 38105 42109 38117 42143
rect 38151 42140 38163 42143
rect 38378 42140 38384 42152
rect 38151 42112 38384 42140
rect 38151 42109 38163 42112
rect 38105 42103 38163 42109
rect 38378 42100 38384 42112
rect 38436 42100 38442 42152
rect 42794 42072 42800 42084
rect 35400 42044 37964 42072
rect 38028 42044 42800 42072
rect 35400 42032 35406 42044
rect 27816 41976 35296 42004
rect 35618 41964 35624 42016
rect 35676 42004 35682 42016
rect 36357 42007 36415 42013
rect 36357 42004 36369 42007
rect 35676 41976 36369 42004
rect 35676 41964 35682 41976
rect 36357 41973 36369 41976
rect 36403 41973 36415 42007
rect 37936 42004 37964 42044
rect 42794 42032 42800 42044
rect 42852 42032 42858 42084
rect 42904 42004 42932 42180
rect 43441 42177 43453 42180
rect 43487 42208 43499 42211
rect 43530 42208 43536 42220
rect 43487 42180 43536 42208
rect 43487 42177 43499 42180
rect 43441 42171 43499 42177
rect 43530 42168 43536 42180
rect 43588 42168 43594 42220
rect 43898 42208 43904 42220
rect 43859 42180 43904 42208
rect 43898 42168 43904 42180
rect 43956 42168 43962 42220
rect 43346 42004 43352 42016
rect 37936 41976 42932 42004
rect 43307 41976 43352 42004
rect 36357 41967 36415 41973
rect 43346 41964 43352 41976
rect 43404 41964 43410 42016
rect 43990 42004 43996 42016
rect 43951 41976 43996 42004
rect 43990 41964 43996 41976
rect 44048 41964 44054 42016
rect 1104 41914 44896 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 44896 41914
rect 1104 41840 44896 41862
rect 3881 41803 3939 41809
rect 3881 41769 3893 41803
rect 3927 41800 3939 41803
rect 3970 41800 3976 41812
rect 3927 41772 3976 41800
rect 3927 41769 3939 41772
rect 3881 41763 3939 41769
rect 3970 41760 3976 41772
rect 4028 41760 4034 41812
rect 4982 41760 4988 41812
rect 5040 41800 5046 41812
rect 10042 41800 10048 41812
rect 5040 41772 6914 41800
rect 10003 41772 10048 41800
rect 5040 41760 5046 41772
rect 2958 41732 2964 41744
rect 2792 41704 2964 41732
rect 2792 41673 2820 41704
rect 2958 41692 2964 41704
rect 3016 41692 3022 41744
rect 6886 41732 6914 41772
rect 10042 41760 10048 41772
rect 10100 41760 10106 41812
rect 14550 41800 14556 41812
rect 14511 41772 14556 41800
rect 14550 41760 14556 41772
rect 14608 41760 14614 41812
rect 22741 41803 22799 41809
rect 22741 41769 22753 41803
rect 22787 41800 22799 41803
rect 22830 41800 22836 41812
rect 22787 41772 22836 41800
rect 22787 41769 22799 41772
rect 22741 41763 22799 41769
rect 22830 41760 22836 41772
rect 22888 41760 22894 41812
rect 23385 41803 23443 41809
rect 23385 41769 23397 41803
rect 23431 41800 23443 41803
rect 23474 41800 23480 41812
rect 23431 41772 23480 41800
rect 23431 41769 23443 41772
rect 23385 41763 23443 41769
rect 23474 41760 23480 41772
rect 23532 41760 23538 41812
rect 24489 41803 24547 41809
rect 24489 41769 24501 41803
rect 24535 41800 24547 41803
rect 24578 41800 24584 41812
rect 24535 41772 24584 41800
rect 24535 41769 24547 41772
rect 24489 41763 24547 41769
rect 24578 41760 24584 41772
rect 24636 41760 24642 41812
rect 28074 41800 28080 41812
rect 28035 41772 28080 41800
rect 28074 41760 28080 41772
rect 28132 41760 28138 41812
rect 34790 41800 34796 41812
rect 34751 41772 34796 41800
rect 34790 41760 34796 41772
rect 34848 41760 34854 41812
rect 37826 41800 37832 41812
rect 37787 41772 37832 41800
rect 37826 41760 37832 41772
rect 37884 41760 37890 41812
rect 38378 41800 38384 41812
rect 38339 41772 38384 41800
rect 38378 41760 38384 41772
rect 38436 41760 38442 41812
rect 39942 41800 39948 41812
rect 39903 41772 39948 41800
rect 39942 41760 39948 41772
rect 40000 41760 40006 41812
rect 12158 41732 12164 41744
rect 6886 41704 12164 41732
rect 12158 41692 12164 41704
rect 12216 41692 12222 41744
rect 14366 41692 14372 41744
rect 14424 41732 14430 41744
rect 15105 41735 15163 41741
rect 15105 41732 15117 41735
rect 14424 41704 15117 41732
rect 14424 41692 14430 41704
rect 15105 41701 15117 41704
rect 15151 41701 15163 41735
rect 15105 41695 15163 41701
rect 30558 41692 30564 41744
rect 30616 41732 30622 41744
rect 42886 41732 42892 41744
rect 30616 41704 42892 41732
rect 30616 41692 30622 41704
rect 42886 41692 42892 41704
rect 42944 41732 42950 41744
rect 43898 41732 43904 41744
rect 42944 41704 43904 41732
rect 42944 41692 42950 41704
rect 43898 41692 43904 41704
rect 43956 41692 43962 41744
rect 2777 41667 2835 41673
rect 2777 41633 2789 41667
rect 2823 41633 2835 41667
rect 2777 41627 2835 41633
rect 2866 41624 2872 41676
rect 2924 41664 2930 41676
rect 3237 41667 3295 41673
rect 3237 41664 3249 41667
rect 2924 41636 3249 41664
rect 2924 41624 2930 41636
rect 3237 41633 3249 41636
rect 3283 41633 3295 41667
rect 5166 41664 5172 41676
rect 5127 41636 5172 41664
rect 3237 41627 3295 41633
rect 5166 41624 5172 41636
rect 5224 41624 5230 41676
rect 6362 41664 6368 41676
rect 6323 41636 6368 41664
rect 6362 41624 6368 41636
rect 6420 41624 6426 41676
rect 6546 41664 6552 41676
rect 6507 41636 6552 41664
rect 6546 41624 6552 41636
rect 6604 41624 6610 41676
rect 27062 41624 27068 41676
rect 27120 41664 27126 41676
rect 35250 41664 35256 41676
rect 27120 41636 35256 41664
rect 27120 41624 27126 41636
rect 35250 41624 35256 41636
rect 35308 41624 35314 41676
rect 35434 41664 35440 41676
rect 35395 41636 35440 41664
rect 35434 41624 35440 41636
rect 35492 41624 35498 41676
rect 35618 41664 35624 41676
rect 35579 41636 35624 41664
rect 35618 41624 35624 41636
rect 35676 41624 35682 41676
rect 36078 41664 36084 41676
rect 36039 41636 36084 41664
rect 36078 41624 36084 41636
rect 36136 41624 36142 41676
rect 42518 41664 42524 41676
rect 42479 41636 42524 41664
rect 42518 41624 42524 41636
rect 42576 41624 42582 41676
rect 43990 41664 43996 41676
rect 43951 41636 43996 41664
rect 43990 41624 43996 41636
rect 44048 41624 44054 41676
rect 44174 41664 44180 41676
rect 44135 41636 44180 41664
rect 44174 41624 44180 41636
rect 44232 41624 44238 41676
rect 3973 41599 4031 41605
rect 3973 41565 3985 41599
rect 4019 41596 4031 41599
rect 4614 41596 4620 41608
rect 4019 41568 4620 41596
rect 4019 41565 4031 41568
rect 3973 41559 4031 41565
rect 4614 41556 4620 41568
rect 4672 41556 4678 41608
rect 10137 41599 10195 41605
rect 10137 41565 10149 41599
rect 10183 41565 10195 41599
rect 10137 41559 10195 41565
rect 11517 41599 11575 41605
rect 11517 41565 11529 41599
rect 11563 41596 11575 41599
rect 12066 41596 12072 41608
rect 11563 41568 12072 41596
rect 11563 41565 11575 41568
rect 11517 41559 11575 41565
rect 3050 41528 3056 41540
rect 3011 41500 3056 41528
rect 3050 41488 3056 41500
rect 3108 41488 3114 41540
rect 10152 41528 10180 41559
rect 12066 41556 12072 41568
rect 12124 41556 12130 41608
rect 14461 41599 14519 41605
rect 14461 41565 14473 41599
rect 14507 41596 14519 41599
rect 14642 41596 14648 41608
rect 14507 41568 14648 41596
rect 14507 41565 14519 41568
rect 14461 41559 14519 41565
rect 14642 41556 14648 41568
rect 14700 41556 14706 41608
rect 22554 41556 22560 41608
rect 22612 41596 22618 41608
rect 22649 41599 22707 41605
rect 22649 41596 22661 41599
rect 22612 41568 22661 41596
rect 22612 41556 22618 41568
rect 22649 41565 22661 41568
rect 22695 41565 22707 41599
rect 22649 41559 22707 41565
rect 22830 41556 22836 41608
rect 22888 41596 22894 41608
rect 23293 41599 23351 41605
rect 23293 41596 23305 41599
rect 22888 41568 23305 41596
rect 22888 41556 22894 41568
rect 23293 41565 23305 41568
rect 23339 41565 23351 41599
rect 24394 41596 24400 41608
rect 24355 41568 24400 41596
rect 23293 41559 23351 41565
rect 24394 41556 24400 41568
rect 24452 41556 24458 41608
rect 28166 41596 28172 41608
rect 26206 41568 28172 41596
rect 10962 41528 10968 41540
rect 10152 41500 10968 41528
rect 10962 41488 10968 41500
rect 11020 41488 11026 41540
rect 12897 41531 12955 41537
rect 12897 41497 12909 41531
rect 12943 41528 12955 41531
rect 12986 41528 12992 41540
rect 12943 41500 12992 41528
rect 12943 41497 12955 41500
rect 12897 41491 12955 41497
rect 12986 41488 12992 41500
rect 13044 41528 13050 41540
rect 26206 41528 26234 41568
rect 28166 41556 28172 41568
rect 28224 41556 28230 41608
rect 34514 41556 34520 41608
rect 34572 41596 34578 41608
rect 34885 41599 34943 41605
rect 34885 41596 34897 41599
rect 34572 41568 34897 41596
rect 34572 41556 34578 41568
rect 34885 41565 34897 41568
rect 34931 41565 34943 41599
rect 37918 41596 37924 41608
rect 37879 41568 37924 41596
rect 34885 41559 34943 41565
rect 37918 41556 37924 41568
rect 37976 41556 37982 41608
rect 39850 41596 39856 41608
rect 39811 41568 39856 41596
rect 39850 41556 39856 41568
rect 39908 41556 39914 41608
rect 13044 41500 26234 41528
rect 13044 41488 13050 41500
rect 43254 41420 43260 41472
rect 43312 41460 43318 41472
rect 44450 41460 44456 41472
rect 43312 41432 44456 41460
rect 43312 41420 43318 41432
rect 44450 41420 44456 41432
rect 44508 41420 44514 41472
rect 1104 41370 44896 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 44896 41370
rect 1104 41296 44896 41318
rect 2961 41259 3019 41265
rect 2961 41225 2973 41259
rect 3007 41256 3019 41259
rect 3050 41256 3056 41268
rect 3007 41228 3056 41256
rect 3007 41225 3019 41228
rect 2961 41219 3019 41225
rect 3050 41216 3056 41228
rect 3108 41216 3114 41268
rect 6454 41256 6460 41268
rect 6415 41228 6460 41256
rect 6454 41216 6460 41228
rect 6512 41216 6518 41268
rect 12526 41256 12532 41268
rect 6886 41228 12532 41256
rect 2317 41191 2375 41197
rect 2317 41157 2329 41191
rect 2363 41188 2375 41191
rect 3142 41188 3148 41200
rect 2363 41160 3148 41188
rect 2363 41157 2375 41160
rect 2317 41151 2375 41157
rect 3142 41148 3148 41160
rect 3200 41148 3206 41200
rect 6886 41188 6914 41228
rect 12526 41216 12532 41228
rect 12584 41216 12590 41268
rect 14185 41259 14243 41265
rect 14185 41225 14197 41259
rect 14231 41256 14243 41259
rect 14458 41256 14464 41268
rect 14231 41228 14464 41256
rect 14231 41225 14243 41228
rect 14185 41219 14243 41225
rect 14458 41216 14464 41228
rect 14516 41216 14522 41268
rect 39850 41256 39856 41268
rect 15304 41228 39856 41256
rect 9306 41188 9312 41200
rect 4724 41160 6914 41188
rect 9048 41160 9312 41188
rect 1765 41123 1823 41129
rect 1765 41089 1777 41123
rect 1811 41120 1823 41123
rect 1854 41120 1860 41132
rect 1811 41092 1860 41120
rect 1811 41089 1823 41092
rect 1765 41083 1823 41089
rect 1854 41080 1860 41092
rect 1912 41080 1918 41132
rect 2409 41123 2467 41129
rect 2409 41120 2421 41123
rect 2332 41092 2421 41120
rect 2332 41064 2360 41092
rect 2409 41089 2421 41092
rect 2455 41089 2467 41123
rect 2409 41083 2467 41089
rect 3053 41123 3111 41129
rect 3053 41089 3065 41123
rect 3099 41089 3111 41123
rect 3053 41083 3111 41089
rect 2314 41012 2320 41064
rect 2372 41012 2378 41064
rect 3068 40984 3096 41083
rect 3234 41080 3240 41132
rect 3292 41120 3298 41132
rect 3513 41123 3571 41129
rect 3513 41120 3525 41123
rect 3292 41092 3525 41120
rect 3292 41080 3298 41092
rect 3513 41089 3525 41092
rect 3559 41089 3571 41123
rect 3513 41083 3571 41089
rect 4724 41064 4752 41160
rect 5445 41123 5503 41129
rect 5445 41089 5457 41123
rect 5491 41120 5503 41123
rect 5626 41120 5632 41132
rect 5491 41092 5632 41120
rect 5491 41089 5503 41092
rect 5445 41083 5503 41089
rect 5626 41080 5632 41092
rect 5684 41080 5690 41132
rect 9048 41129 9076 41160
rect 9306 41148 9312 41160
rect 9364 41188 9370 41200
rect 15304 41188 15332 41228
rect 39850 41216 39856 41228
rect 39908 41216 39914 41268
rect 41386 41228 43576 41256
rect 41386 41188 41414 41228
rect 9364 41160 15332 41188
rect 22066 41160 41414 41188
rect 41693 41191 41751 41197
rect 9364 41148 9370 41160
rect 6549 41123 6607 41129
rect 6549 41089 6561 41123
rect 6595 41120 6607 41123
rect 9033 41123 9091 41129
rect 6595 41092 6684 41120
rect 6595 41089 6607 41092
rect 6549 41083 6607 41089
rect 6656 41064 6684 41092
rect 9033 41089 9045 41123
rect 9079 41089 9091 41123
rect 10686 41120 10692 41132
rect 10647 41092 10692 41120
rect 9033 41083 9091 41089
rect 10686 41080 10692 41092
rect 10744 41080 10750 41132
rect 11054 41080 11060 41132
rect 11112 41120 11118 41132
rect 11885 41123 11943 41129
rect 11885 41120 11897 41123
rect 11112 41092 11897 41120
rect 11112 41080 11118 41092
rect 11885 41089 11897 41092
rect 11931 41120 11943 41123
rect 12066 41120 12072 41132
rect 11931 41092 12072 41120
rect 11931 41089 11943 41092
rect 11885 41083 11943 41089
rect 12066 41080 12072 41092
rect 12124 41080 12130 41132
rect 13998 41080 14004 41132
rect 14056 41120 14062 41132
rect 14093 41123 14151 41129
rect 14093 41120 14105 41123
rect 14056 41092 14105 41120
rect 14056 41080 14062 41092
rect 14093 41089 14105 41092
rect 14139 41089 14151 41123
rect 14093 41083 14151 41089
rect 14642 41080 14648 41132
rect 14700 41120 14706 41132
rect 22066 41120 22094 41160
rect 41693 41157 41705 41191
rect 41739 41188 41751 41191
rect 43441 41191 43499 41197
rect 43441 41188 43453 41191
rect 41739 41160 43453 41188
rect 41739 41157 41751 41160
rect 41693 41151 41751 41157
rect 43441 41157 43453 41160
rect 43487 41157 43499 41191
rect 43441 41151 43499 41157
rect 32490 41120 32496 41132
rect 14700 41092 22094 41120
rect 32451 41092 32496 41120
rect 14700 41080 14706 41092
rect 32490 41080 32496 41092
rect 32548 41080 32554 41132
rect 32582 41080 32588 41132
rect 32640 41120 32646 41132
rect 32769 41123 32827 41129
rect 32640 41092 32685 41120
rect 32640 41080 32646 41092
rect 32769 41089 32781 41123
rect 32815 41120 32827 41123
rect 33042 41120 33048 41132
rect 32815 41092 33048 41120
rect 32815 41089 32827 41092
rect 32769 41083 32827 41089
rect 33042 41080 33048 41092
rect 33100 41080 33106 41132
rect 33410 41120 33416 41132
rect 33371 41092 33416 41120
rect 33410 41080 33416 41092
rect 33468 41080 33474 41132
rect 43349 41123 43407 41129
rect 43349 41089 43361 41123
rect 43395 41120 43407 41123
rect 43548 41120 43576 41228
rect 43395 41092 43576 41120
rect 43395 41089 43407 41092
rect 43349 41083 43407 41089
rect 43456 41064 43484 41092
rect 4706 41052 4712 41064
rect 4667 41024 4712 41052
rect 4706 41012 4712 41024
rect 4764 41012 4770 41064
rect 6638 41012 6644 41064
rect 6696 41052 6702 41064
rect 9582 41052 9588 41064
rect 6696 41024 6914 41052
rect 9543 41024 9588 41052
rect 6696 41012 6702 41024
rect 4798 40984 4804 40996
rect 3068 40956 4804 40984
rect 4798 40944 4804 40956
rect 4856 40944 4862 40996
rect 6886 40984 6914 41024
rect 9582 41012 9588 41024
rect 9640 41012 9646 41064
rect 36446 41052 36452 41064
rect 10704 41024 36452 41052
rect 10704 40984 10732 41024
rect 36446 41012 36452 41024
rect 36504 41012 36510 41064
rect 41325 41055 41383 41061
rect 41325 41021 41337 41055
rect 41371 41052 41383 41055
rect 41506 41052 41512 41064
rect 41371 41024 41512 41052
rect 41371 41021 41383 41024
rect 41325 41015 41383 41021
rect 41506 41012 41512 41024
rect 41564 41012 41570 41064
rect 41877 41055 41935 41061
rect 41877 41021 41889 41055
rect 41923 41052 41935 41055
rect 42705 41055 42763 41061
rect 42705 41052 42717 41055
rect 41923 41024 42717 41052
rect 41923 41021 41935 41024
rect 41877 41015 41935 41021
rect 42705 41021 42717 41024
rect 42751 41021 42763 41055
rect 42705 41015 42763 41021
rect 43438 41012 43444 41064
rect 43496 41012 43502 41064
rect 6886 40956 10732 40984
rect 10873 40987 10931 40993
rect 10873 40953 10885 40987
rect 10919 40984 10931 40987
rect 11054 40984 11060 40996
rect 10919 40956 11060 40984
rect 10919 40953 10931 40956
rect 10873 40947 10931 40953
rect 11054 40944 11060 40956
rect 11112 40944 11118 40996
rect 30558 40984 30564 40996
rect 11900 40956 30564 40984
rect 9582 40876 9588 40928
rect 9640 40916 9646 40928
rect 11900 40916 11928 40956
rect 30558 40944 30564 40956
rect 30616 40944 30622 40996
rect 9640 40888 11928 40916
rect 9640 40876 9646 40888
rect 13262 40876 13268 40928
rect 13320 40916 13326 40928
rect 13357 40919 13415 40925
rect 13357 40916 13369 40919
rect 13320 40888 13369 40916
rect 13320 40876 13326 40888
rect 13357 40885 13369 40888
rect 13403 40916 13415 40919
rect 22830 40916 22836 40928
rect 13403 40888 22836 40916
rect 13403 40885 13415 40888
rect 13357 40879 13415 40885
rect 22830 40876 22836 40888
rect 22888 40916 22894 40928
rect 23382 40916 23388 40928
rect 22888 40888 23388 40916
rect 22888 40876 22894 40888
rect 23382 40876 23388 40888
rect 23440 40876 23446 40928
rect 32953 40919 33011 40925
rect 32953 40885 32965 40919
rect 32999 40916 33011 40919
rect 33318 40916 33324 40928
rect 32999 40888 33324 40916
rect 32999 40885 33011 40888
rect 32953 40879 33011 40885
rect 33318 40876 33324 40888
rect 33376 40876 33382 40928
rect 33594 40916 33600 40928
rect 33555 40888 33600 40916
rect 33594 40876 33600 40888
rect 33652 40876 33658 40928
rect 44174 40916 44180 40928
rect 44135 40888 44180 40916
rect 44174 40876 44180 40888
rect 44232 40876 44238 40928
rect 1104 40826 44896 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 44896 40826
rect 1104 40752 44896 40774
rect 2866 40712 2872 40724
rect 2827 40684 2872 40712
rect 2866 40672 2872 40684
rect 2924 40672 2930 40724
rect 13449 40715 13507 40721
rect 13449 40681 13461 40715
rect 13495 40712 13507 40715
rect 14090 40712 14096 40724
rect 13495 40684 14096 40712
rect 13495 40681 13507 40684
rect 13449 40675 13507 40681
rect 14090 40672 14096 40684
rect 14148 40672 14154 40724
rect 32306 40712 32312 40724
rect 32219 40684 32312 40712
rect 32306 40672 32312 40684
rect 32364 40712 32370 40724
rect 32490 40712 32496 40724
rect 32364 40684 32496 40712
rect 32364 40672 32370 40684
rect 32490 40672 32496 40684
rect 32548 40672 32554 40724
rect 2314 40604 2320 40656
rect 2372 40644 2378 40656
rect 37277 40647 37335 40653
rect 2372 40616 12204 40644
rect 2372 40604 2378 40616
rect 10686 40576 10692 40588
rect 3896 40548 10692 40576
rect 3896 40520 3924 40548
rect 10686 40536 10692 40548
rect 10744 40536 10750 40588
rect 12176 40585 12204 40616
rect 37277 40613 37289 40647
rect 37323 40644 37335 40647
rect 37366 40644 37372 40656
rect 37323 40616 37372 40644
rect 37323 40613 37335 40616
rect 37277 40607 37335 40613
rect 37366 40604 37372 40616
rect 37424 40604 37430 40656
rect 40678 40604 40684 40656
rect 40736 40644 40742 40656
rect 40773 40647 40831 40653
rect 40773 40644 40785 40647
rect 40736 40616 40785 40644
rect 40736 40604 40742 40616
rect 40773 40613 40785 40616
rect 40819 40613 40831 40647
rect 40773 40607 40831 40613
rect 12161 40579 12219 40585
rect 12161 40545 12173 40579
rect 12207 40545 12219 40579
rect 12161 40539 12219 40545
rect 27433 40579 27491 40585
rect 27433 40545 27445 40579
rect 27479 40576 27491 40579
rect 28902 40576 28908 40588
rect 27479 40548 28908 40576
rect 27479 40545 27491 40548
rect 27433 40539 27491 40545
rect 28902 40536 28908 40548
rect 28960 40536 28966 40588
rect 43254 40576 43260 40588
rect 43215 40548 43260 40576
rect 43254 40536 43260 40548
rect 43312 40536 43318 40588
rect 43346 40536 43352 40588
rect 43404 40576 43410 40588
rect 43993 40579 44051 40585
rect 43993 40576 44005 40579
rect 43404 40548 44005 40576
rect 43404 40536 43410 40548
rect 43993 40545 44005 40548
rect 44039 40545 44051 40579
rect 44174 40576 44180 40588
rect 44135 40548 44180 40576
rect 43993 40539 44051 40545
rect 44174 40536 44180 40548
rect 44232 40536 44238 40588
rect 1946 40468 1952 40520
rect 2004 40508 2010 40520
rect 2041 40511 2099 40517
rect 2041 40508 2053 40511
rect 2004 40480 2053 40508
rect 2004 40468 2010 40480
rect 2041 40477 2053 40480
rect 2087 40477 2099 40511
rect 2041 40471 2099 40477
rect 3602 40468 3608 40520
rect 3660 40508 3666 40520
rect 3878 40508 3884 40520
rect 3660 40480 3884 40508
rect 3660 40468 3666 40480
rect 3878 40468 3884 40480
rect 3936 40468 3942 40520
rect 4617 40511 4675 40517
rect 4617 40508 4629 40511
rect 4080 40480 4629 40508
rect 4080 40381 4108 40480
rect 4617 40477 4629 40480
rect 4663 40508 4675 40511
rect 5626 40508 5632 40520
rect 4663 40480 5632 40508
rect 4663 40477 4675 40480
rect 4617 40471 4675 40477
rect 5626 40468 5632 40480
rect 5684 40508 5690 40520
rect 6917 40511 6975 40517
rect 6917 40508 6929 40511
rect 5684 40480 6929 40508
rect 5684 40468 5690 40480
rect 6917 40477 6929 40480
rect 6963 40477 6975 40511
rect 6917 40471 6975 40477
rect 8846 40468 8852 40520
rect 8904 40508 8910 40520
rect 9306 40508 9312 40520
rect 8904 40480 9312 40508
rect 8904 40468 8910 40480
rect 9306 40468 9312 40480
rect 9364 40468 9370 40520
rect 11977 40511 12035 40517
rect 10060 40480 11376 40508
rect 7466 40440 7472 40452
rect 7379 40412 7472 40440
rect 7466 40400 7472 40412
rect 7524 40440 7530 40452
rect 10060 40440 10088 40480
rect 7524 40412 10088 40440
rect 7524 40400 7530 40412
rect 10134 40400 10140 40452
rect 10192 40440 10198 40452
rect 11348 40440 11376 40480
rect 11977 40477 11989 40511
rect 12023 40508 12035 40511
rect 12066 40508 12072 40520
rect 12023 40480 12072 40508
rect 12023 40477 12035 40480
rect 11977 40471 12035 40477
rect 12066 40468 12072 40480
rect 12124 40468 12130 40520
rect 27617 40511 27675 40517
rect 27617 40477 27629 40511
rect 27663 40477 27675 40511
rect 31110 40508 31116 40520
rect 31071 40480 31116 40508
rect 27617 40471 27675 40477
rect 14642 40440 14648 40452
rect 10192 40412 11192 40440
rect 11348 40412 14648 40440
rect 10192 40400 10198 40412
rect 4065 40375 4123 40381
rect 4065 40341 4077 40375
rect 4111 40341 4123 40375
rect 5902 40372 5908 40384
rect 5863 40344 5908 40372
rect 4065 40335 4123 40341
rect 5902 40332 5908 40344
rect 5960 40332 5966 40384
rect 11164 40372 11192 40412
rect 14642 40400 14648 40412
rect 14700 40400 14706 40452
rect 26418 40400 26424 40452
rect 26476 40440 26482 40452
rect 27632 40440 27660 40471
rect 31110 40468 31116 40480
rect 31168 40468 31174 40520
rect 32122 40508 32128 40520
rect 32083 40480 32128 40508
rect 32122 40468 32128 40480
rect 32180 40468 32186 40520
rect 34149 40511 34207 40517
rect 34149 40508 34161 40511
rect 32232 40480 34161 40508
rect 26476 40412 27660 40440
rect 26476 40400 26482 40412
rect 30742 40400 30748 40452
rect 30800 40440 30806 40452
rect 32232 40440 32260 40480
rect 34149 40477 34161 40480
rect 34195 40477 34207 40511
rect 34149 40471 34207 40477
rect 35069 40511 35127 40517
rect 35069 40477 35081 40511
rect 35115 40508 35127 40511
rect 35342 40508 35348 40520
rect 35115 40480 35348 40508
rect 35115 40477 35127 40480
rect 35069 40471 35127 40477
rect 35342 40468 35348 40480
rect 35400 40468 35406 40520
rect 37001 40511 37059 40517
rect 37001 40477 37013 40511
rect 37047 40508 37059 40511
rect 37734 40508 37740 40520
rect 37047 40480 37740 40508
rect 37047 40477 37059 40480
rect 37001 40471 37059 40477
rect 37734 40468 37740 40480
rect 37792 40468 37798 40520
rect 39301 40511 39359 40517
rect 39301 40477 39313 40511
rect 39347 40508 39359 40511
rect 39942 40508 39948 40520
rect 39347 40480 39948 40508
rect 39347 40477 39359 40480
rect 39301 40471 39359 40477
rect 39942 40468 39948 40480
rect 40000 40468 40006 40520
rect 40034 40468 40040 40520
rect 40092 40508 40098 40520
rect 40494 40508 40500 40520
rect 40092 40480 40137 40508
rect 40455 40480 40500 40508
rect 40092 40468 40098 40480
rect 40494 40468 40500 40480
rect 40552 40468 40558 40520
rect 30800 40412 32260 40440
rect 30800 40400 30806 40412
rect 33594 40400 33600 40452
rect 33652 40440 33658 40452
rect 33882 40443 33940 40449
rect 33882 40440 33894 40443
rect 33652 40412 33894 40440
rect 33652 40400 33658 40412
rect 33882 40409 33894 40412
rect 33928 40409 33940 40443
rect 37274 40440 37280 40452
rect 37235 40412 37280 40440
rect 33882 40403 33940 40409
rect 37274 40400 37280 40412
rect 37332 40400 37338 40452
rect 39056 40443 39114 40449
rect 39056 40409 39068 40443
rect 39102 40440 39114 40443
rect 40770 40440 40776 40452
rect 39102 40412 39896 40440
rect 40731 40412 40776 40440
rect 39102 40409 39114 40412
rect 39056 40403 39114 40409
rect 20806 40372 20812 40384
rect 11164 40344 20812 40372
rect 20806 40332 20812 40344
rect 20864 40332 20870 40384
rect 27801 40375 27859 40381
rect 27801 40341 27813 40375
rect 27847 40372 27859 40375
rect 28074 40372 28080 40384
rect 27847 40344 28080 40372
rect 27847 40341 27859 40344
rect 27801 40335 27859 40341
rect 28074 40332 28080 40344
rect 28132 40332 28138 40384
rect 30929 40375 30987 40381
rect 30929 40341 30941 40375
rect 30975 40372 30987 40375
rect 31018 40372 31024 40384
rect 30975 40344 31024 40372
rect 30975 40341 30987 40344
rect 30929 40335 30987 40341
rect 31018 40332 31024 40344
rect 31076 40332 31082 40384
rect 32769 40375 32827 40381
rect 32769 40341 32781 40375
rect 32815 40372 32827 40375
rect 33042 40372 33048 40384
rect 32815 40344 33048 40372
rect 32815 40341 32827 40344
rect 32769 40335 32827 40341
rect 33042 40332 33048 40344
rect 33100 40332 33106 40384
rect 35250 40372 35256 40384
rect 35211 40344 35256 40372
rect 35250 40332 35256 40344
rect 35308 40332 35314 40384
rect 37093 40375 37151 40381
rect 37093 40341 37105 40375
rect 37139 40372 37151 40375
rect 37642 40372 37648 40384
rect 37139 40344 37648 40372
rect 37139 40341 37151 40344
rect 37093 40335 37151 40341
rect 37642 40332 37648 40344
rect 37700 40332 37706 40384
rect 37921 40375 37979 40381
rect 37921 40341 37933 40375
rect 37967 40372 37979 40375
rect 39206 40372 39212 40384
rect 37967 40344 39212 40372
rect 37967 40341 37979 40344
rect 37921 40335 37979 40341
rect 39206 40332 39212 40344
rect 39264 40332 39270 40384
rect 39868 40381 39896 40412
rect 40770 40400 40776 40412
rect 40828 40400 40834 40452
rect 39853 40375 39911 40381
rect 39853 40341 39865 40375
rect 39899 40341 39911 40375
rect 40586 40372 40592 40384
rect 40547 40344 40592 40372
rect 39853 40335 39911 40341
rect 40586 40332 40592 40344
rect 40644 40332 40650 40384
rect 1104 40282 44896 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 44896 40282
rect 1104 40208 44896 40230
rect 4614 40128 4620 40180
rect 4672 40168 4678 40180
rect 13078 40168 13084 40180
rect 4672 40140 13084 40168
rect 4672 40128 4678 40140
rect 13078 40128 13084 40140
rect 13136 40128 13142 40180
rect 27430 40128 27436 40180
rect 27488 40168 27494 40180
rect 28353 40171 28411 40177
rect 28353 40168 28365 40171
rect 27488 40140 28365 40168
rect 27488 40128 27494 40140
rect 28353 40137 28365 40140
rect 28399 40137 28411 40171
rect 31110 40168 31116 40180
rect 31071 40140 31116 40168
rect 28353 40131 28411 40137
rect 31110 40128 31116 40140
rect 31168 40128 31174 40180
rect 32582 40168 32588 40180
rect 32140 40140 32588 40168
rect 2133 40103 2191 40109
rect 2133 40069 2145 40103
rect 2179 40100 2191 40103
rect 2866 40100 2872 40112
rect 2179 40072 2872 40100
rect 2179 40069 2191 40072
rect 2133 40063 2191 40069
rect 2866 40060 2872 40072
rect 2924 40060 2930 40112
rect 5626 40100 5632 40112
rect 4724 40072 5632 40100
rect 1946 40032 1952 40044
rect 1907 40004 1952 40032
rect 1946 39992 1952 40004
rect 2004 39992 2010 40044
rect 4724 40041 4752 40072
rect 5626 40060 5632 40072
rect 5684 40060 5690 40112
rect 12066 40100 12072 40112
rect 11992 40072 12072 40100
rect 11992 40041 12020 40072
rect 12066 40060 12072 40072
rect 12124 40060 12130 40112
rect 29822 40100 29828 40112
rect 29783 40072 29828 40100
rect 29822 40060 29828 40072
rect 29880 40060 29886 40112
rect 30041 40103 30099 40109
rect 30041 40069 30053 40103
rect 30087 40100 30099 40103
rect 31294 40100 31300 40112
rect 30087 40072 31300 40100
rect 30087 40069 30099 40072
rect 30041 40063 30099 40069
rect 31294 40060 31300 40072
rect 31352 40060 31358 40112
rect 32140 40109 32168 40140
rect 32582 40128 32588 40140
rect 32640 40128 32646 40180
rect 33410 40128 33416 40180
rect 33468 40168 33474 40180
rect 33505 40171 33563 40177
rect 33505 40168 33517 40171
rect 33468 40140 33517 40168
rect 33468 40128 33474 40140
rect 33505 40137 33517 40140
rect 33551 40137 33563 40171
rect 33505 40131 33563 40137
rect 37642 40128 37648 40180
rect 37700 40168 37706 40180
rect 38657 40171 38715 40177
rect 38657 40168 38669 40171
rect 37700 40140 38669 40168
rect 37700 40128 37706 40140
rect 38657 40137 38669 40140
rect 38703 40137 38715 40171
rect 38657 40131 38715 40137
rect 32125 40103 32183 40109
rect 32125 40069 32137 40103
rect 32171 40069 32183 40103
rect 32125 40063 32183 40069
rect 32341 40103 32399 40109
rect 32341 40069 32353 40103
rect 32387 40100 32399 40103
rect 33042 40100 33048 40112
rect 32387 40072 33048 40100
rect 32387 40069 32399 40072
rect 32341 40063 32399 40069
rect 33042 40060 33048 40072
rect 33100 40060 33106 40112
rect 33321 40103 33379 40109
rect 33321 40069 33333 40103
rect 33367 40100 33379 40103
rect 34514 40100 34520 40112
rect 33367 40072 34520 40100
rect 33367 40069 33379 40072
rect 33321 40063 33379 40069
rect 34514 40060 34520 40072
rect 34572 40060 34578 40112
rect 35250 40060 35256 40112
rect 35308 40100 35314 40112
rect 35630 40103 35688 40109
rect 35630 40100 35642 40103
rect 35308 40072 35642 40100
rect 35308 40060 35314 40072
rect 35630 40069 35642 40072
rect 35676 40069 35688 40103
rect 39482 40100 39488 40112
rect 39443 40072 39488 40100
rect 35630 40063 35688 40069
rect 39482 40060 39488 40072
rect 39540 40060 39546 40112
rect 40678 40060 40684 40112
rect 40736 40109 40742 40112
rect 40736 40103 40800 40109
rect 40736 40069 40754 40103
rect 40788 40069 40800 40103
rect 40736 40063 40800 40069
rect 40736 40060 40742 40063
rect 4709 40035 4767 40041
rect 4709 40001 4721 40035
rect 4755 40001 4767 40035
rect 4709 39995 4767 40001
rect 11977 40035 12035 40041
rect 11977 40001 11989 40035
rect 12023 40001 12035 40035
rect 11977 39995 12035 40001
rect 18960 40035 19018 40041
rect 18960 40001 18972 40035
rect 19006 40032 19018 40035
rect 19242 40032 19248 40044
rect 19006 40004 19248 40032
rect 19006 40001 19018 40004
rect 18960 39995 19018 40001
rect 19242 39992 19248 40004
rect 19300 39992 19306 40044
rect 20530 40032 20536 40044
rect 20491 40004 20536 40032
rect 20530 39992 20536 40004
rect 20588 39992 20594 40044
rect 24296 40035 24354 40041
rect 24296 40001 24308 40035
rect 24342 40032 24354 40035
rect 24578 40032 24584 40044
rect 24342 40004 24584 40032
rect 24342 40001 24354 40004
rect 24296 39995 24354 40001
rect 24578 39992 24584 40004
rect 24636 39992 24642 40044
rect 27062 39992 27068 40044
rect 27120 40032 27126 40044
rect 27229 40035 27287 40041
rect 27229 40032 27241 40035
rect 27120 40004 27241 40032
rect 27120 39992 27126 40004
rect 27229 40001 27241 40004
rect 27275 40001 27287 40035
rect 27229 39995 27287 40001
rect 30282 39992 30288 40044
rect 30340 40032 30346 40044
rect 30653 40035 30711 40041
rect 30653 40032 30665 40035
rect 30340 40004 30665 40032
rect 30340 39992 30346 40004
rect 30653 40001 30665 40004
rect 30699 40032 30711 40035
rect 30699 40004 31754 40032
rect 30699 40001 30711 40004
rect 30653 39995 30711 40001
rect 31726 39976 31754 40004
rect 37366 39992 37372 40044
rect 37424 40032 37430 40044
rect 37533 40035 37591 40041
rect 37533 40032 37545 40035
rect 37424 40004 37545 40032
rect 37424 39992 37430 40004
rect 37533 40001 37545 40004
rect 37579 40001 37591 40035
rect 37533 39995 37591 40001
rect 2774 39964 2780 39976
rect 2735 39936 2780 39964
rect 2774 39924 2780 39936
rect 2832 39924 2838 39976
rect 4614 39924 4620 39976
rect 4672 39964 4678 39976
rect 4893 39967 4951 39973
rect 4893 39964 4905 39967
rect 4672 39936 4905 39964
rect 4672 39924 4678 39936
rect 4893 39933 4905 39936
rect 4939 39933 4951 39967
rect 12158 39964 12164 39976
rect 12119 39936 12164 39964
rect 4893 39927 4951 39933
rect 12158 39924 12164 39936
rect 12216 39924 12222 39976
rect 16390 39924 16396 39976
rect 16448 39964 16454 39976
rect 18690 39964 18696 39976
rect 16448 39936 18696 39964
rect 16448 39924 16454 39936
rect 18690 39924 18696 39936
rect 18748 39924 18754 39976
rect 24029 39967 24087 39973
rect 24029 39933 24041 39967
rect 24075 39933 24087 39967
rect 26970 39964 26976 39976
rect 26931 39936 26976 39964
rect 24029 39927 24087 39933
rect 19978 39788 19984 39840
rect 20036 39828 20042 39840
rect 20073 39831 20131 39837
rect 20073 39828 20085 39831
rect 20036 39800 20085 39828
rect 20036 39788 20042 39800
rect 20073 39797 20085 39800
rect 20119 39797 20131 39831
rect 20714 39828 20720 39840
rect 20675 39800 20720 39828
rect 20073 39791 20131 39797
rect 20714 39788 20720 39800
rect 20772 39788 20778 39840
rect 24044 39828 24072 39927
rect 26970 39924 26976 39936
rect 27028 39924 27034 39976
rect 31726 39964 31760 39976
rect 31667 39936 31760 39964
rect 31754 39924 31760 39936
rect 31812 39964 31818 39976
rect 32306 39964 32312 39976
rect 31812 39936 32312 39964
rect 31812 39924 31818 39936
rect 32306 39924 32312 39936
rect 32364 39924 32370 39976
rect 35897 39967 35955 39973
rect 35897 39933 35909 39967
rect 35943 39964 35955 39967
rect 36078 39964 36084 39976
rect 35943 39936 36084 39964
rect 35943 39933 35955 39936
rect 35897 39927 35955 39933
rect 36078 39924 36084 39936
rect 36136 39964 36142 39976
rect 37277 39967 37335 39973
rect 37277 39964 37289 39967
rect 36136 39936 37289 39964
rect 36136 39924 36142 39936
rect 37277 39933 37289 39936
rect 37323 39933 37335 39967
rect 39942 39964 39948 39976
rect 37277 39927 37335 39933
rect 38304 39936 39948 39964
rect 26988 39896 27016 39924
rect 24964 39868 27016 39896
rect 31021 39899 31079 39905
rect 24302 39828 24308 39840
rect 24044 39800 24308 39828
rect 24302 39788 24308 39800
rect 24360 39828 24366 39840
rect 24964 39828 24992 39868
rect 31021 39865 31033 39899
rect 31067 39896 31079 39899
rect 31478 39896 31484 39908
rect 31067 39868 31484 39896
rect 31067 39865 31079 39868
rect 31021 39859 31079 39865
rect 31478 39856 31484 39868
rect 31536 39856 31542 39908
rect 32493 39899 32551 39905
rect 32493 39865 32505 39899
rect 32539 39896 32551 39899
rect 32950 39896 32956 39908
rect 32539 39868 32956 39896
rect 32539 39865 32551 39868
rect 32493 39859 32551 39865
rect 32950 39856 32956 39868
rect 33008 39856 33014 39908
rect 24360 39800 24992 39828
rect 24360 39788 24366 39800
rect 25314 39788 25320 39840
rect 25372 39828 25378 39840
rect 25409 39831 25467 39837
rect 25409 39828 25421 39831
rect 25372 39800 25421 39828
rect 25372 39788 25378 39800
rect 25409 39797 25421 39800
rect 25455 39797 25467 39831
rect 30006 39828 30012 39840
rect 29967 39800 30012 39828
rect 25409 39791 25467 39797
rect 30006 39788 30012 39800
rect 30064 39788 30070 39840
rect 30098 39788 30104 39840
rect 30156 39828 30162 39840
rect 30193 39831 30251 39837
rect 30193 39828 30205 39831
rect 30156 39800 30205 39828
rect 30156 39788 30162 39800
rect 30193 39797 30205 39800
rect 30239 39797 30251 39831
rect 32306 39828 32312 39840
rect 32267 39800 32312 39828
rect 30193 39791 30251 39797
rect 32306 39788 32312 39800
rect 32364 39788 32370 39840
rect 33318 39828 33324 39840
rect 33279 39800 33324 39828
rect 33318 39788 33324 39800
rect 33376 39788 33382 39840
rect 33962 39788 33968 39840
rect 34020 39828 34026 39840
rect 34517 39831 34575 39837
rect 34517 39828 34529 39831
rect 34020 39800 34529 39828
rect 34020 39788 34026 39800
rect 34517 39797 34529 39800
rect 34563 39797 34575 39831
rect 37292 39828 37320 39927
rect 38304 39828 38332 39936
rect 39942 39924 39948 39936
rect 40000 39964 40006 39976
rect 40497 39967 40555 39973
rect 40497 39964 40509 39967
rect 40000 39936 40509 39964
rect 40000 39924 40006 39936
rect 40497 39933 40509 39936
rect 40543 39933 40555 39967
rect 40497 39927 40555 39933
rect 38930 39856 38936 39908
rect 38988 39896 38994 39908
rect 39117 39899 39175 39905
rect 39117 39896 39129 39899
rect 38988 39868 39129 39896
rect 38988 39856 38994 39868
rect 39117 39865 39129 39868
rect 39163 39865 39175 39899
rect 39117 39859 39175 39865
rect 39669 39899 39727 39905
rect 39669 39865 39681 39899
rect 39715 39896 39727 39899
rect 40034 39896 40040 39908
rect 39715 39868 40040 39896
rect 39715 39865 39727 39868
rect 39669 39859 39727 39865
rect 40034 39856 40040 39868
rect 40092 39856 40098 39908
rect 37292 39800 38332 39828
rect 34517 39791 34575 39797
rect 39390 39788 39396 39840
rect 39448 39828 39454 39840
rect 39485 39831 39543 39837
rect 39485 39828 39497 39831
rect 39448 39800 39497 39828
rect 39448 39788 39454 39800
rect 39485 39797 39497 39800
rect 39531 39797 39543 39831
rect 41874 39828 41880 39840
rect 41835 39800 41880 39828
rect 39485 39791 39543 39797
rect 41874 39788 41880 39800
rect 41932 39788 41938 39840
rect 43809 39831 43867 39837
rect 43809 39797 43821 39831
rect 43855 39828 43867 39831
rect 44174 39828 44180 39840
rect 43855 39800 44180 39828
rect 43855 39797 43867 39800
rect 43809 39791 43867 39797
rect 44174 39788 44180 39800
rect 44232 39788 44238 39840
rect 1104 39738 44896 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 44896 39738
rect 1104 39664 44896 39686
rect 2866 39624 2872 39636
rect 2827 39596 2872 39624
rect 2866 39584 2872 39596
rect 2924 39584 2930 39636
rect 3786 39624 3792 39636
rect 3747 39596 3792 39624
rect 3786 39584 3792 39596
rect 3844 39584 3850 39636
rect 19242 39624 19248 39636
rect 19203 39596 19248 39624
rect 19242 39584 19248 39596
rect 19300 39584 19306 39636
rect 24578 39624 24584 39636
rect 24539 39596 24584 39624
rect 24578 39584 24584 39596
rect 24636 39584 24642 39636
rect 27062 39624 27068 39636
rect 27023 39596 27068 39624
rect 27062 39584 27068 39596
rect 27120 39584 27126 39636
rect 28902 39624 28908 39636
rect 28863 39596 28908 39624
rect 28902 39584 28908 39596
rect 28960 39584 28966 39636
rect 32122 39624 32128 39636
rect 32083 39596 32128 39624
rect 32122 39584 32128 39596
rect 32180 39584 32186 39636
rect 34149 39627 34207 39633
rect 34149 39593 34161 39627
rect 34195 39624 34207 39627
rect 35069 39627 35127 39633
rect 35069 39624 35081 39627
rect 34195 39596 35081 39624
rect 34195 39593 34207 39596
rect 34149 39587 34207 39593
rect 35069 39593 35081 39596
rect 35115 39593 35127 39627
rect 35069 39587 35127 39593
rect 35253 39627 35311 39633
rect 35253 39593 35265 39627
rect 35299 39624 35311 39627
rect 35342 39624 35348 39636
rect 35299 39596 35348 39624
rect 35299 39593 35311 39596
rect 35253 39587 35311 39593
rect 35342 39584 35348 39596
rect 35400 39584 35406 39636
rect 37274 39584 37280 39636
rect 37332 39624 37338 39636
rect 37369 39627 37427 39633
rect 37369 39624 37381 39627
rect 37332 39596 37381 39624
rect 37332 39584 37338 39596
rect 37369 39593 37381 39596
rect 37415 39593 37427 39627
rect 38930 39624 38936 39636
rect 38891 39596 38936 39624
rect 37369 39587 37427 39593
rect 38930 39584 38936 39596
rect 38988 39584 38994 39636
rect 39117 39627 39175 39633
rect 39117 39593 39129 39627
rect 39163 39624 39175 39627
rect 39206 39624 39212 39636
rect 39163 39596 39212 39624
rect 39163 39593 39175 39596
rect 39117 39587 39175 39593
rect 39206 39584 39212 39596
rect 39264 39584 39270 39636
rect 39482 39584 39488 39636
rect 39540 39624 39546 39636
rect 39853 39627 39911 39633
rect 39853 39624 39865 39627
rect 39540 39596 39865 39624
rect 39540 39584 39546 39596
rect 39853 39593 39865 39596
rect 39899 39593 39911 39627
rect 39853 39587 39911 39593
rect 40770 39584 40776 39636
rect 40828 39624 40834 39636
rect 40865 39627 40923 39633
rect 40865 39624 40877 39627
rect 40828 39596 40877 39624
rect 40828 39584 40834 39596
rect 40865 39593 40877 39596
rect 40911 39593 40923 39627
rect 40865 39587 40923 39593
rect 32582 39516 32588 39568
rect 32640 39556 32646 39568
rect 32677 39559 32735 39565
rect 32677 39556 32689 39559
rect 32640 39528 32689 39556
rect 32640 39516 32646 39528
rect 32677 39525 32689 39528
rect 32723 39525 32735 39559
rect 32677 39519 32735 39525
rect 34514 39516 34520 39568
rect 34572 39556 34578 39568
rect 39390 39556 39396 39568
rect 34572 39528 39396 39556
rect 34572 39516 34578 39528
rect 39390 39516 39396 39528
rect 39448 39516 39454 39568
rect 40957 39559 41015 39565
rect 40957 39525 40969 39559
rect 41003 39556 41015 39559
rect 41046 39556 41052 39568
rect 41003 39528 41052 39556
rect 41003 39525 41015 39528
rect 40957 39519 41015 39525
rect 10134 39488 10140 39500
rect 2976 39460 10140 39488
rect 2976 39429 3004 39460
rect 10134 39448 10140 39460
rect 10192 39448 10198 39500
rect 18690 39448 18696 39500
rect 18748 39488 18754 39500
rect 20441 39491 20499 39497
rect 20441 39488 20453 39491
rect 18748 39460 20453 39488
rect 18748 39448 18754 39460
rect 20441 39457 20453 39460
rect 20487 39457 20499 39491
rect 20441 39451 20499 39457
rect 25961 39491 26019 39497
rect 25961 39457 25973 39491
rect 26007 39488 26019 39491
rect 26418 39488 26424 39500
rect 26007 39460 26424 39488
rect 26007 39457 26019 39460
rect 25961 39451 26019 39457
rect 2961 39423 3019 39429
rect 2961 39389 2973 39423
rect 3007 39389 3019 39423
rect 4798 39420 4804 39432
rect 4759 39392 4804 39420
rect 2961 39383 3019 39389
rect 4798 39380 4804 39392
rect 4856 39380 4862 39432
rect 5626 39420 5632 39432
rect 5587 39392 5632 39420
rect 5626 39380 5632 39392
rect 5684 39380 5690 39432
rect 19429 39423 19487 39429
rect 19429 39389 19441 39423
rect 19475 39389 19487 39423
rect 19429 39383 19487 39389
rect 19521 39423 19579 39429
rect 19521 39389 19533 39423
rect 19567 39420 19579 39423
rect 19978 39420 19984 39432
rect 19567 39392 19984 39420
rect 19567 39389 19579 39392
rect 19521 39383 19579 39389
rect 19444 39352 19472 39383
rect 19978 39380 19984 39392
rect 20036 39380 20042 39432
rect 20456 39420 20484 39451
rect 26418 39448 26424 39460
rect 26476 39448 26482 39500
rect 26789 39491 26847 39497
rect 26789 39457 26801 39491
rect 26835 39488 26847 39491
rect 27430 39488 27436 39500
rect 26835 39460 27436 39488
rect 26835 39457 26847 39460
rect 26789 39451 26847 39457
rect 27430 39448 27436 39460
rect 27488 39448 27494 39500
rect 30742 39488 30748 39500
rect 30703 39460 30748 39488
rect 30742 39448 30748 39460
rect 30800 39448 30806 39500
rect 37277 39491 37335 39497
rect 37277 39488 37289 39491
rect 31772 39460 37289 39488
rect 21634 39420 21640 39432
rect 20456 39392 21640 39420
rect 21634 39380 21640 39392
rect 21692 39380 21698 39432
rect 22922 39380 22928 39432
rect 22980 39420 22986 39432
rect 24397 39423 24455 39429
rect 24397 39420 24409 39423
rect 22980 39392 24409 39420
rect 22980 39380 22986 39392
rect 24397 39389 24409 39392
rect 24443 39389 24455 39423
rect 24397 39383 24455 39389
rect 24673 39423 24731 39429
rect 24673 39389 24685 39423
rect 24719 39420 24731 39423
rect 25498 39420 25504 39432
rect 24719 39392 25504 39420
rect 24719 39389 24731 39392
rect 24673 39383 24731 39389
rect 25498 39380 25504 39392
rect 25556 39380 25562 39432
rect 25590 39380 25596 39432
rect 25648 39420 25654 39432
rect 25777 39423 25835 39429
rect 25648 39392 25693 39420
rect 25648 39380 25654 39392
rect 25777 39389 25789 39423
rect 25823 39389 25835 39423
rect 26878 39420 26884 39432
rect 26839 39392 26884 39420
rect 25777 39383 25835 39389
rect 20438 39352 20444 39364
rect 19444 39324 20444 39352
rect 20438 39312 20444 39324
rect 20496 39312 20502 39364
rect 20714 39361 20720 39364
rect 20708 39352 20720 39361
rect 20675 39324 20720 39352
rect 20708 39315 20720 39324
rect 20714 39312 20720 39315
rect 20772 39312 20778 39364
rect 24486 39352 24492 39364
rect 24447 39324 24492 39352
rect 24486 39312 24492 39324
rect 24544 39312 24550 39364
rect 25406 39312 25412 39364
rect 25464 39352 25470 39364
rect 25792 39352 25820 39383
rect 26878 39380 26884 39392
rect 26936 39380 26942 39432
rect 26970 39380 26976 39432
rect 27028 39420 27034 39432
rect 27525 39423 27583 39429
rect 27525 39420 27537 39423
rect 27028 39392 27537 39420
rect 27028 39380 27034 39392
rect 27525 39389 27537 39392
rect 27571 39420 27583 39423
rect 29454 39420 29460 39432
rect 27571 39392 29460 39420
rect 27571 39389 27583 39392
rect 27525 39383 27583 39389
rect 29454 39380 29460 39392
rect 29512 39380 29518 39432
rect 30282 39420 30288 39432
rect 30243 39392 30288 39420
rect 30282 39380 30288 39392
rect 30340 39380 30346 39432
rect 31018 39429 31024 39432
rect 31012 39420 31024 39429
rect 30979 39392 31024 39420
rect 31012 39383 31024 39392
rect 31018 39380 31024 39383
rect 31076 39380 31082 39432
rect 31478 39380 31484 39432
rect 31536 39420 31542 39432
rect 31772 39420 31800 39460
rect 37277 39457 37289 39460
rect 37323 39457 37335 39491
rect 37277 39451 37335 39457
rect 37461 39491 37519 39497
rect 37461 39457 37473 39491
rect 37507 39488 37519 39491
rect 37734 39488 37740 39500
rect 37507 39460 37740 39488
rect 37507 39457 37519 39460
rect 37461 39451 37519 39457
rect 31536 39392 31800 39420
rect 31536 39380 31542 39392
rect 32122 39380 32128 39432
rect 32180 39420 32186 39432
rect 32861 39423 32919 39429
rect 32861 39420 32873 39423
rect 32180 39392 32873 39420
rect 32180 39380 32186 39392
rect 32861 39389 32873 39392
rect 32907 39389 32919 39423
rect 32861 39383 32919 39389
rect 32950 39380 32956 39432
rect 33008 39420 33014 39432
rect 33781 39423 33839 39429
rect 33781 39420 33793 39423
rect 33008 39392 33793 39420
rect 33008 39380 33014 39392
rect 33781 39389 33793 39392
rect 33827 39389 33839 39423
rect 33962 39420 33968 39432
rect 33923 39392 33968 39420
rect 33781 39383 33839 39389
rect 33962 39380 33968 39392
rect 34020 39380 34026 39432
rect 34698 39420 34704 39432
rect 34659 39392 34704 39420
rect 34698 39380 34704 39392
rect 34756 39380 34762 39432
rect 25464 39324 25820 39352
rect 27792 39355 27850 39361
rect 25464 39312 25470 39324
rect 27792 39321 27804 39355
rect 27838 39352 27850 39355
rect 27890 39352 27896 39364
rect 27838 39324 27896 39352
rect 27838 39321 27850 39324
rect 27792 39315 27850 39321
rect 27890 39312 27896 39324
rect 27948 39312 27954 39364
rect 30101 39355 30159 39361
rect 30101 39321 30113 39355
rect 30147 39352 30159 39355
rect 30834 39352 30840 39364
rect 30147 39324 30840 39352
rect 30147 39321 30159 39324
rect 30101 39315 30159 39321
rect 30834 39312 30840 39324
rect 30892 39312 30898 39364
rect 33318 39352 33324 39364
rect 32968 39324 33324 39352
rect 19889 39287 19947 39293
rect 19889 39253 19901 39287
rect 19935 39284 19947 39287
rect 20070 39284 20076 39296
rect 19935 39256 20076 39284
rect 19935 39253 19947 39256
rect 19889 39247 19947 39253
rect 20070 39244 20076 39256
rect 20128 39244 20134 39296
rect 20806 39244 20812 39296
rect 20864 39284 20870 39296
rect 21821 39287 21879 39293
rect 21821 39284 21833 39287
rect 20864 39256 21833 39284
rect 20864 39244 20870 39256
rect 21821 39253 21833 39256
rect 21867 39253 21879 39287
rect 21821 39247 21879 39253
rect 29917 39287 29975 39293
rect 29917 39253 29929 39287
rect 29963 39284 29975 39287
rect 30006 39284 30012 39296
rect 29963 39256 30012 39284
rect 29963 39253 29975 39256
rect 29917 39247 29975 39253
rect 30006 39244 30012 39256
rect 30064 39284 30070 39296
rect 31846 39284 31852 39296
rect 30064 39256 31852 39284
rect 30064 39244 30070 39256
rect 31846 39244 31852 39256
rect 31904 39244 31910 39296
rect 32968 39293 32996 39324
rect 33318 39312 33324 39324
rect 33376 39352 33382 39364
rect 33980 39352 34008 39380
rect 33376 39324 34008 39352
rect 33376 39312 33382 39324
rect 32953 39287 33011 39293
rect 32953 39253 32965 39287
rect 32999 39253 33011 39287
rect 32953 39247 33011 39253
rect 33042 39244 33048 39296
rect 33100 39284 33106 39296
rect 33226 39284 33232 39296
rect 33100 39256 33145 39284
rect 33187 39256 33232 39284
rect 33100 39244 33106 39256
rect 33226 39244 33232 39256
rect 33284 39244 33290 39296
rect 34514 39244 34520 39296
rect 34572 39284 34578 39296
rect 35069 39287 35127 39293
rect 35069 39284 35081 39287
rect 34572 39256 35081 39284
rect 34572 39244 34578 39256
rect 35069 39253 35081 39256
rect 35115 39253 35127 39287
rect 37292 39284 37320 39451
rect 37734 39448 37740 39460
rect 37792 39448 37798 39500
rect 40770 39488 40776 39500
rect 39132 39460 40356 39488
rect 40731 39460 40776 39488
rect 37553 39423 37611 39429
rect 37553 39389 37565 39423
rect 37599 39420 37611 39423
rect 37642 39420 37648 39432
rect 37599 39392 37648 39420
rect 37599 39389 37611 39392
rect 37553 39383 37611 39389
rect 37642 39380 37648 39392
rect 37700 39380 37706 39432
rect 39132 39361 39160 39460
rect 39206 39380 39212 39432
rect 39264 39420 39270 39432
rect 39666 39420 39672 39432
rect 39264 39392 39672 39420
rect 39264 39380 39270 39392
rect 39666 39380 39672 39392
rect 39724 39420 39730 39432
rect 40328 39429 40356 39460
rect 40770 39448 40776 39460
rect 40828 39448 40834 39500
rect 40037 39423 40095 39429
rect 40037 39420 40049 39423
rect 39724 39392 40049 39420
rect 39724 39380 39730 39392
rect 40037 39389 40049 39392
rect 40083 39389 40095 39423
rect 40037 39383 40095 39389
rect 40313 39423 40371 39429
rect 40313 39389 40325 39423
rect 40359 39420 40371 39423
rect 40494 39420 40500 39432
rect 40359 39392 40500 39420
rect 40359 39389 40371 39392
rect 40313 39383 40371 39389
rect 40494 39380 40500 39392
rect 40552 39420 40558 39432
rect 40972 39420 41000 39519
rect 41046 39516 41052 39528
rect 41104 39516 41110 39568
rect 42702 39488 42708 39500
rect 42663 39460 42708 39488
rect 42702 39448 42708 39460
rect 42760 39448 42766 39500
rect 44174 39488 44180 39500
rect 44135 39460 44180 39488
rect 44174 39448 44180 39460
rect 44232 39448 44238 39500
rect 40552 39392 41000 39420
rect 41049 39423 41107 39429
rect 40552 39380 40558 39392
rect 41049 39389 41061 39423
rect 41095 39389 41107 39423
rect 41049 39383 41107 39389
rect 41693 39423 41751 39429
rect 41693 39389 41705 39423
rect 41739 39420 41751 39423
rect 41874 39420 41880 39432
rect 41739 39392 41880 39420
rect 41739 39389 41751 39392
rect 41693 39383 41751 39389
rect 39101 39355 39160 39361
rect 39101 39321 39113 39355
rect 39147 39324 39160 39355
rect 39298 39352 39304 39364
rect 39259 39324 39304 39352
rect 39147 39321 39159 39324
rect 39101 39315 39159 39321
rect 39298 39312 39304 39324
rect 39356 39352 39362 39364
rect 40221 39355 40279 39361
rect 40221 39352 40233 39355
rect 39356 39324 40233 39352
rect 39356 39312 39362 39324
rect 40221 39321 40233 39324
rect 40267 39352 40279 39355
rect 40586 39352 40592 39364
rect 40267 39324 40592 39352
rect 40267 39321 40279 39324
rect 40221 39315 40279 39321
rect 40586 39312 40592 39324
rect 40644 39352 40650 39364
rect 41064 39352 41092 39383
rect 41874 39380 41880 39392
rect 41932 39380 41938 39432
rect 40644 39324 41414 39352
rect 40644 39312 40650 39324
rect 37550 39284 37556 39296
rect 37292 39256 37556 39284
rect 35069 39247 35127 39253
rect 37550 39244 37556 39256
rect 37608 39284 37614 39296
rect 40770 39284 40776 39296
rect 37608 39256 40776 39284
rect 37608 39244 37614 39256
rect 40770 39244 40776 39256
rect 40828 39244 40834 39296
rect 41386 39284 41414 39324
rect 43438 39312 43444 39364
rect 43496 39352 43502 39364
rect 43993 39355 44051 39361
rect 43993 39352 44005 39355
rect 43496 39324 44005 39352
rect 43496 39312 43502 39324
rect 43993 39321 44005 39324
rect 44039 39321 44051 39355
rect 43993 39315 44051 39321
rect 41509 39287 41567 39293
rect 41509 39284 41521 39287
rect 41386 39256 41521 39284
rect 41509 39253 41521 39256
rect 41555 39253 41567 39287
rect 41509 39247 41567 39253
rect 1104 39194 44896 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 44896 39194
rect 1104 39120 44896 39142
rect 20349 39083 20407 39089
rect 20349 39049 20361 39083
rect 20395 39080 20407 39083
rect 20530 39080 20536 39092
rect 20395 39052 20536 39080
rect 20395 39049 20407 39052
rect 20349 39043 20407 39049
rect 20530 39040 20536 39052
rect 20588 39040 20594 39092
rect 24486 39040 24492 39092
rect 24544 39080 24550 39092
rect 24673 39083 24731 39089
rect 24673 39080 24685 39083
rect 24544 39052 24685 39080
rect 24544 39040 24550 39052
rect 24673 39049 24685 39052
rect 24719 39049 24731 39083
rect 24673 39043 24731 39049
rect 26329 39083 26387 39089
rect 26329 39049 26341 39083
rect 26375 39080 26387 39083
rect 26878 39080 26884 39092
rect 26375 39052 26884 39080
rect 26375 39049 26387 39052
rect 26329 39043 26387 39049
rect 26878 39040 26884 39052
rect 26936 39040 26942 39092
rect 27890 39080 27896 39092
rect 27851 39052 27896 39080
rect 27890 39040 27896 39052
rect 27948 39040 27954 39092
rect 30834 39080 30840 39092
rect 30795 39052 30840 39080
rect 30834 39040 30840 39052
rect 30892 39040 30898 39092
rect 31294 39080 31300 39092
rect 31255 39052 31300 39080
rect 31294 39040 31300 39052
rect 31352 39040 31358 39092
rect 43438 39080 43444 39092
rect 35866 39052 41414 39080
rect 43399 39052 43444 39080
rect 25406 39012 25412 39024
rect 19352 38984 25412 39012
rect 16853 38947 16911 38953
rect 16853 38913 16865 38947
rect 16899 38913 16911 38947
rect 16853 38907 16911 38913
rect 16758 38836 16764 38888
rect 16816 38876 16822 38888
rect 16868 38876 16896 38907
rect 16942 38904 16948 38956
rect 17000 38944 17006 38956
rect 17129 38947 17187 38953
rect 17000 38916 17045 38944
rect 17000 38904 17006 38916
rect 17129 38913 17141 38947
rect 17175 38944 17187 38947
rect 18414 38944 18420 38956
rect 17175 38916 18420 38944
rect 17175 38913 17187 38916
rect 17129 38907 17187 38913
rect 18414 38904 18420 38916
rect 18472 38944 18478 38956
rect 19352 38953 19380 38984
rect 25406 38972 25412 38984
rect 25464 38972 25470 39024
rect 25590 38972 25596 39024
rect 25648 39012 25654 39024
rect 26973 39015 27031 39021
rect 26973 39012 26985 39015
rect 25648 38984 26985 39012
rect 25648 38972 25654 38984
rect 26973 38981 26985 38984
rect 27019 38981 27031 39015
rect 26973 38975 27031 38981
rect 28166 38972 28172 39024
rect 28224 39012 28230 39024
rect 28224 38984 30512 39012
rect 28224 38972 28230 38984
rect 19061 38947 19119 38953
rect 19061 38944 19073 38947
rect 18472 38916 19073 38944
rect 18472 38904 18478 38916
rect 19061 38913 19073 38916
rect 19107 38913 19119 38947
rect 19061 38907 19119 38913
rect 19337 38947 19395 38953
rect 19337 38913 19349 38947
rect 19383 38913 19395 38947
rect 19337 38907 19395 38913
rect 19521 38947 19579 38953
rect 19521 38913 19533 38947
rect 19567 38944 19579 38947
rect 20070 38944 20076 38956
rect 19567 38916 20076 38944
rect 19567 38913 19579 38916
rect 19521 38907 19579 38913
rect 20070 38904 20076 38916
rect 20128 38944 20134 38956
rect 22186 38953 22192 38956
rect 20165 38947 20223 38953
rect 20165 38944 20177 38947
rect 20128 38916 20177 38944
rect 20128 38904 20134 38916
rect 20165 38913 20177 38916
rect 20211 38913 20223 38947
rect 20165 38907 20223 38913
rect 22180 38907 22192 38953
rect 22244 38944 22250 38956
rect 24394 38944 24400 38956
rect 22244 38916 22280 38944
rect 24355 38916 24400 38944
rect 22186 38904 22192 38907
rect 22244 38904 22250 38916
rect 24394 38904 24400 38916
rect 24452 38944 24458 38956
rect 25133 38947 25191 38953
rect 25133 38944 25145 38947
rect 24452 38916 25145 38944
rect 24452 38904 24458 38916
rect 25133 38913 25145 38916
rect 25179 38913 25191 38947
rect 25314 38944 25320 38956
rect 25275 38916 25320 38944
rect 25133 38907 25191 38913
rect 25314 38904 25320 38916
rect 25372 38904 25378 38956
rect 25501 38947 25559 38953
rect 25501 38913 25513 38947
rect 25547 38944 25559 38947
rect 25866 38944 25872 38956
rect 25547 38916 25872 38944
rect 25547 38913 25559 38916
rect 25501 38907 25559 38913
rect 25866 38904 25872 38916
rect 25924 38944 25930 38956
rect 25961 38947 26019 38953
rect 25961 38944 25973 38947
rect 25924 38916 25973 38944
rect 25924 38904 25930 38916
rect 25961 38913 25973 38916
rect 26007 38913 26019 38947
rect 27154 38944 27160 38956
rect 27115 38916 27160 38944
rect 25961 38907 26019 38913
rect 27154 38904 27160 38916
rect 27212 38904 27218 38956
rect 28074 38944 28080 38956
rect 28035 38916 28080 38944
rect 28074 38904 28080 38916
rect 28132 38904 28138 38956
rect 29454 38944 29460 38956
rect 29415 38916 29460 38944
rect 29454 38904 29460 38916
rect 29512 38904 29518 38956
rect 29730 38953 29736 38956
rect 29724 38907 29736 38953
rect 29788 38944 29794 38956
rect 29788 38916 29824 38944
rect 29730 38904 29736 38907
rect 29788 38904 29794 38916
rect 19981 38879 20039 38885
rect 16816 38848 19472 38876
rect 16816 38836 16822 38848
rect 16850 38740 16856 38752
rect 16811 38712 16856 38740
rect 16850 38700 16856 38712
rect 16908 38700 16914 38752
rect 19153 38743 19211 38749
rect 19153 38709 19165 38743
rect 19199 38740 19211 38743
rect 19334 38740 19340 38752
rect 19199 38712 19340 38740
rect 19199 38709 19211 38712
rect 19153 38703 19211 38709
rect 19334 38700 19340 38712
rect 19392 38700 19398 38752
rect 19444 38740 19472 38848
rect 19981 38845 19993 38879
rect 20027 38876 20039 38879
rect 20806 38876 20812 38888
rect 20027 38848 20812 38876
rect 20027 38845 20039 38848
rect 19981 38839 20039 38845
rect 20806 38836 20812 38848
rect 20864 38836 20870 38888
rect 21634 38836 21640 38888
rect 21692 38876 21698 38888
rect 21913 38879 21971 38885
rect 21913 38876 21925 38879
rect 21692 38848 21925 38876
rect 21692 38836 21698 38848
rect 21913 38845 21925 38848
rect 21959 38845 21971 38879
rect 21913 38839 21971 38845
rect 24673 38879 24731 38885
rect 24673 38845 24685 38879
rect 24719 38876 24731 38879
rect 25332 38876 25360 38904
rect 24719 38848 25360 38876
rect 26053 38879 26111 38885
rect 24719 38845 24731 38848
rect 24673 38839 24731 38845
rect 26053 38845 26065 38879
rect 26099 38845 26111 38879
rect 27430 38876 27436 38888
rect 27391 38848 27436 38876
rect 26053 38839 26111 38845
rect 23293 38811 23351 38817
rect 23293 38777 23305 38811
rect 23339 38808 23351 38811
rect 26068 38808 26096 38839
rect 27430 38836 27436 38848
rect 27488 38836 27494 38888
rect 30484 38876 30512 38984
rect 30852 38944 30880 39040
rect 32582 39012 32588 39024
rect 31312 38984 32588 39012
rect 31312 38953 31340 38984
rect 32582 38972 32588 38984
rect 32640 38972 32646 39024
rect 32861 39015 32919 39021
rect 32861 38981 32873 39015
rect 32907 39012 32919 39015
rect 33410 39012 33416 39024
rect 32907 38984 33416 39012
rect 32907 38981 32919 38984
rect 32861 38975 32919 38981
rect 33410 38972 33416 38984
rect 33468 38972 33474 39024
rect 31297 38947 31355 38953
rect 31297 38944 31309 38947
rect 30852 38916 31309 38944
rect 31297 38913 31309 38916
rect 31343 38913 31355 38947
rect 31297 38907 31355 38913
rect 31481 38947 31539 38953
rect 31481 38913 31493 38947
rect 31527 38944 31539 38947
rect 31754 38944 31760 38956
rect 31527 38916 31760 38944
rect 31527 38913 31539 38916
rect 31481 38907 31539 38913
rect 31754 38904 31760 38916
rect 31812 38904 31818 38956
rect 31846 38904 31852 38956
rect 31904 38944 31910 38956
rect 33137 38947 33195 38953
rect 33137 38944 33149 38947
rect 31904 38916 33149 38944
rect 31904 38904 31910 38916
rect 33137 38913 33149 38916
rect 33183 38913 33195 38947
rect 33318 38944 33324 38956
rect 33279 38916 33324 38944
rect 33137 38907 33195 38913
rect 33318 38904 33324 38916
rect 33376 38904 33382 38956
rect 34054 38944 34060 38956
rect 34015 38916 34060 38944
rect 34054 38904 34060 38916
rect 34112 38904 34118 38956
rect 35866 38876 35894 39052
rect 39761 39015 39819 39021
rect 39761 39012 39773 39015
rect 38856 38984 39773 39012
rect 38856 38956 38884 38984
rect 39761 38981 39773 38984
rect 39807 38981 39819 39015
rect 39761 38975 39819 38981
rect 36725 38947 36783 38953
rect 36725 38913 36737 38947
rect 36771 38944 36783 38947
rect 37274 38944 37280 38956
rect 36771 38916 37280 38944
rect 36771 38913 36783 38916
rect 36725 38907 36783 38913
rect 37274 38904 37280 38916
rect 37332 38904 37338 38956
rect 37366 38904 37372 38956
rect 37424 38944 37430 38956
rect 37461 38947 37519 38953
rect 37461 38944 37473 38947
rect 37424 38916 37473 38944
rect 37424 38904 37430 38916
rect 37461 38913 37473 38916
rect 37507 38913 37519 38947
rect 37642 38944 37648 38956
rect 37603 38916 37648 38944
rect 37461 38907 37519 38913
rect 37642 38904 37648 38916
rect 37700 38904 37706 38956
rect 37734 38904 37740 38956
rect 37792 38944 37798 38956
rect 38838 38944 38844 38956
rect 37792 38916 37837 38944
rect 38751 38916 38844 38944
rect 37792 38904 37798 38916
rect 38838 38904 38844 38916
rect 38896 38904 38902 38956
rect 38930 38904 38936 38956
rect 38988 38944 38994 38956
rect 38988 38916 39033 38944
rect 38988 38904 38994 38916
rect 39298 38904 39304 38956
rect 39356 38944 39362 38956
rect 39577 38947 39635 38953
rect 39577 38944 39589 38947
rect 39356 38916 39589 38944
rect 39356 38904 39362 38916
rect 39577 38913 39589 38916
rect 39623 38913 39635 38947
rect 39577 38907 39635 38913
rect 39666 38904 39672 38956
rect 39724 38944 39730 38956
rect 39853 38947 39911 38953
rect 39853 38944 39865 38947
rect 39724 38916 39865 38944
rect 39724 38904 39730 38916
rect 39853 38913 39865 38916
rect 39899 38913 39911 38947
rect 39853 38907 39911 38913
rect 39945 38947 40003 38953
rect 39945 38913 39957 38947
rect 39991 38913 40003 38947
rect 41386 38944 41414 39052
rect 43438 39040 43444 39052
rect 43496 39040 43502 39092
rect 43162 38944 43168 38956
rect 41386 38916 43168 38944
rect 39945 38907 40003 38913
rect 39114 38876 39120 38888
rect 30484 38848 35894 38876
rect 39075 38848 39120 38876
rect 39114 38836 39120 38848
rect 39172 38836 39178 38888
rect 39960 38876 39988 38907
rect 43162 38904 43168 38916
rect 43220 38944 43226 38956
rect 43349 38947 43407 38953
rect 43349 38944 43361 38947
rect 43220 38916 43361 38944
rect 43220 38904 43226 38916
rect 43349 38913 43361 38916
rect 43395 38913 43407 38947
rect 43349 38907 43407 38913
rect 40770 38876 40776 38888
rect 39960 38848 40776 38876
rect 40770 38836 40776 38848
rect 40828 38836 40834 38888
rect 41046 38876 41052 38888
rect 41007 38848 41052 38876
rect 41046 38836 41052 38848
rect 41104 38836 41110 38888
rect 27341 38811 27399 38817
rect 27341 38808 27353 38811
rect 23339 38780 27353 38808
rect 23339 38777 23351 38780
rect 23293 38771 23351 38777
rect 27341 38777 27353 38780
rect 27387 38808 27399 38811
rect 27798 38808 27804 38820
rect 27387 38780 27804 38808
rect 27387 38777 27399 38780
rect 27341 38771 27399 38777
rect 27798 38768 27804 38780
rect 27856 38768 27862 38820
rect 37734 38768 37740 38820
rect 37792 38808 37798 38820
rect 40034 38808 40040 38820
rect 37792 38780 40040 38808
rect 37792 38768 37798 38780
rect 40034 38768 40040 38780
rect 40092 38808 40098 38820
rect 40129 38811 40187 38817
rect 40129 38808 40141 38811
rect 40092 38780 40141 38808
rect 40092 38768 40098 38780
rect 40129 38777 40141 38780
rect 40175 38777 40187 38811
rect 40129 38771 40187 38777
rect 22922 38740 22928 38752
rect 19444 38712 22928 38740
rect 22922 38700 22928 38712
rect 22980 38700 22986 38752
rect 24489 38743 24547 38749
rect 24489 38709 24501 38743
rect 24535 38740 24547 38743
rect 25038 38740 25044 38752
rect 24535 38712 25044 38740
rect 24535 38709 24547 38712
rect 24489 38703 24547 38709
rect 25038 38700 25044 38712
rect 25096 38740 25102 38752
rect 25961 38743 26019 38749
rect 25961 38740 25973 38743
rect 25096 38712 25973 38740
rect 25096 38700 25102 38712
rect 25961 38709 25973 38712
rect 26007 38709 26019 38743
rect 33042 38740 33048 38752
rect 33003 38712 33048 38740
rect 25961 38703 26019 38709
rect 33042 38700 33048 38712
rect 33100 38700 33106 38752
rect 33502 38740 33508 38752
rect 33463 38712 33508 38740
rect 33502 38700 33508 38712
rect 33560 38700 33566 38752
rect 34146 38700 34152 38752
rect 34204 38740 34210 38752
rect 34241 38743 34299 38749
rect 34241 38740 34253 38743
rect 34204 38712 34253 38740
rect 34204 38700 34210 38712
rect 34241 38709 34253 38712
rect 34287 38709 34299 38743
rect 34241 38703 34299 38709
rect 36354 38700 36360 38752
rect 36412 38740 36418 38752
rect 36541 38743 36599 38749
rect 36541 38740 36553 38743
rect 36412 38712 36553 38740
rect 36412 38700 36418 38712
rect 36541 38709 36553 38712
rect 36587 38709 36599 38743
rect 36541 38703 36599 38709
rect 37277 38743 37335 38749
rect 37277 38709 37289 38743
rect 37323 38740 37335 38743
rect 37458 38740 37464 38752
rect 37323 38712 37464 38740
rect 37323 38709 37335 38712
rect 37277 38703 37335 38709
rect 37458 38700 37464 38712
rect 37516 38700 37522 38752
rect 39025 38743 39083 38749
rect 39025 38709 39037 38743
rect 39071 38740 39083 38743
rect 39850 38740 39856 38752
rect 39071 38712 39856 38740
rect 39071 38709 39083 38712
rect 39025 38703 39083 38709
rect 39850 38700 39856 38712
rect 39908 38700 39914 38752
rect 44174 38740 44180 38752
rect 44135 38712 44180 38740
rect 44174 38700 44180 38712
rect 44232 38700 44238 38752
rect 1104 38650 44896 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 44896 38650
rect 1104 38576 44896 38598
rect 19334 38536 19340 38548
rect 19295 38508 19340 38536
rect 19334 38496 19340 38508
rect 19392 38496 19398 38548
rect 22186 38536 22192 38548
rect 22147 38508 22192 38536
rect 22186 38496 22192 38508
rect 22244 38496 22250 38548
rect 29730 38496 29736 38548
rect 29788 38536 29794 38548
rect 29917 38539 29975 38545
rect 29917 38536 29929 38539
rect 29788 38508 29929 38536
rect 29788 38496 29794 38508
rect 29917 38505 29929 38508
rect 29963 38505 29975 38539
rect 29917 38499 29975 38505
rect 34974 38468 34980 38480
rect 34935 38440 34980 38468
rect 34974 38428 34980 38440
rect 35032 38428 35038 38480
rect 19705 38403 19763 38409
rect 19705 38369 19717 38403
rect 19751 38400 19763 38403
rect 20254 38400 20260 38412
rect 19751 38372 20260 38400
rect 19751 38369 19763 38372
rect 19705 38363 19763 38369
rect 20254 38360 20260 38372
rect 20312 38360 20318 38412
rect 21634 38400 21640 38412
rect 21595 38372 21640 38400
rect 21634 38360 21640 38372
rect 21692 38360 21698 38412
rect 25314 38360 25320 38412
rect 25372 38400 25378 38412
rect 25372 38372 26556 38400
rect 25372 38360 25378 38372
rect 15838 38292 15844 38344
rect 15896 38332 15902 38344
rect 16301 38335 16359 38341
rect 16301 38332 16313 38335
rect 15896 38304 16313 38332
rect 15896 38292 15902 38304
rect 16301 38301 16313 38304
rect 16347 38332 16359 38335
rect 16390 38332 16396 38344
rect 16347 38304 16396 38332
rect 16347 38301 16359 38304
rect 16301 38295 16359 38301
rect 16390 38292 16396 38304
rect 16448 38292 16454 38344
rect 16568 38335 16626 38341
rect 16568 38301 16580 38335
rect 16614 38332 16626 38335
rect 16850 38332 16856 38344
rect 16614 38304 16856 38332
rect 16614 38301 16626 38304
rect 16568 38295 16626 38301
rect 16850 38292 16856 38304
rect 16908 38292 16914 38344
rect 19521 38335 19579 38341
rect 19521 38301 19533 38335
rect 19567 38301 19579 38335
rect 19521 38295 19579 38301
rect 19797 38335 19855 38341
rect 19797 38301 19809 38335
rect 19843 38332 19855 38335
rect 20070 38332 20076 38344
rect 19843 38304 20076 38332
rect 19843 38301 19855 38304
rect 19797 38295 19855 38301
rect 19426 38224 19432 38276
rect 19484 38264 19490 38276
rect 19536 38264 19564 38295
rect 20070 38292 20076 38304
rect 20128 38292 20134 38344
rect 21542 38292 21548 38344
rect 21600 38332 21606 38344
rect 22097 38335 22155 38341
rect 22097 38332 22109 38335
rect 21600 38304 22109 38332
rect 21600 38292 21606 38304
rect 22097 38301 22109 38304
rect 22143 38301 22155 38335
rect 22097 38295 22155 38301
rect 22281 38335 22339 38341
rect 22281 38301 22293 38335
rect 22327 38301 22339 38335
rect 22281 38295 22339 38301
rect 22833 38335 22891 38341
rect 22833 38301 22845 38335
rect 22879 38332 22891 38335
rect 23014 38332 23020 38344
rect 22879 38304 23020 38332
rect 22879 38301 22891 38304
rect 22833 38295 22891 38301
rect 20346 38264 20352 38276
rect 19484 38236 20352 38264
rect 19484 38224 19490 38236
rect 20346 38224 20352 38236
rect 20404 38224 20410 38276
rect 21266 38224 21272 38276
rect 21324 38264 21330 38276
rect 21370 38267 21428 38273
rect 21370 38264 21382 38267
rect 21324 38236 21382 38264
rect 21324 38224 21330 38236
rect 21370 38233 21382 38236
rect 21416 38233 21428 38267
rect 22296 38264 22324 38295
rect 23014 38292 23020 38304
rect 23072 38292 23078 38344
rect 25593 38335 25651 38341
rect 25593 38301 25605 38335
rect 25639 38301 25651 38335
rect 25866 38332 25872 38344
rect 25827 38304 25872 38332
rect 25593 38295 25651 38301
rect 24762 38264 24768 38276
rect 22296 38236 24768 38264
rect 21370 38227 21428 38233
rect 24762 38224 24768 38236
rect 24820 38224 24826 38276
rect 25608 38264 25636 38295
rect 25866 38292 25872 38304
rect 25924 38292 25930 38344
rect 26528 38341 26556 38372
rect 33226 38360 33232 38412
rect 33284 38400 33290 38412
rect 33321 38403 33379 38409
rect 33321 38400 33333 38403
rect 33284 38372 33333 38400
rect 33284 38360 33290 38372
rect 33321 38369 33333 38372
rect 33367 38369 33379 38403
rect 36078 38400 36084 38412
rect 36039 38372 36084 38400
rect 33321 38363 33379 38369
rect 36078 38360 36084 38372
rect 36136 38360 36142 38412
rect 37642 38360 37648 38412
rect 37700 38400 37706 38412
rect 38473 38403 38531 38409
rect 38473 38400 38485 38403
rect 37700 38372 38485 38400
rect 37700 38360 37706 38372
rect 38473 38369 38485 38372
rect 38519 38369 38531 38403
rect 38473 38363 38531 38369
rect 38565 38403 38623 38409
rect 38565 38369 38577 38403
rect 38611 38400 38623 38403
rect 38654 38400 38660 38412
rect 38611 38372 38660 38400
rect 38611 38369 38623 38372
rect 38565 38363 38623 38369
rect 38654 38360 38660 38372
rect 38712 38400 38718 38412
rect 38838 38400 38844 38412
rect 38712 38372 38844 38400
rect 38712 38360 38718 38372
rect 38838 38360 38844 38372
rect 38896 38360 38902 38412
rect 39942 38360 39948 38412
rect 40000 38400 40006 38412
rect 40497 38403 40555 38409
rect 40497 38400 40509 38403
rect 40000 38372 40509 38400
rect 40000 38360 40006 38372
rect 40497 38369 40509 38372
rect 40543 38369 40555 38403
rect 42702 38400 42708 38412
rect 42663 38372 42708 38400
rect 40497 38363 40555 38369
rect 42702 38360 42708 38372
rect 42760 38360 42766 38412
rect 44174 38400 44180 38412
rect 44135 38372 44180 38400
rect 44174 38360 44180 38372
rect 44232 38360 44238 38412
rect 26513 38335 26571 38341
rect 26513 38301 26525 38335
rect 26559 38301 26571 38335
rect 30098 38332 30104 38344
rect 30059 38304 30104 38332
rect 26513 38295 26571 38301
rect 30098 38292 30104 38304
rect 30156 38292 30162 38344
rect 33597 38335 33655 38341
rect 33597 38301 33609 38335
rect 33643 38332 33655 38335
rect 34698 38332 34704 38344
rect 33643 38304 34704 38332
rect 33643 38301 33655 38304
rect 33597 38295 33655 38301
rect 34698 38292 34704 38304
rect 34756 38292 34762 38344
rect 34790 38292 34796 38344
rect 34848 38332 34854 38344
rect 36354 38341 36360 38344
rect 34977 38335 35035 38341
rect 34977 38332 34989 38335
rect 34848 38304 34989 38332
rect 34848 38292 34854 38304
rect 34977 38301 34989 38304
rect 35023 38301 35035 38335
rect 36348 38332 36360 38341
rect 36315 38304 36360 38332
rect 34977 38295 35035 38301
rect 36348 38295 36360 38304
rect 36354 38292 36360 38295
rect 36412 38292 36418 38344
rect 38197 38335 38255 38341
rect 38197 38332 38209 38335
rect 37476 38304 38209 38332
rect 26234 38264 26240 38276
rect 25608 38236 26240 38264
rect 26234 38224 26240 38236
rect 26292 38224 26298 38276
rect 27154 38264 27160 38276
rect 26436 38236 27160 38264
rect 17310 38156 17316 38208
rect 17368 38196 17374 38208
rect 17681 38199 17739 38205
rect 17681 38196 17693 38199
rect 17368 38168 17693 38196
rect 17368 38156 17374 38168
rect 17681 38165 17693 38168
rect 17727 38165 17739 38199
rect 20254 38196 20260 38208
rect 20215 38168 20260 38196
rect 17681 38159 17739 38165
rect 20254 38156 20260 38168
rect 20312 38156 20318 38208
rect 22922 38156 22928 38208
rect 22980 38196 22986 38208
rect 23017 38199 23075 38205
rect 23017 38196 23029 38199
rect 22980 38168 23029 38196
rect 22980 38156 22986 38168
rect 23017 38165 23029 38168
rect 23063 38165 23075 38199
rect 23017 38159 23075 38165
rect 24946 38156 24952 38208
rect 25004 38196 25010 38208
rect 25409 38199 25467 38205
rect 25409 38196 25421 38199
rect 25004 38168 25421 38196
rect 25004 38156 25010 38168
rect 25409 38165 25421 38168
rect 25455 38196 25467 38199
rect 25498 38196 25504 38208
rect 25455 38168 25504 38196
rect 25455 38165 25467 38168
rect 25409 38159 25467 38165
rect 25498 38156 25504 38168
rect 25556 38156 25562 38208
rect 25777 38199 25835 38205
rect 25777 38165 25789 38199
rect 25823 38196 25835 38199
rect 26142 38196 26148 38208
rect 25823 38168 26148 38196
rect 25823 38165 25835 38168
rect 25777 38159 25835 38165
rect 26142 38156 26148 38168
rect 26200 38196 26206 38208
rect 26436 38196 26464 38236
rect 27154 38224 27160 38236
rect 27212 38224 27218 38276
rect 26200 38168 26464 38196
rect 26605 38199 26663 38205
rect 26200 38156 26206 38168
rect 26605 38165 26617 38199
rect 26651 38196 26663 38199
rect 27982 38196 27988 38208
rect 26651 38168 27988 38196
rect 26651 38165 26663 38168
rect 26605 38159 26663 38165
rect 27982 38156 27988 38168
rect 28040 38196 28046 38208
rect 28810 38196 28816 38208
rect 28040 38168 28816 38196
rect 28040 38156 28046 38168
rect 28810 38156 28816 38168
rect 28868 38156 28874 38208
rect 34146 38156 34152 38208
rect 34204 38196 34210 38208
rect 34793 38199 34851 38205
rect 34793 38196 34805 38199
rect 34204 38168 34805 38196
rect 34204 38156 34210 38168
rect 34793 38165 34805 38168
rect 34839 38165 34851 38199
rect 34793 38159 34851 38165
rect 37366 38156 37372 38208
rect 37424 38196 37430 38208
rect 37476 38205 37504 38304
rect 38197 38301 38209 38304
rect 38243 38301 38255 38335
rect 39850 38332 39856 38344
rect 39811 38304 39856 38332
rect 38197 38295 38255 38301
rect 39850 38292 39856 38304
rect 39908 38292 39914 38344
rect 40034 38332 40040 38344
rect 39995 38304 40040 38332
rect 40034 38292 40040 38304
rect 40092 38292 40098 38344
rect 38682 38267 38740 38273
rect 38682 38233 38694 38267
rect 38728 38264 38740 38267
rect 39666 38264 39672 38276
rect 38728 38236 39672 38264
rect 38728 38233 38740 38236
rect 38682 38227 38740 38233
rect 39666 38224 39672 38236
rect 39724 38224 39730 38276
rect 40764 38267 40822 38273
rect 40764 38233 40776 38267
rect 40810 38264 40822 38267
rect 41138 38264 41144 38276
rect 40810 38236 41144 38264
rect 40810 38233 40822 38236
rect 40764 38227 40822 38233
rect 41138 38224 41144 38236
rect 41196 38224 41202 38276
rect 43622 38224 43628 38276
rect 43680 38264 43686 38276
rect 43993 38267 44051 38273
rect 43993 38264 44005 38267
rect 43680 38236 44005 38264
rect 43680 38224 43686 38236
rect 43993 38233 44005 38236
rect 44039 38233 44051 38267
rect 43993 38227 44051 38233
rect 37461 38199 37519 38205
rect 37461 38196 37473 38199
rect 37424 38168 37473 38196
rect 37424 38156 37430 38168
rect 37461 38165 37473 38168
rect 37507 38165 37519 38199
rect 38838 38196 38844 38208
rect 38799 38168 38844 38196
rect 37461 38159 37519 38165
rect 38838 38156 38844 38168
rect 38896 38156 38902 38208
rect 39574 38156 39580 38208
rect 39632 38196 39638 38208
rect 39945 38199 40003 38205
rect 39945 38196 39957 38199
rect 39632 38168 39957 38196
rect 39632 38156 39638 38168
rect 39945 38165 39957 38168
rect 39991 38165 40003 38199
rect 39945 38159 40003 38165
rect 41598 38156 41604 38208
rect 41656 38196 41662 38208
rect 41877 38199 41935 38205
rect 41877 38196 41889 38199
rect 41656 38168 41889 38196
rect 41656 38156 41662 38168
rect 41877 38165 41889 38168
rect 41923 38196 41935 38199
rect 42426 38196 42432 38208
rect 41923 38168 42432 38196
rect 41923 38165 41935 38168
rect 41877 38159 41935 38165
rect 42426 38156 42432 38168
rect 42484 38156 42490 38208
rect 1104 38106 44896 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 44896 38106
rect 1104 38032 44896 38054
rect 16942 37952 16948 38004
rect 17000 37992 17006 38004
rect 17313 37995 17371 38001
rect 17313 37992 17325 37995
rect 17000 37964 17325 37992
rect 17000 37952 17006 37964
rect 17313 37961 17325 37964
rect 17359 37961 17371 37995
rect 18414 37992 18420 38004
rect 18375 37964 18420 37992
rect 17313 37955 17371 37961
rect 18414 37952 18420 37964
rect 18472 37992 18478 38004
rect 19334 37992 19340 38004
rect 18472 37964 19340 37992
rect 18472 37952 18478 37964
rect 19334 37952 19340 37964
rect 19392 37952 19398 38004
rect 20438 37952 20444 38004
rect 20496 37992 20502 38004
rect 20533 37995 20591 38001
rect 20533 37992 20545 37995
rect 20496 37964 20545 37992
rect 20496 37952 20502 37964
rect 20533 37961 20545 37964
rect 20579 37961 20591 37995
rect 21266 37992 21272 38004
rect 21227 37964 21272 37992
rect 20533 37955 20591 37961
rect 21266 37952 21272 37964
rect 21324 37952 21330 38004
rect 33226 37952 33232 38004
rect 33284 37992 33290 38004
rect 33413 37995 33471 38001
rect 33413 37992 33425 37995
rect 33284 37964 33425 37992
rect 33284 37952 33290 37964
rect 33413 37961 33425 37964
rect 33459 37961 33471 37995
rect 33413 37955 33471 37961
rect 34054 37952 34060 38004
rect 34112 37992 34118 38004
rect 34241 37995 34299 38001
rect 34241 37992 34253 37995
rect 34112 37964 34253 37992
rect 34112 37952 34118 37964
rect 34241 37961 34253 37964
rect 34287 37961 34299 37995
rect 37274 37992 37280 38004
rect 37235 37964 37280 37992
rect 34241 37955 34299 37961
rect 37274 37952 37280 37964
rect 37332 37952 37338 38004
rect 38473 37995 38531 38001
rect 37384 37964 38424 37992
rect 4798 37884 4804 37936
rect 4856 37924 4862 37936
rect 37384 37924 37412 37964
rect 4856 37896 37412 37924
rect 37445 37927 37503 37933
rect 4856 37884 4862 37896
rect 37445 37893 37457 37927
rect 37491 37924 37503 37927
rect 37645 37927 37703 37933
rect 37491 37893 37504 37924
rect 37445 37887 37504 37893
rect 37645 37893 37657 37927
rect 37691 37893 37703 37927
rect 37645 37887 37703 37893
rect 17037 37859 17095 37865
rect 17037 37825 17049 37859
rect 17083 37856 17095 37859
rect 17586 37856 17592 37868
rect 17083 37828 17592 37856
rect 17083 37825 17095 37828
rect 17037 37819 17095 37825
rect 17586 37816 17592 37828
rect 17644 37816 17650 37868
rect 18598 37856 18604 37868
rect 18559 37828 18604 37856
rect 18598 37816 18604 37828
rect 18656 37816 18662 37868
rect 18785 37859 18843 37865
rect 18785 37825 18797 37859
rect 18831 37825 18843 37859
rect 18785 37819 18843 37825
rect 17310 37788 17316 37800
rect 17271 37760 17316 37788
rect 17310 37748 17316 37760
rect 17368 37748 17374 37800
rect 18800 37720 18828 37819
rect 18874 37816 18880 37868
rect 18932 37856 18938 37868
rect 18932 37828 19472 37856
rect 18932 37816 18938 37828
rect 19334 37788 19340 37800
rect 19295 37760 19340 37788
rect 19334 37748 19340 37760
rect 19392 37748 19398 37800
rect 19444 37788 19472 37828
rect 19518 37816 19524 37868
rect 19576 37856 19582 37868
rect 20165 37859 20223 37865
rect 19576 37828 19621 37856
rect 19576 37816 19582 37828
rect 20165 37825 20177 37859
rect 20211 37825 20223 37859
rect 20165 37819 20223 37825
rect 20993 37859 21051 37865
rect 20993 37825 21005 37859
rect 21039 37825 21051 37859
rect 20993 37819 21051 37825
rect 20180 37788 20208 37819
rect 19444 37760 20208 37788
rect 20254 37748 20260 37800
rect 20312 37788 20318 37800
rect 20312 37760 20357 37788
rect 20312 37748 20318 37760
rect 19426 37720 19432 37732
rect 18800 37692 19432 37720
rect 19426 37680 19432 37692
rect 19484 37680 19490 37732
rect 19705 37723 19763 37729
rect 19705 37689 19717 37723
rect 19751 37720 19763 37723
rect 21008 37720 21036 37819
rect 21634 37816 21640 37868
rect 21692 37856 21698 37868
rect 23198 37865 23204 37868
rect 22925 37859 22983 37865
rect 22925 37856 22937 37859
rect 21692 37828 22937 37856
rect 21692 37816 21698 37828
rect 22925 37825 22937 37828
rect 22971 37825 22983 37859
rect 23192 37856 23204 37865
rect 23159 37828 23204 37856
rect 22925 37819 22983 37825
rect 23192 37819 23204 37828
rect 23198 37816 23204 37819
rect 23256 37816 23262 37868
rect 25041 37859 25099 37865
rect 25041 37825 25053 37859
rect 25087 37856 25099 37859
rect 25498 37856 25504 37868
rect 25087 37828 25504 37856
rect 25087 37825 25099 37828
rect 25041 37819 25099 37825
rect 25498 37816 25504 37828
rect 25556 37816 25562 37868
rect 25593 37859 25651 37865
rect 25593 37825 25605 37859
rect 25639 37856 25651 37859
rect 26234 37856 26240 37868
rect 25639 37828 26240 37856
rect 25639 37825 25651 37828
rect 25593 37819 25651 37825
rect 26234 37816 26240 37828
rect 26292 37816 26298 37868
rect 27341 37859 27399 37865
rect 27341 37825 27353 37859
rect 27387 37856 27399 37859
rect 27798 37856 27804 37868
rect 27387 37828 27804 37856
rect 27387 37825 27399 37828
rect 27341 37819 27399 37825
rect 27798 37816 27804 37828
rect 27856 37856 27862 37868
rect 28077 37859 28135 37865
rect 28077 37856 28089 37859
rect 27856 37828 28089 37856
rect 27856 37816 27862 37828
rect 28077 37825 28089 37828
rect 28123 37825 28135 37859
rect 28077 37819 28135 37825
rect 31481 37859 31539 37865
rect 31481 37825 31493 37859
rect 31527 37856 31539 37859
rect 32030 37856 32036 37868
rect 31527 37828 32036 37856
rect 31527 37825 31539 37828
rect 31481 37819 31539 37825
rect 32030 37816 32036 37828
rect 32088 37816 32094 37868
rect 32125 37859 32183 37865
rect 32125 37825 32137 37859
rect 32171 37825 32183 37859
rect 32125 37819 32183 37825
rect 21269 37791 21327 37797
rect 21269 37757 21281 37791
rect 21315 37788 21327 37791
rect 21450 37788 21456 37800
rect 21315 37760 21456 37788
rect 21315 37757 21327 37760
rect 21269 37751 21327 37757
rect 21450 37748 21456 37760
rect 21508 37748 21514 37800
rect 24394 37788 24400 37800
rect 24307 37760 24400 37788
rect 24320 37729 24348 37760
rect 24394 37748 24400 37760
rect 24452 37788 24458 37800
rect 24670 37788 24676 37800
rect 24452 37760 24676 37788
rect 24452 37748 24458 37760
rect 24670 37748 24676 37760
rect 24728 37788 24734 37800
rect 24765 37791 24823 37797
rect 24765 37788 24777 37791
rect 24728 37760 24777 37788
rect 24728 37748 24734 37760
rect 24765 37757 24777 37760
rect 24811 37757 24823 37791
rect 25869 37791 25927 37797
rect 25869 37788 25881 37791
rect 24765 37751 24823 37757
rect 25056 37760 25881 37788
rect 19751 37692 21036 37720
rect 24305 37723 24363 37729
rect 19751 37689 19763 37692
rect 19705 37683 19763 37689
rect 24305 37689 24317 37723
rect 24351 37689 24363 37723
rect 24305 37683 24363 37689
rect 25056 37664 25084 37760
rect 25869 37757 25881 37760
rect 25915 37757 25927 37791
rect 25869 37751 25927 37757
rect 27617 37791 27675 37797
rect 27617 37757 27629 37791
rect 27663 37788 27675 37791
rect 27706 37788 27712 37800
rect 27663 37760 27712 37788
rect 27663 37757 27675 37760
rect 27617 37751 27675 37757
rect 27706 37748 27712 37760
rect 27764 37788 27770 37800
rect 28902 37788 28908 37800
rect 27764 37760 28908 37788
rect 27764 37748 27770 37760
rect 28902 37748 28908 37760
rect 28960 37748 28966 37800
rect 32140 37788 32168 37819
rect 32214 37816 32220 37868
rect 32272 37856 32278 37868
rect 32398 37856 32404 37868
rect 32272 37828 32317 37856
rect 32359 37828 32404 37856
rect 32272 37816 32278 37828
rect 32398 37816 32404 37828
rect 32456 37816 32462 37868
rect 33410 37816 33416 37868
rect 33468 37856 33474 37868
rect 33505 37859 33563 37865
rect 33505 37856 33517 37859
rect 33468 37828 33517 37856
rect 33468 37816 33474 37828
rect 33505 37825 33517 37828
rect 33551 37825 33563 37859
rect 33505 37819 33563 37825
rect 33594 37816 33600 37868
rect 33652 37856 33658 37868
rect 33781 37859 33839 37865
rect 33652 37828 33697 37856
rect 33652 37816 33658 37828
rect 33781 37825 33793 37859
rect 33827 37856 33839 37859
rect 34054 37856 34060 37868
rect 33827 37828 34060 37856
rect 33827 37825 33839 37828
rect 33781 37819 33839 37825
rect 34054 37816 34060 37828
rect 34112 37816 34118 37868
rect 34974 37816 34980 37868
rect 35032 37856 35038 37868
rect 35354 37859 35412 37865
rect 35354 37856 35366 37859
rect 35032 37828 35366 37856
rect 35032 37816 35038 37828
rect 35354 37825 35366 37828
rect 35400 37825 35412 37859
rect 35354 37819 35412 37825
rect 37274 37816 37280 37868
rect 37332 37854 37338 37868
rect 37476 37854 37504 37887
rect 37332 37826 37504 37854
rect 37332 37816 37338 37826
rect 32490 37788 32496 37800
rect 32140 37760 32496 37788
rect 32490 37748 32496 37760
rect 32548 37748 32554 37800
rect 35621 37791 35679 37797
rect 35621 37757 35633 37791
rect 35667 37788 35679 37791
rect 36078 37788 36084 37800
rect 35667 37760 36084 37788
rect 35667 37757 35679 37760
rect 35621 37751 35679 37757
rect 36078 37748 36084 37760
rect 36136 37748 36142 37800
rect 27430 37720 27436 37732
rect 27391 37692 27436 37720
rect 27430 37680 27436 37692
rect 27488 37680 27494 37732
rect 32674 37680 32680 37732
rect 32732 37720 32738 37732
rect 37660 37720 37688 37887
rect 38396 37856 38424 37964
rect 38473 37961 38485 37995
rect 38519 37992 38531 37995
rect 38654 37992 38660 38004
rect 38519 37964 38660 37992
rect 38519 37961 38531 37964
rect 38473 37955 38531 37961
rect 38654 37952 38660 37964
rect 38712 37952 38718 38004
rect 41138 37992 41144 38004
rect 41099 37964 41144 37992
rect 41138 37952 41144 37964
rect 41196 37952 41202 38004
rect 42705 37995 42763 38001
rect 42705 37992 42717 37995
rect 41248 37964 42717 37992
rect 39574 37884 39580 37936
rect 39632 37933 39638 37936
rect 39632 37924 39644 37933
rect 39632 37896 39677 37924
rect 39632 37887 39644 37896
rect 39632 37884 39638 37887
rect 39853 37859 39911 37865
rect 38396 37828 39804 37856
rect 39776 37788 39804 37828
rect 39853 37825 39865 37859
rect 39899 37856 39911 37859
rect 39942 37856 39948 37868
rect 39899 37828 39948 37856
rect 39899 37825 39911 37828
rect 39853 37819 39911 37825
rect 39942 37816 39948 37828
rect 40000 37816 40006 37868
rect 41046 37856 41052 37868
rect 41007 37828 41052 37856
rect 41046 37816 41052 37828
rect 41104 37816 41110 37868
rect 41248 37865 41276 37964
rect 42705 37961 42717 37964
rect 42751 37961 42763 37995
rect 43622 37992 43628 38004
rect 43583 37964 43628 37992
rect 42705 37955 42763 37961
rect 43622 37952 43628 37964
rect 43680 37952 43686 38004
rect 43254 37924 43260 37936
rect 41892 37896 43260 37924
rect 41892 37865 41920 37896
rect 43254 37884 43260 37896
rect 43312 37884 43318 37936
rect 41233 37859 41291 37865
rect 41233 37825 41245 37859
rect 41279 37825 41291 37859
rect 41233 37819 41291 37825
rect 41693 37859 41751 37865
rect 41693 37825 41705 37859
rect 41739 37825 41751 37859
rect 41693 37819 41751 37825
rect 41877 37859 41935 37865
rect 41877 37825 41889 37859
rect 41923 37825 41935 37859
rect 42426 37856 42432 37868
rect 42387 37828 42432 37856
rect 41877 37819 41935 37825
rect 41708 37788 41736 37819
rect 42426 37816 42432 37828
rect 42484 37816 42490 37868
rect 43533 37859 43591 37865
rect 43533 37825 43545 37859
rect 43579 37856 43591 37859
rect 43714 37856 43720 37868
rect 43579 37828 43720 37856
rect 43579 37825 43591 37828
rect 43533 37819 43591 37825
rect 43714 37816 43720 37828
rect 43772 37816 43778 37868
rect 42521 37791 42579 37797
rect 42521 37788 42533 37791
rect 39776 37760 41414 37788
rect 41708 37760 42533 37788
rect 32732 37692 33364 37720
rect 32732 37680 32738 37692
rect 2133 37655 2191 37661
rect 2133 37621 2145 37655
rect 2179 37652 2191 37655
rect 3234 37652 3240 37664
rect 2179 37624 3240 37652
rect 2179 37621 2191 37624
rect 2133 37615 2191 37621
rect 3234 37612 3240 37624
rect 3292 37612 3298 37664
rect 17126 37652 17132 37664
rect 17087 37624 17132 37652
rect 17126 37612 17132 37624
rect 17184 37612 17190 37664
rect 19518 37612 19524 37664
rect 19576 37652 19582 37664
rect 20165 37655 20223 37661
rect 20165 37652 20177 37655
rect 19576 37624 20177 37652
rect 19576 37612 19582 37624
rect 20165 37621 20177 37624
rect 20211 37621 20223 37655
rect 20165 37615 20223 37621
rect 20254 37612 20260 37664
rect 20312 37652 20318 37664
rect 21085 37655 21143 37661
rect 21085 37652 21097 37655
rect 20312 37624 21097 37652
rect 20312 37612 20318 37624
rect 21085 37621 21097 37624
rect 21131 37621 21143 37655
rect 24854 37652 24860 37664
rect 24815 37624 24860 37652
rect 21085 37615 21143 37621
rect 24854 37612 24860 37624
rect 24912 37612 24918 37664
rect 24949 37655 25007 37661
rect 24949 37621 24961 37655
rect 24995 37652 25007 37655
rect 25038 37652 25044 37664
rect 24995 37624 25044 37652
rect 24995 37621 25007 37624
rect 24949 37615 25007 37621
rect 25038 37612 25044 37624
rect 25096 37612 25102 37664
rect 26326 37612 26332 37664
rect 26384 37652 26390 37664
rect 27341 37655 27399 37661
rect 27341 37652 27353 37655
rect 26384 37624 27353 37652
rect 26384 37612 26390 37624
rect 27341 37621 27353 37624
rect 27387 37621 27399 37655
rect 27341 37615 27399 37621
rect 27522 37612 27528 37664
rect 27580 37652 27586 37664
rect 28169 37655 28227 37661
rect 28169 37652 28181 37655
rect 27580 37624 28181 37652
rect 27580 37612 27586 37624
rect 28169 37621 28181 37624
rect 28215 37621 28227 37655
rect 31294 37652 31300 37664
rect 31255 37624 31300 37652
rect 28169 37615 28227 37621
rect 31294 37612 31300 37624
rect 31352 37612 31358 37664
rect 32582 37652 32588 37664
rect 32543 37624 32588 37652
rect 32582 37612 32588 37624
rect 32640 37612 32646 37664
rect 33042 37612 33048 37664
rect 33100 37652 33106 37664
rect 33229 37655 33287 37661
rect 33229 37652 33241 37655
rect 33100 37624 33241 37652
rect 33100 37612 33106 37624
rect 33229 37621 33241 37624
rect 33275 37621 33287 37655
rect 33336 37652 33364 37692
rect 35866 37692 37688 37720
rect 41386 37720 41414 37760
rect 42444 37732 42472 37760
rect 42521 37757 42533 37760
rect 42567 37757 42579 37791
rect 42521 37751 42579 37757
rect 42702 37748 42708 37800
rect 42760 37788 42766 37800
rect 42886 37788 42892 37800
rect 42760 37760 42892 37788
rect 42760 37748 42766 37760
rect 42886 37748 42892 37760
rect 42944 37748 42950 37800
rect 41386 37692 42380 37720
rect 35866 37652 35894 37692
rect 37458 37652 37464 37664
rect 33336 37624 35894 37652
rect 37419 37624 37464 37652
rect 33229 37615 33287 37621
rect 37458 37612 37464 37624
rect 37516 37612 37522 37664
rect 41877 37655 41935 37661
rect 41877 37621 41889 37655
rect 41923 37652 41935 37655
rect 42242 37652 42248 37664
rect 41923 37624 42248 37652
rect 41923 37621 41935 37624
rect 41877 37615 41935 37621
rect 42242 37612 42248 37624
rect 42300 37612 42306 37664
rect 42352 37652 42380 37692
rect 42426 37680 42432 37732
rect 42484 37680 42490 37732
rect 43714 37652 43720 37664
rect 42352 37624 43720 37652
rect 43714 37612 43720 37624
rect 43772 37612 43778 37664
rect 1104 37562 44896 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 44896 37562
rect 1104 37488 44896 37510
rect 18509 37451 18567 37457
rect 18509 37417 18521 37451
rect 18555 37448 18567 37451
rect 18874 37448 18880 37460
rect 18555 37420 18880 37448
rect 18555 37417 18567 37420
rect 18509 37411 18567 37417
rect 18874 37408 18880 37420
rect 18932 37408 18938 37460
rect 23198 37408 23204 37460
rect 23256 37448 23262 37460
rect 23385 37451 23443 37457
rect 23385 37448 23397 37451
rect 23256 37420 23397 37448
rect 23256 37408 23262 37420
rect 23385 37417 23397 37420
rect 23431 37417 23443 37451
rect 25222 37448 25228 37460
rect 23385 37411 23443 37417
rect 23492 37420 25228 37448
rect 19518 37312 19524 37324
rect 19479 37284 19524 37312
rect 19518 37272 19524 37284
rect 19576 37272 19582 37324
rect 23492 37321 23520 37420
rect 25222 37408 25228 37420
rect 25280 37408 25286 37460
rect 25590 37408 25596 37460
rect 25648 37448 25654 37460
rect 25869 37451 25927 37457
rect 25869 37448 25881 37451
rect 25648 37420 25881 37448
rect 25648 37408 25654 37420
rect 25869 37417 25881 37420
rect 25915 37417 25927 37451
rect 25869 37411 25927 37417
rect 32030 37408 32036 37460
rect 32088 37448 32094 37460
rect 32493 37451 32551 37457
rect 32493 37448 32505 37451
rect 32088 37420 32505 37448
rect 32088 37408 32094 37420
rect 32493 37417 32505 37420
rect 32539 37417 32551 37451
rect 32674 37448 32680 37460
rect 32635 37420 32680 37448
rect 32493 37411 32551 37417
rect 32674 37408 32680 37420
rect 32732 37408 32738 37460
rect 33410 37408 33416 37460
rect 33468 37448 33474 37460
rect 33505 37451 33563 37457
rect 33505 37448 33517 37451
rect 33468 37420 33517 37448
rect 33468 37408 33474 37420
rect 33505 37417 33517 37420
rect 33551 37417 33563 37451
rect 33505 37411 33563 37417
rect 34790 37408 34796 37460
rect 34848 37448 34854 37460
rect 34885 37451 34943 37457
rect 34885 37448 34897 37451
rect 34848 37420 34897 37448
rect 34848 37408 34854 37420
rect 34885 37417 34897 37420
rect 34931 37417 34943 37451
rect 37274 37448 37280 37460
rect 37235 37420 37280 37448
rect 34885 37411 34943 37417
rect 37274 37408 37280 37420
rect 37332 37408 37338 37460
rect 41690 37448 41696 37460
rect 41651 37420 41696 37448
rect 41690 37408 41696 37420
rect 41748 37408 41754 37460
rect 42702 37448 42708 37460
rect 42444 37420 42708 37448
rect 23753 37383 23811 37389
rect 23753 37349 23765 37383
rect 23799 37380 23811 37383
rect 25038 37380 25044 37392
rect 23799 37352 25044 37380
rect 23799 37349 23811 37352
rect 23753 37343 23811 37349
rect 25038 37340 25044 37352
rect 25096 37380 25102 37392
rect 25096 37352 26004 37380
rect 25096 37340 25102 37352
rect 23477 37315 23535 37321
rect 23477 37281 23489 37315
rect 23523 37281 23535 37315
rect 23477 37275 23535 37281
rect 23569 37315 23627 37321
rect 23569 37281 23581 37315
rect 23615 37312 23627 37315
rect 24854 37312 24860 37324
rect 23615 37284 24860 37312
rect 23615 37281 23627 37284
rect 23569 37275 23627 37281
rect 24854 37272 24860 37284
rect 24912 37272 24918 37324
rect 24946 37272 24952 37324
rect 25004 37312 25010 37324
rect 25976 37321 26004 37352
rect 27430 37340 27436 37392
rect 27488 37380 27494 37392
rect 42444 37380 42472 37420
rect 42702 37408 42708 37420
rect 42760 37408 42766 37460
rect 27488 37352 28672 37380
rect 27488 37340 27494 37352
rect 25961 37315 26019 37321
rect 25004 37284 25049 37312
rect 25004 37272 25010 37284
rect 25961 37281 25973 37315
rect 26007 37281 26019 37315
rect 25961 37275 26019 37281
rect 27522 37272 27528 37324
rect 27580 37272 27586 37324
rect 27982 37312 27988 37324
rect 27632 37284 27988 37312
rect 1394 37244 1400 37256
rect 1355 37216 1400 37244
rect 1394 37204 1400 37216
rect 1452 37204 1458 37256
rect 3234 37204 3240 37256
rect 3292 37244 3298 37256
rect 3292 37216 3337 37244
rect 3292 37204 3298 37216
rect 17310 37204 17316 37256
rect 17368 37244 17374 37256
rect 17770 37244 17776 37256
rect 17368 37216 17776 37244
rect 17368 37204 17374 37216
rect 17770 37204 17776 37216
rect 17828 37244 17834 37256
rect 18325 37247 18383 37253
rect 18325 37244 18337 37247
rect 17828 37216 18337 37244
rect 17828 37204 17834 37216
rect 18325 37213 18337 37216
rect 18371 37213 18383 37247
rect 18325 37207 18383 37213
rect 18598 37204 18604 37256
rect 18656 37244 18662 37256
rect 19245 37247 19303 37253
rect 19245 37244 19257 37247
rect 18656 37216 19257 37244
rect 18656 37204 18662 37216
rect 19245 37213 19257 37216
rect 19291 37213 19303 37247
rect 19245 37207 19303 37213
rect 20162 37204 20168 37256
rect 20220 37244 20226 37256
rect 20530 37244 20536 37256
rect 20220 37216 20536 37244
rect 20220 37204 20226 37216
rect 20530 37204 20536 37216
rect 20588 37244 20594 37256
rect 20993 37247 21051 37253
rect 20993 37244 21005 37247
rect 20588 37216 21005 37244
rect 20588 37204 20594 37216
rect 20993 37213 21005 37216
rect 21039 37213 21051 37247
rect 20993 37207 21051 37213
rect 23845 37247 23903 37253
rect 23845 37213 23857 37247
rect 23891 37244 23903 37247
rect 24670 37244 24676 37256
rect 23891 37216 24676 37244
rect 23891 37213 23903 37216
rect 23845 37207 23903 37213
rect 24670 37204 24676 37216
rect 24728 37204 24734 37256
rect 24762 37204 24768 37256
rect 24820 37244 24826 37256
rect 25041 37247 25099 37253
rect 24820 37216 24865 37244
rect 24820 37204 24826 37216
rect 25041 37213 25053 37247
rect 25087 37244 25099 37247
rect 26145 37247 26203 37253
rect 26145 37244 26157 37247
rect 25087 37216 26157 37244
rect 25087 37213 25099 37216
rect 25041 37207 25099 37213
rect 26145 37213 26157 37216
rect 26191 37244 26203 37247
rect 27428 37247 27486 37253
rect 27428 37244 27440 37247
rect 26191 37216 27440 37244
rect 26191 37213 26203 37216
rect 26145 37207 26203 37213
rect 27428 37213 27440 37216
rect 27474 37244 27486 37247
rect 27540 37244 27568 37272
rect 27632 37253 27660 37284
rect 27982 37272 27988 37284
rect 28040 37272 28046 37324
rect 28644 37321 28672 37352
rect 39132 37352 42472 37380
rect 39132 37324 39160 37352
rect 28353 37315 28411 37321
rect 28353 37281 28365 37315
rect 28399 37281 28411 37315
rect 28353 37275 28411 37281
rect 28629 37315 28687 37321
rect 28629 37281 28641 37315
rect 28675 37281 28687 37315
rect 33042 37312 33048 37324
rect 33003 37284 33048 37312
rect 28629 37275 28687 37281
rect 27474 37216 27568 37244
rect 27617 37247 27675 37253
rect 27474 37213 27486 37216
rect 27428 37207 27486 37213
rect 27617 37213 27629 37247
rect 27663 37213 27675 37247
rect 27617 37207 27675 37213
rect 27800 37247 27858 37253
rect 27800 37213 27812 37247
rect 27846 37213 27858 37247
rect 27800 37207 27858 37213
rect 27893 37247 27951 37253
rect 27893 37213 27905 37247
rect 27939 37244 27951 37247
rect 28368 37244 28396 37275
rect 33042 37272 33048 37284
rect 33100 37272 33106 37324
rect 33873 37315 33931 37321
rect 33873 37312 33885 37315
rect 33152 37284 33885 37312
rect 27939 37216 28396 37244
rect 27939 37213 27951 37216
rect 27893 37207 27951 37213
rect 2682 37136 2688 37188
rect 2740 37176 2746 37188
rect 3053 37179 3111 37185
rect 3053 37176 3065 37179
rect 2740 37148 3065 37176
rect 2740 37136 2746 37148
rect 3053 37145 3065 37148
rect 3099 37145 3111 37179
rect 3053 37139 3111 37145
rect 17586 37136 17592 37188
rect 17644 37176 17650 37188
rect 18141 37179 18199 37185
rect 18141 37176 18153 37179
rect 17644 37148 18153 37176
rect 17644 37136 17650 37148
rect 18141 37145 18153 37148
rect 18187 37145 18199 37179
rect 25866 37176 25872 37188
rect 25827 37148 25872 37176
rect 18141 37139 18199 37145
rect 25866 37136 25872 37148
rect 25924 37136 25930 37188
rect 27522 37176 27528 37188
rect 27483 37148 27528 37176
rect 27522 37136 27528 37148
rect 27580 37136 27586 37188
rect 21085 37111 21143 37117
rect 21085 37077 21097 37111
rect 21131 37108 21143 37111
rect 21174 37108 21180 37120
rect 21131 37080 21180 37108
rect 21131 37077 21143 37080
rect 21085 37071 21143 37077
rect 21174 37068 21180 37080
rect 21232 37068 21238 37120
rect 25409 37111 25467 37117
rect 25409 37077 25421 37111
rect 25455 37108 25467 37111
rect 26329 37111 26387 37117
rect 26329 37108 26341 37111
rect 25455 37080 26341 37108
rect 25455 37077 25467 37080
rect 25409 37071 25467 37077
rect 26329 37077 26341 37080
rect 26375 37077 26387 37111
rect 27246 37108 27252 37120
rect 27207 37080 27252 37108
rect 26329 37071 26387 37077
rect 27246 37068 27252 37080
rect 27304 37068 27310 37120
rect 27614 37068 27620 37120
rect 27672 37108 27678 37120
rect 27815 37108 27843 37207
rect 28442 37204 28448 37256
rect 28500 37244 28506 37256
rect 28721 37247 28779 37253
rect 28721 37244 28733 37247
rect 28500 37216 28733 37244
rect 28500 37204 28506 37216
rect 28721 37213 28733 37216
rect 28767 37213 28779 37247
rect 28721 37207 28779 37213
rect 30653 37247 30711 37253
rect 30653 37213 30665 37247
rect 30699 37244 30711 37247
rect 30742 37244 30748 37256
rect 30699 37216 30748 37244
rect 30699 37213 30711 37216
rect 30653 37207 30711 37213
rect 30742 37204 30748 37216
rect 30800 37204 30806 37256
rect 30920 37247 30978 37253
rect 30920 37213 30932 37247
rect 30966 37244 30978 37247
rect 31294 37244 31300 37256
rect 30966 37216 31300 37244
rect 30966 37213 30978 37216
rect 30920 37207 30978 37213
rect 31294 37204 31300 37216
rect 31352 37204 31358 37256
rect 33152 37244 33180 37284
rect 33873 37281 33885 37284
rect 33919 37281 33931 37315
rect 33873 37275 33931 37281
rect 34977 37315 35035 37321
rect 34977 37281 34989 37315
rect 35023 37312 35035 37315
rect 35342 37312 35348 37324
rect 35023 37284 35348 37312
rect 35023 37281 35035 37284
rect 34977 37275 35035 37281
rect 35342 37272 35348 37284
rect 35400 37312 35406 37324
rect 39114 37312 39120 37324
rect 35400 37284 39120 37312
rect 35400 37272 35406 37284
rect 39114 37272 39120 37284
rect 39172 37272 39178 37324
rect 41598 37312 41604 37324
rect 41559 37284 41604 37312
rect 41598 37272 41604 37284
rect 41656 37272 41662 37324
rect 32784 37216 33180 37244
rect 33689 37247 33747 37253
rect 32582 37136 32588 37188
rect 32640 37176 32646 37188
rect 32677 37179 32735 37185
rect 32677 37176 32689 37179
rect 32640 37148 32689 37176
rect 32640 37136 32646 37148
rect 32677 37145 32689 37148
rect 32723 37145 32735 37179
rect 32677 37139 32735 37145
rect 28718 37108 28724 37120
rect 27672 37080 28724 37108
rect 27672 37068 27678 37080
rect 28718 37068 28724 37080
rect 28776 37068 28782 37120
rect 32033 37111 32091 37117
rect 32033 37077 32045 37111
rect 32079 37108 32091 37111
rect 32398 37108 32404 37120
rect 32079 37080 32404 37108
rect 32079 37077 32091 37080
rect 32033 37071 32091 37077
rect 32398 37068 32404 37080
rect 32456 37108 32462 37120
rect 32784 37108 32812 37216
rect 33689 37213 33701 37247
rect 33735 37213 33747 37247
rect 33689 37207 33747 37213
rect 32950 37136 32956 37188
rect 33008 37176 33014 37188
rect 33704 37176 33732 37207
rect 34146 37204 34152 37256
rect 34204 37244 34210 37256
rect 34701 37247 34759 37253
rect 34701 37244 34713 37247
rect 34204 37216 34713 37244
rect 34204 37204 34210 37216
rect 34701 37213 34713 37216
rect 34747 37213 34759 37247
rect 34701 37207 34759 37213
rect 34790 37204 34796 37256
rect 34848 37244 34854 37256
rect 37277 37247 37335 37253
rect 34848 37216 34893 37244
rect 34848 37204 34854 37216
rect 37277 37213 37289 37247
rect 37323 37244 37335 37247
rect 37366 37244 37372 37256
rect 37323 37216 37372 37244
rect 37323 37213 37335 37216
rect 37277 37207 37335 37213
rect 37366 37204 37372 37216
rect 37424 37204 37430 37256
rect 39298 37244 39304 37256
rect 39259 37216 39304 37244
rect 39298 37204 39304 37216
rect 39356 37204 39362 37256
rect 41414 37204 41420 37256
rect 41472 37244 41478 37256
rect 42429 37247 42487 37253
rect 42429 37244 42441 37247
rect 41472 37216 41517 37244
rect 41800 37216 42441 37244
rect 41472 37204 41478 37216
rect 33008 37148 33732 37176
rect 37001 37179 37059 37185
rect 33008 37136 33014 37148
rect 37001 37145 37013 37179
rect 37047 37145 37059 37179
rect 37001 37139 37059 37145
rect 37185 37179 37243 37185
rect 37185 37145 37197 37179
rect 37231 37176 37243 37179
rect 37642 37176 37648 37188
rect 37231 37148 37648 37176
rect 37231 37145 37243 37148
rect 37185 37139 37243 37145
rect 32456 37080 32812 37108
rect 37016 37108 37044 37139
rect 37642 37136 37648 37148
rect 37700 37136 37706 37188
rect 39942 37136 39948 37188
rect 40000 37176 40006 37188
rect 41800 37176 41828 37216
rect 42429 37213 42441 37216
rect 42475 37213 42487 37247
rect 42429 37207 42487 37213
rect 40000 37148 41828 37176
rect 40000 37136 40006 37148
rect 41874 37136 41880 37188
rect 41932 37176 41938 37188
rect 41932 37148 41977 37176
rect 41932 37136 41938 37148
rect 42242 37136 42248 37188
rect 42300 37176 42306 37188
rect 42674 37179 42732 37185
rect 42674 37176 42686 37179
rect 42300 37148 42686 37176
rect 42300 37136 42306 37148
rect 42674 37145 42686 37148
rect 42720 37145 42732 37179
rect 42674 37139 42732 37145
rect 37734 37108 37740 37120
rect 37016 37080 37740 37108
rect 32456 37068 32462 37080
rect 37734 37068 37740 37080
rect 37792 37068 37798 37120
rect 38930 37068 38936 37120
rect 38988 37108 38994 37120
rect 39117 37111 39175 37117
rect 39117 37108 39129 37111
rect 38988 37080 39129 37108
rect 38988 37068 38994 37080
rect 39117 37077 39129 37080
rect 39163 37077 39175 37111
rect 39117 37071 39175 37077
rect 40218 37068 40224 37120
rect 40276 37108 40282 37120
rect 41233 37111 41291 37117
rect 41233 37108 41245 37111
rect 40276 37080 41245 37108
rect 40276 37068 40282 37080
rect 41233 37077 41245 37080
rect 41279 37077 41291 37111
rect 43806 37108 43812 37120
rect 43767 37080 43812 37108
rect 41233 37071 41291 37077
rect 43806 37068 43812 37080
rect 43864 37068 43870 37120
rect 1104 37018 44896 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 44896 37018
rect 1104 36944 44896 36966
rect 2682 36904 2688 36916
rect 2643 36876 2688 36904
rect 2682 36864 2688 36876
rect 2740 36864 2746 36916
rect 18693 36907 18751 36913
rect 18693 36873 18705 36907
rect 18739 36904 18751 36907
rect 20254 36904 20260 36916
rect 18739 36876 20260 36904
rect 18739 36873 18751 36876
rect 18693 36867 18751 36873
rect 20254 36864 20260 36876
rect 20312 36864 20318 36916
rect 20346 36864 20352 36916
rect 20404 36904 20410 36916
rect 24302 36904 24308 36916
rect 20404 36876 22324 36904
rect 24263 36876 24308 36904
rect 20404 36864 20410 36876
rect 17589 36839 17647 36845
rect 17589 36836 17601 36839
rect 16868 36808 17601 36836
rect 2777 36771 2835 36777
rect 2777 36737 2789 36771
rect 2823 36768 2835 36771
rect 7926 36768 7932 36780
rect 2823 36740 7932 36768
rect 2823 36737 2835 36740
rect 2777 36731 2835 36737
rect 7926 36728 7932 36740
rect 7984 36728 7990 36780
rect 16868 36777 16896 36808
rect 17589 36805 17601 36808
rect 17635 36805 17647 36839
rect 17589 36799 17647 36805
rect 18601 36839 18659 36845
rect 18601 36805 18613 36839
rect 18647 36836 18659 36839
rect 18874 36836 18880 36848
rect 18647 36808 18880 36836
rect 18647 36805 18659 36808
rect 18601 36799 18659 36805
rect 18874 36796 18880 36808
rect 18932 36796 18938 36848
rect 18969 36839 19027 36845
rect 18969 36805 18981 36839
rect 19015 36836 19027 36839
rect 19334 36836 19340 36848
rect 19015 36808 19340 36836
rect 19015 36805 19027 36808
rect 18969 36799 19027 36805
rect 19334 36796 19340 36808
rect 19392 36836 19398 36848
rect 21174 36836 21180 36848
rect 19392 36808 21180 36836
rect 19392 36796 19398 36808
rect 21174 36796 21180 36808
rect 21232 36796 21238 36848
rect 22002 36796 22008 36848
rect 22060 36836 22066 36848
rect 22296 36836 22324 36876
rect 24302 36864 24308 36876
rect 24360 36864 24366 36916
rect 25409 36907 25467 36913
rect 25409 36873 25421 36907
rect 25455 36873 25467 36907
rect 25409 36867 25467 36873
rect 23750 36836 23756 36848
rect 22060 36808 22232 36836
rect 22060 36796 22066 36808
rect 16853 36771 16911 36777
rect 16853 36737 16865 36771
rect 16899 36737 16911 36771
rect 16853 36731 16911 36737
rect 17129 36771 17187 36777
rect 17129 36737 17141 36771
rect 17175 36737 17187 36771
rect 17129 36731 17187 36737
rect 17865 36771 17923 36777
rect 17865 36737 17877 36771
rect 17911 36768 17923 36771
rect 18414 36768 18420 36780
rect 17911 36740 18420 36768
rect 17911 36737 17923 36740
rect 17865 36731 17923 36737
rect 16761 36703 16819 36709
rect 16761 36669 16773 36703
rect 16807 36700 16819 36703
rect 17144 36700 17172 36731
rect 18414 36728 18420 36740
rect 18472 36728 18478 36780
rect 19613 36771 19671 36777
rect 19613 36737 19625 36771
rect 19659 36768 19671 36771
rect 20254 36768 20260 36780
rect 19659 36740 20260 36768
rect 19659 36737 19671 36740
rect 19613 36731 19671 36737
rect 20254 36728 20260 36740
rect 20312 36728 20318 36780
rect 20438 36768 20444 36780
rect 20399 36740 20444 36768
rect 20438 36728 20444 36740
rect 20496 36728 20502 36780
rect 20622 36768 20628 36780
rect 20583 36740 20628 36768
rect 20622 36728 20628 36740
rect 20680 36728 20686 36780
rect 20714 36728 20720 36780
rect 20772 36768 20778 36780
rect 20993 36771 21051 36777
rect 20772 36740 20817 36768
rect 20772 36728 20778 36740
rect 20993 36737 21005 36771
rect 21039 36737 21051 36771
rect 20993 36731 21051 36737
rect 17586 36700 17592 36712
rect 16807 36672 16896 36700
rect 17144 36672 17592 36700
rect 16807 36669 16819 36672
rect 16761 36663 16819 36669
rect 16868 36644 16896 36672
rect 17586 36660 17592 36672
rect 17644 36660 17650 36712
rect 20806 36660 20812 36712
rect 20864 36700 20870 36712
rect 20901 36703 20959 36709
rect 20901 36700 20913 36703
rect 20864 36672 20913 36700
rect 20864 36660 20870 36672
rect 20901 36669 20913 36672
rect 20947 36669 20959 36703
rect 21008 36700 21036 36731
rect 21726 36728 21732 36780
rect 21784 36768 21790 36780
rect 22204 36777 22232 36808
rect 22296 36808 23756 36836
rect 22296 36777 22324 36808
rect 23750 36796 23756 36808
rect 23808 36796 23814 36848
rect 25424 36836 25452 36867
rect 30742 36864 30748 36916
rect 30800 36904 30806 36916
rect 30926 36904 30932 36916
rect 30800 36876 30932 36904
rect 30800 36864 30806 36876
rect 30926 36864 30932 36876
rect 30984 36904 30990 36916
rect 33229 36907 33287 36913
rect 33229 36904 33241 36907
rect 30984 36876 33241 36904
rect 30984 36864 30990 36876
rect 25424 36808 28672 36836
rect 22097 36771 22155 36777
rect 22097 36768 22109 36771
rect 21784 36740 22109 36768
rect 21784 36728 21790 36740
rect 22097 36737 22109 36740
rect 22143 36737 22155 36771
rect 22097 36731 22155 36737
rect 22189 36771 22247 36777
rect 22189 36737 22201 36771
rect 22235 36737 22247 36771
rect 22189 36731 22247 36737
rect 22281 36771 22339 36777
rect 22281 36737 22293 36771
rect 22327 36737 22339 36771
rect 22281 36731 22339 36737
rect 22465 36771 22523 36777
rect 22465 36737 22477 36771
rect 22511 36737 22523 36771
rect 22465 36731 22523 36737
rect 22370 36700 22376 36712
rect 21008 36672 22376 36700
rect 20901 36663 20959 36669
rect 16850 36592 16856 36644
rect 16908 36592 16914 36644
rect 17037 36635 17095 36641
rect 17037 36601 17049 36635
rect 17083 36632 17095 36635
rect 17126 36632 17132 36644
rect 17083 36604 17132 36632
rect 17083 36601 17095 36604
rect 17037 36595 17095 36601
rect 17126 36592 17132 36604
rect 17184 36632 17190 36644
rect 17773 36635 17831 36641
rect 17773 36632 17785 36635
rect 17184 36604 17785 36632
rect 17184 36592 17190 36604
rect 17773 36601 17785 36604
rect 17819 36632 17831 36635
rect 18785 36635 18843 36641
rect 18785 36632 18797 36635
rect 17819 36604 18797 36632
rect 17819 36601 17831 36604
rect 17773 36595 17831 36601
rect 18785 36601 18797 36604
rect 18831 36632 18843 36635
rect 19426 36632 19432 36644
rect 18831 36604 19432 36632
rect 18831 36601 18843 36604
rect 18785 36595 18843 36601
rect 19426 36592 19432 36604
rect 19484 36592 19490 36644
rect 19886 36592 19892 36644
rect 19944 36632 19950 36644
rect 20916 36632 20944 36663
rect 22370 36660 22376 36672
rect 22428 36660 22434 36712
rect 21910 36632 21916 36644
rect 19944 36604 21916 36632
rect 19944 36592 19950 36604
rect 21910 36592 21916 36604
rect 21968 36592 21974 36644
rect 22480 36632 22508 36731
rect 23658 36728 23664 36780
rect 23716 36768 23722 36780
rect 24213 36771 24271 36777
rect 24213 36768 24225 36771
rect 23716 36740 24225 36768
rect 23716 36728 23722 36740
rect 24213 36737 24225 36740
rect 24259 36737 24271 36771
rect 25038 36768 25044 36780
rect 24999 36740 25044 36768
rect 24213 36731 24271 36737
rect 25038 36728 25044 36740
rect 25096 36728 25102 36780
rect 26326 36768 26332 36780
rect 26287 36740 26332 36768
rect 26326 36728 26332 36740
rect 26384 36728 26390 36780
rect 26418 36728 26424 36780
rect 26476 36768 26482 36780
rect 27706 36777 27712 36780
rect 27704 36768 27712 36777
rect 26476 36740 26521 36768
rect 27667 36740 27712 36768
rect 26476 36728 26482 36740
rect 27704 36731 27712 36740
rect 27706 36728 27712 36731
rect 27764 36728 27770 36780
rect 27801 36771 27859 36777
rect 27801 36737 27813 36771
rect 27847 36737 27859 36771
rect 27801 36731 27859 36737
rect 24670 36660 24676 36712
rect 24728 36700 24734 36712
rect 24949 36703 25007 36709
rect 24949 36700 24961 36703
rect 24728 36672 24961 36700
rect 24728 36660 24734 36672
rect 24949 36669 24961 36672
rect 24995 36669 25007 36703
rect 24949 36663 25007 36669
rect 26050 36660 26056 36712
rect 26108 36700 26114 36712
rect 26145 36703 26203 36709
rect 26145 36700 26157 36703
rect 26108 36672 26157 36700
rect 26108 36660 26114 36672
rect 26145 36669 26157 36672
rect 26191 36669 26203 36703
rect 26145 36663 26203 36669
rect 26326 36632 26332 36644
rect 22480 36604 26332 36632
rect 26326 36592 26332 36604
rect 26384 36592 26390 36644
rect 16666 36564 16672 36576
rect 16627 36536 16672 36564
rect 16666 36524 16672 36536
rect 16724 36524 16730 36576
rect 18414 36524 18420 36576
rect 18472 36564 18478 36576
rect 18877 36567 18935 36573
rect 18877 36564 18889 36567
rect 18472 36536 18889 36564
rect 18472 36524 18478 36536
rect 18877 36533 18889 36536
rect 18923 36564 18935 36567
rect 19521 36567 19579 36573
rect 19521 36564 19533 36567
rect 18923 36536 19533 36564
rect 18923 36533 18935 36536
rect 18877 36527 18935 36533
rect 19521 36533 19533 36536
rect 19567 36533 19579 36567
rect 20806 36564 20812 36576
rect 20767 36536 20812 36564
rect 19521 36527 19579 36533
rect 20806 36524 20812 36536
rect 20864 36524 20870 36576
rect 21821 36567 21879 36573
rect 21821 36533 21833 36567
rect 21867 36564 21879 36567
rect 22186 36564 22192 36576
rect 21867 36536 22192 36564
rect 21867 36533 21879 36536
rect 21821 36527 21879 36533
rect 22186 36524 22192 36536
rect 22244 36524 22250 36576
rect 26142 36524 26148 36576
rect 26200 36564 26206 36576
rect 26237 36567 26295 36573
rect 26237 36564 26249 36567
rect 26200 36536 26249 36564
rect 26200 36524 26206 36536
rect 26237 36533 26249 36536
rect 26283 36533 26295 36567
rect 26237 36527 26295 36533
rect 27430 36524 27436 36576
rect 27488 36564 27494 36576
rect 27525 36567 27583 36573
rect 27525 36564 27537 36567
rect 27488 36536 27537 36564
rect 27488 36524 27494 36536
rect 27525 36533 27537 36536
rect 27571 36533 27583 36567
rect 27816 36564 27844 36731
rect 27890 36728 27896 36780
rect 27948 36768 27954 36780
rect 28074 36768 28080 36780
rect 27948 36740 27993 36768
rect 28035 36740 28080 36768
rect 27948 36728 27954 36740
rect 28074 36728 28080 36740
rect 28132 36728 28138 36780
rect 28644 36777 28672 36808
rect 28718 36796 28724 36848
rect 28776 36836 28782 36848
rect 28776 36808 28948 36836
rect 28776 36796 28782 36808
rect 28169 36771 28227 36777
rect 28169 36737 28181 36771
rect 28215 36737 28227 36771
rect 28169 36731 28227 36737
rect 28629 36771 28687 36777
rect 28629 36737 28641 36771
rect 28675 36737 28687 36771
rect 28810 36768 28816 36780
rect 28771 36740 28816 36768
rect 28629 36731 28687 36737
rect 28184 36700 28212 36731
rect 28810 36728 28816 36740
rect 28868 36728 28874 36780
rect 28920 36777 28948 36808
rect 31220 36777 31248 36876
rect 33229 36873 33241 36876
rect 33275 36873 33287 36907
rect 33229 36867 33287 36873
rect 28905 36771 28963 36777
rect 28905 36737 28917 36771
rect 28951 36737 28963 36771
rect 28905 36731 28963 36737
rect 29181 36771 29239 36777
rect 29181 36737 29193 36771
rect 29227 36737 29239 36771
rect 29181 36731 29239 36737
rect 30949 36771 31007 36777
rect 30949 36737 30961 36771
rect 30995 36768 31007 36771
rect 31205 36771 31263 36777
rect 30995 36740 31156 36768
rect 30995 36737 31007 36740
rect 30949 36731 31007 36737
rect 28721 36703 28779 36709
rect 28721 36700 28733 36703
rect 28184 36672 28733 36700
rect 28721 36669 28733 36672
rect 28767 36669 28779 36703
rect 29196 36700 29224 36731
rect 28721 36663 28779 36669
rect 28828 36672 29224 36700
rect 31128 36700 31156 36740
rect 31205 36737 31217 36771
rect 31251 36737 31263 36771
rect 32306 36768 32312 36780
rect 32267 36740 32312 36768
rect 31205 36731 31263 36737
rect 32306 36728 32312 36740
rect 32364 36728 32370 36780
rect 32125 36703 32183 36709
rect 32125 36700 32137 36703
rect 31128 36672 32137 36700
rect 28350 36564 28356 36576
rect 27816 36536 28356 36564
rect 27525 36527 27583 36533
rect 28350 36524 28356 36536
rect 28408 36564 28414 36576
rect 28828 36564 28856 36672
rect 32125 36669 32137 36672
rect 32171 36669 32183 36703
rect 32125 36663 32183 36669
rect 32585 36703 32643 36709
rect 32585 36669 32597 36703
rect 32631 36700 32643 36703
rect 32950 36700 32956 36712
rect 32631 36672 32956 36700
rect 32631 36669 32643 36672
rect 32585 36663 32643 36669
rect 32214 36632 32220 36644
rect 31726 36604 32220 36632
rect 28408 36536 28856 36564
rect 28408 36524 28414 36536
rect 28902 36524 28908 36576
rect 28960 36564 28966 36576
rect 29089 36567 29147 36573
rect 29089 36564 29101 36567
rect 28960 36536 29101 36564
rect 28960 36524 28966 36536
rect 29089 36533 29101 36536
rect 29135 36533 29147 36567
rect 29089 36527 29147 36533
rect 29825 36567 29883 36573
rect 29825 36533 29837 36567
rect 29871 36564 29883 36567
rect 31294 36564 31300 36576
rect 29871 36536 31300 36564
rect 29871 36533 29883 36536
rect 29825 36527 29883 36533
rect 31294 36524 31300 36536
rect 31352 36564 31358 36576
rect 31726 36564 31754 36604
rect 32214 36592 32220 36604
rect 32272 36632 32278 36644
rect 32600 36632 32628 36663
rect 32950 36660 32956 36672
rect 33008 36660 33014 36712
rect 33244 36700 33272 36867
rect 34146 36864 34152 36916
rect 34204 36904 34210 36916
rect 34977 36907 35035 36913
rect 34977 36904 34989 36907
rect 34204 36876 34989 36904
rect 34204 36864 34210 36876
rect 34977 36873 34989 36876
rect 35023 36873 35035 36907
rect 34977 36867 35035 36873
rect 40770 36864 40776 36916
rect 40828 36904 40834 36916
rect 41325 36907 41383 36913
rect 41325 36904 41337 36907
rect 40828 36876 41337 36904
rect 40828 36864 40834 36876
rect 41325 36873 41337 36876
rect 41371 36873 41383 36907
rect 41598 36904 41604 36916
rect 41559 36876 41604 36904
rect 41325 36867 41383 36873
rect 41598 36864 41604 36876
rect 41656 36864 41662 36916
rect 41690 36864 41696 36916
rect 41748 36904 41754 36916
rect 42426 36904 42432 36916
rect 41748 36876 41793 36904
rect 42387 36876 42432 36904
rect 41748 36864 41754 36876
rect 42426 36864 42432 36876
rect 42484 36864 42490 36916
rect 43254 36904 43260 36916
rect 43215 36876 43260 36904
rect 43254 36864 43260 36876
rect 43312 36864 43318 36916
rect 34241 36839 34299 36845
rect 34241 36805 34253 36839
rect 34287 36836 34299 36839
rect 34514 36836 34520 36848
rect 34287 36808 34520 36836
rect 34287 36805 34299 36808
rect 34241 36799 34299 36805
rect 34514 36796 34520 36808
rect 34572 36796 34578 36848
rect 35986 36836 35992 36848
rect 34624 36808 35992 36836
rect 33321 36771 33379 36777
rect 33321 36737 33333 36771
rect 33367 36768 33379 36771
rect 34624 36768 34652 36808
rect 35986 36796 35992 36808
rect 36044 36836 36050 36848
rect 37369 36839 37427 36845
rect 37369 36836 37381 36839
rect 36044 36808 37381 36836
rect 36044 36796 36050 36808
rect 37369 36805 37381 36808
rect 37415 36805 37427 36839
rect 37369 36799 37427 36805
rect 37553 36839 37611 36845
rect 37553 36805 37565 36839
rect 37599 36836 37611 36839
rect 39942 36836 39948 36848
rect 37599 36808 39948 36836
rect 37599 36805 37611 36808
rect 37553 36799 37611 36805
rect 38672 36780 38700 36808
rect 39942 36796 39948 36808
rect 40000 36796 40006 36848
rect 41414 36796 41420 36848
rect 41472 36836 41478 36848
rect 41472 36808 41920 36836
rect 41472 36796 41478 36808
rect 33367 36740 34652 36768
rect 33367 36737 33379 36740
rect 33321 36731 33379 36737
rect 34698 36728 34704 36780
rect 34756 36768 34762 36780
rect 34885 36771 34943 36777
rect 34885 36768 34897 36771
rect 34756 36740 34897 36768
rect 34756 36728 34762 36740
rect 34885 36737 34897 36740
rect 34931 36737 34943 36771
rect 34885 36731 34943 36737
rect 35161 36771 35219 36777
rect 35161 36737 35173 36771
rect 35207 36768 35219 36771
rect 35434 36768 35440 36780
rect 35207 36740 35440 36768
rect 35207 36737 35219 36740
rect 35161 36731 35219 36737
rect 35434 36728 35440 36740
rect 35492 36728 35498 36780
rect 38654 36768 38660 36780
rect 38567 36740 38660 36768
rect 38654 36728 38660 36740
rect 38712 36728 38718 36780
rect 38930 36777 38936 36780
rect 38924 36768 38936 36777
rect 38891 36740 38936 36768
rect 38924 36731 38936 36740
rect 38930 36728 38936 36731
rect 38988 36728 38994 36780
rect 41892 36777 41920 36808
rect 41966 36796 41972 36848
rect 42024 36836 42030 36848
rect 42581 36839 42639 36845
rect 42581 36836 42593 36839
rect 42024 36808 42593 36836
rect 42024 36796 42030 36808
rect 42581 36805 42593 36808
rect 42627 36805 42639 36839
rect 42581 36799 42639 36805
rect 42797 36839 42855 36845
rect 42797 36805 42809 36839
rect 42843 36805 42855 36839
rect 42797 36799 42855 36805
rect 41509 36771 41567 36777
rect 41509 36737 41521 36771
rect 41555 36737 41567 36771
rect 41509 36731 41567 36737
rect 41877 36771 41935 36777
rect 41877 36737 41889 36771
rect 41923 36768 41935 36771
rect 42812 36768 42840 36799
rect 43533 36771 43591 36777
rect 43533 36768 43545 36771
rect 41923 36740 43545 36768
rect 41923 36737 41935 36740
rect 41877 36731 41935 36737
rect 43533 36737 43545 36740
rect 43579 36768 43591 36771
rect 43806 36768 43812 36780
rect 43579 36740 43812 36768
rect 43579 36737 43591 36740
rect 43533 36731 43591 36737
rect 36170 36700 36176 36712
rect 33244 36672 36176 36700
rect 36170 36660 36176 36672
rect 36228 36660 36234 36712
rect 41524 36700 41552 36731
rect 43806 36728 43812 36740
rect 43864 36728 43870 36780
rect 41966 36700 41972 36712
rect 41524 36672 41972 36700
rect 41966 36660 41972 36672
rect 42024 36660 42030 36712
rect 42886 36660 42892 36712
rect 42944 36700 42950 36712
rect 43257 36703 43315 36709
rect 43257 36700 43269 36703
rect 42944 36672 43269 36700
rect 42944 36660 42950 36672
rect 43257 36669 43269 36672
rect 43303 36669 43315 36703
rect 43257 36663 43315 36669
rect 32272 36604 32628 36632
rect 33873 36635 33931 36641
rect 32272 36592 32278 36604
rect 33873 36601 33885 36635
rect 33919 36601 33931 36635
rect 35345 36635 35403 36641
rect 35345 36632 35357 36635
rect 33873 36595 33931 36601
rect 34256 36604 35357 36632
rect 32490 36564 32496 36576
rect 31352 36536 31754 36564
rect 32451 36536 32496 36564
rect 31352 36524 31358 36536
rect 32490 36524 32496 36536
rect 32548 36564 32554 36576
rect 33888 36564 33916 36595
rect 34256 36573 34284 36604
rect 35345 36601 35357 36604
rect 35391 36601 35403 36635
rect 35345 36595 35403 36601
rect 42058 36592 42064 36644
rect 42116 36632 42122 36644
rect 43441 36635 43499 36641
rect 43441 36632 43453 36635
rect 42116 36604 43453 36632
rect 42116 36592 42122 36604
rect 43441 36601 43453 36604
rect 43487 36601 43499 36635
rect 43441 36595 43499 36601
rect 32548 36536 33916 36564
rect 34241 36567 34299 36573
rect 32548 36524 32554 36536
rect 34241 36533 34253 36567
rect 34287 36533 34299 36567
rect 34241 36527 34299 36533
rect 34425 36567 34483 36573
rect 34425 36533 34437 36567
rect 34471 36564 34483 36567
rect 34790 36564 34796 36576
rect 34471 36536 34796 36564
rect 34471 36533 34483 36536
rect 34425 36527 34483 36533
rect 34790 36524 34796 36536
rect 34848 36524 34854 36576
rect 40034 36564 40040 36576
rect 39995 36536 40040 36564
rect 40034 36524 40040 36536
rect 40092 36524 40098 36576
rect 41690 36524 41696 36576
rect 41748 36564 41754 36576
rect 42613 36567 42671 36573
rect 42613 36564 42625 36567
rect 41748 36536 42625 36564
rect 41748 36524 41754 36536
rect 42613 36533 42625 36536
rect 42659 36533 42671 36567
rect 44174 36564 44180 36576
rect 44135 36536 44180 36564
rect 42613 36527 42671 36533
rect 44174 36524 44180 36536
rect 44232 36524 44238 36576
rect 1104 36474 44896 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 44896 36474
rect 1104 36400 44896 36422
rect 18598 36360 18604 36372
rect 18559 36332 18604 36360
rect 18598 36320 18604 36332
rect 18656 36320 18662 36372
rect 20530 36360 20536 36372
rect 20180 36332 20536 36360
rect 20070 36292 20076 36304
rect 20031 36264 20076 36292
rect 20070 36252 20076 36264
rect 20128 36252 20134 36304
rect 20180 36301 20208 36332
rect 20530 36320 20536 36332
rect 20588 36360 20594 36372
rect 21542 36360 21548 36372
rect 20588 36332 21548 36360
rect 20588 36320 20594 36332
rect 21542 36320 21548 36332
rect 21600 36320 21606 36372
rect 21637 36363 21695 36369
rect 21637 36329 21649 36363
rect 21683 36360 21695 36363
rect 21726 36360 21732 36372
rect 21683 36332 21732 36360
rect 21683 36329 21695 36332
rect 21637 36323 21695 36329
rect 21726 36320 21732 36332
rect 21784 36320 21790 36372
rect 22094 36320 22100 36372
rect 22152 36360 22158 36372
rect 26234 36360 26240 36372
rect 22152 36332 22197 36360
rect 26195 36332 26240 36360
rect 22152 36320 22158 36332
rect 26234 36320 26240 36332
rect 26292 36320 26298 36372
rect 27246 36320 27252 36372
rect 27304 36360 27310 36372
rect 27798 36360 27804 36372
rect 27304 36332 27804 36360
rect 27304 36320 27310 36332
rect 27798 36320 27804 36332
rect 27856 36320 27862 36372
rect 31113 36363 31171 36369
rect 31113 36329 31125 36363
rect 31159 36360 31171 36363
rect 32306 36360 32312 36372
rect 31159 36332 32312 36360
rect 31159 36329 31171 36332
rect 31113 36323 31171 36329
rect 32306 36320 32312 36332
rect 32364 36320 32370 36372
rect 33594 36320 33600 36372
rect 33652 36360 33658 36372
rect 33965 36363 34023 36369
rect 33965 36360 33977 36363
rect 33652 36332 33977 36360
rect 33652 36320 33658 36332
rect 33965 36329 33977 36332
rect 34011 36360 34023 36363
rect 34238 36360 34244 36372
rect 34011 36332 34244 36360
rect 34011 36329 34023 36332
rect 33965 36323 34023 36329
rect 34238 36320 34244 36332
rect 34296 36360 34302 36372
rect 34793 36363 34851 36369
rect 34793 36360 34805 36363
rect 34296 36332 34805 36360
rect 34296 36320 34302 36332
rect 34793 36329 34805 36332
rect 34839 36360 34851 36363
rect 35434 36360 35440 36372
rect 34839 36332 35440 36360
rect 34839 36329 34851 36332
rect 34793 36323 34851 36329
rect 35434 36320 35440 36332
rect 35492 36320 35498 36372
rect 39117 36363 39175 36369
rect 39117 36329 39129 36363
rect 39163 36360 39175 36363
rect 40034 36360 40040 36372
rect 39163 36332 40040 36360
rect 39163 36329 39175 36332
rect 39117 36323 39175 36329
rect 40034 36320 40040 36332
rect 40092 36320 40098 36372
rect 40218 36360 40224 36372
rect 40179 36332 40224 36360
rect 40218 36320 40224 36332
rect 40276 36320 40282 36372
rect 20165 36295 20223 36301
rect 20165 36261 20177 36295
rect 20211 36261 20223 36295
rect 21818 36292 21824 36304
rect 20165 36255 20223 36261
rect 20272 36264 21824 36292
rect 18690 36224 18696 36236
rect 18651 36196 18696 36224
rect 18690 36184 18696 36196
rect 18748 36184 18754 36236
rect 15838 36116 15844 36168
rect 15896 36156 15902 36168
rect 15933 36159 15991 36165
rect 15933 36156 15945 36159
rect 15896 36128 15945 36156
rect 15896 36116 15902 36128
rect 15933 36125 15945 36128
rect 15979 36125 15991 36159
rect 15933 36119 15991 36125
rect 16200 36159 16258 36165
rect 16200 36125 16212 36159
rect 16246 36156 16258 36159
rect 16666 36156 16672 36168
rect 16246 36128 16672 36156
rect 16246 36125 16258 36128
rect 16200 36119 16258 36125
rect 16666 36116 16672 36128
rect 16724 36116 16730 36168
rect 17770 36156 17776 36168
rect 17731 36128 17776 36156
rect 17770 36116 17776 36128
rect 17828 36116 17834 36168
rect 18414 36156 18420 36168
rect 18375 36128 18420 36156
rect 18414 36116 18420 36128
rect 18472 36116 18478 36168
rect 18509 36159 18567 36165
rect 18509 36125 18521 36159
rect 18555 36156 18567 36159
rect 19797 36159 19855 36165
rect 19797 36156 19809 36159
rect 18555 36128 19809 36156
rect 18555 36125 18567 36128
rect 18509 36119 18567 36125
rect 19797 36125 19809 36128
rect 19843 36125 19855 36159
rect 19797 36119 19855 36125
rect 19886 36116 19892 36168
rect 19944 36156 19950 36168
rect 20272 36165 20300 36264
rect 21818 36252 21824 36264
rect 21876 36252 21882 36304
rect 26326 36252 26332 36304
rect 26384 36292 26390 36304
rect 26384 36264 27200 36292
rect 26384 36252 26390 36264
rect 20806 36184 20812 36236
rect 20864 36224 20870 36236
rect 20864 36196 22784 36224
rect 20864 36184 20870 36196
rect 19981 36159 20039 36165
rect 19981 36156 19993 36159
rect 19944 36128 19993 36156
rect 19944 36116 19950 36128
rect 19981 36125 19993 36128
rect 20027 36125 20039 36159
rect 19981 36119 20039 36125
rect 20257 36159 20315 36165
rect 20257 36125 20269 36159
rect 20303 36125 20315 36159
rect 20990 36156 20996 36168
rect 20951 36128 20996 36156
rect 20257 36119 20315 36125
rect 20990 36116 20996 36128
rect 21048 36116 21054 36168
rect 21086 36159 21144 36165
rect 21086 36125 21098 36159
rect 21132 36125 21144 36159
rect 21086 36119 21144 36125
rect 17586 36088 17592 36100
rect 17328 36060 17592 36088
rect 17328 36029 17356 36060
rect 17586 36048 17592 36060
rect 17644 36088 17650 36100
rect 18598 36088 18604 36100
rect 17644 36060 18604 36088
rect 17644 36048 17650 36060
rect 18598 36048 18604 36060
rect 18656 36048 18662 36100
rect 20714 36048 20720 36100
rect 20772 36088 20778 36100
rect 21101 36088 21129 36119
rect 21174 36116 21180 36168
rect 21232 36156 21238 36168
rect 21458 36159 21516 36165
rect 21458 36156 21470 36159
rect 21232 36128 21470 36156
rect 21232 36116 21238 36128
rect 21458 36125 21470 36128
rect 21504 36125 21516 36159
rect 21458 36119 21516 36125
rect 22002 36116 22008 36168
rect 22060 36156 22066 36168
rect 22235 36159 22293 36165
rect 22235 36156 22247 36159
rect 22060 36128 22247 36156
rect 22060 36116 22066 36128
rect 22235 36125 22247 36128
rect 22281 36125 22293 36159
rect 22235 36119 22293 36125
rect 22370 36116 22376 36168
rect 22428 36156 22434 36168
rect 22646 36156 22652 36168
rect 22428 36128 22473 36156
rect 22607 36128 22652 36156
rect 22428 36116 22434 36128
rect 22646 36116 22652 36128
rect 22704 36116 22710 36168
rect 22756 36165 22784 36196
rect 22741 36159 22799 36165
rect 22741 36125 22753 36159
rect 22787 36125 22799 36159
rect 23474 36156 23480 36168
rect 23435 36128 23480 36156
rect 22741 36119 22799 36125
rect 23474 36116 23480 36128
rect 23532 36116 23538 36168
rect 25685 36159 25743 36165
rect 25685 36125 25697 36159
rect 25731 36125 25743 36159
rect 26142 36156 26148 36168
rect 26103 36128 26148 36156
rect 25685 36119 25743 36125
rect 20772 36060 21129 36088
rect 21269 36091 21327 36097
rect 20772 36048 20778 36060
rect 21269 36057 21281 36091
rect 21315 36057 21327 36091
rect 21269 36051 21327 36057
rect 21361 36091 21419 36097
rect 21361 36057 21373 36091
rect 21407 36088 21419 36091
rect 21910 36088 21916 36100
rect 21407 36060 21916 36088
rect 21407 36057 21419 36060
rect 21361 36051 21419 36057
rect 17313 36023 17371 36029
rect 17313 35989 17325 36023
rect 17359 35989 17371 36023
rect 17313 35983 17371 35989
rect 17865 36023 17923 36029
rect 17865 35989 17877 36023
rect 17911 36020 17923 36023
rect 20622 36020 20628 36032
rect 17911 35992 20628 36020
rect 17911 35989 17923 35992
rect 17865 35983 17923 35989
rect 20622 35980 20628 35992
rect 20680 36020 20686 36032
rect 21284 36020 21312 36051
rect 21910 36048 21916 36060
rect 21968 36048 21974 36100
rect 22465 36091 22523 36097
rect 22465 36057 22477 36091
rect 22511 36057 22523 36091
rect 25700 36088 25728 36119
rect 26142 36116 26148 36128
rect 26200 36116 26206 36168
rect 26326 36156 26332 36168
rect 26287 36128 26332 36156
rect 26326 36116 26332 36128
rect 26384 36116 26390 36168
rect 27172 36165 27200 36264
rect 27522 36252 27528 36304
rect 27580 36292 27586 36304
rect 27706 36292 27712 36304
rect 27580 36264 27712 36292
rect 27580 36252 27586 36264
rect 27706 36252 27712 36264
rect 27764 36292 27770 36304
rect 27764 36264 28304 36292
rect 27764 36252 27770 36264
rect 27157 36159 27215 36165
rect 27157 36125 27169 36159
rect 27203 36125 27215 36159
rect 27320 36159 27378 36165
rect 27320 36156 27332 36159
rect 27157 36119 27215 36125
rect 27264 36128 27332 36156
rect 26050 36088 26056 36100
rect 25700 36060 26056 36088
rect 22465 36051 22523 36057
rect 20680 35992 21312 36020
rect 20680 35980 20686 35992
rect 21542 35980 21548 36032
rect 21600 36020 21606 36032
rect 22480 36020 22508 36051
rect 26050 36048 26056 36060
rect 26108 36088 26114 36100
rect 27264 36088 27292 36128
rect 27320 36125 27332 36128
rect 27366 36125 27378 36159
rect 27430 36154 27436 36206
rect 27488 36154 27494 36206
rect 27545 36159 27603 36165
rect 27545 36158 27557 36159
rect 27320 36119 27378 36125
rect 27436 36122 27448 36154
rect 27482 36122 27494 36154
rect 27540 36128 27557 36158
rect 27436 36116 27494 36122
rect 27545 36125 27557 36128
rect 27591 36158 27603 36159
rect 27591 36156 27660 36158
rect 27798 36156 27804 36168
rect 27591 36130 27804 36156
rect 27591 36125 27603 36130
rect 27632 36128 27804 36130
rect 27545 36119 27603 36125
rect 27798 36116 27804 36128
rect 27856 36116 27862 36168
rect 28276 36165 28304 36264
rect 32490 36252 32496 36304
rect 32548 36292 32554 36304
rect 33781 36295 33839 36301
rect 33781 36292 33793 36295
rect 32548 36264 33793 36292
rect 32548 36252 32554 36264
rect 33781 36261 33793 36264
rect 33827 36261 33839 36295
rect 33781 36255 33839 36261
rect 38013 36295 38071 36301
rect 38013 36261 38025 36295
rect 38059 36292 38071 36295
rect 38746 36292 38752 36304
rect 38059 36264 38752 36292
rect 38059 36261 38071 36264
rect 38013 36255 38071 36261
rect 38746 36252 38752 36264
rect 38804 36292 38810 36304
rect 39301 36295 39359 36301
rect 38804 36264 39160 36292
rect 38804 36252 38810 36264
rect 33321 36227 33379 36233
rect 33321 36193 33333 36227
rect 33367 36224 33379 36227
rect 34514 36224 34520 36236
rect 33367 36196 34520 36224
rect 33367 36193 33379 36196
rect 33321 36187 33379 36193
rect 34514 36184 34520 36196
rect 34572 36184 34578 36236
rect 36170 36224 36176 36236
rect 36131 36196 36176 36224
rect 36170 36184 36176 36196
rect 36228 36224 36234 36236
rect 36633 36227 36691 36233
rect 36633 36224 36645 36227
rect 36228 36196 36645 36224
rect 36228 36184 36234 36196
rect 36633 36193 36645 36196
rect 36679 36193 36691 36227
rect 36633 36187 36691 36193
rect 38657 36227 38715 36233
rect 38657 36193 38669 36227
rect 38703 36224 38715 36227
rect 38838 36224 38844 36236
rect 38703 36196 38844 36224
rect 38703 36193 38715 36196
rect 38657 36187 38715 36193
rect 38838 36184 38844 36196
rect 38896 36184 38902 36236
rect 28261 36159 28319 36165
rect 28261 36125 28273 36159
rect 28307 36125 28319 36159
rect 28261 36119 28319 36125
rect 30929 36159 30987 36165
rect 30929 36125 30941 36159
rect 30975 36156 30987 36159
rect 31018 36156 31024 36168
rect 30975 36128 31024 36156
rect 30975 36125 30987 36128
rect 30929 36119 30987 36125
rect 31018 36116 31024 36128
rect 31076 36116 31082 36168
rect 31294 36156 31300 36168
rect 31255 36128 31300 36156
rect 31294 36116 31300 36128
rect 31352 36116 31358 36168
rect 31389 36159 31447 36165
rect 31389 36125 31401 36159
rect 31435 36156 31447 36159
rect 32490 36156 32496 36168
rect 31435 36128 32496 36156
rect 31435 36125 31447 36128
rect 31389 36119 31447 36125
rect 32490 36116 32496 36128
rect 32548 36116 32554 36168
rect 38749 36159 38807 36165
rect 38749 36125 38761 36159
rect 38795 36156 38807 36159
rect 38930 36156 38936 36168
rect 38795 36128 38936 36156
rect 38795 36125 38807 36128
rect 38749 36119 38807 36125
rect 38930 36116 38936 36128
rect 38988 36116 38994 36168
rect 39132 36165 39160 36264
rect 39301 36261 39313 36295
rect 39347 36261 39359 36295
rect 40052 36292 40080 36320
rect 40494 36292 40500 36304
rect 40052 36264 40500 36292
rect 39301 36255 39359 36261
rect 39316 36224 39344 36255
rect 40494 36252 40500 36264
rect 40552 36252 40558 36304
rect 40512 36224 40540 36252
rect 41049 36227 41107 36233
rect 41049 36224 41061 36227
rect 39316 36196 40264 36224
rect 40512 36196 41061 36224
rect 39117 36159 39175 36165
rect 39117 36125 39129 36159
rect 39163 36125 39175 36159
rect 40034 36156 40040 36168
rect 39995 36128 40040 36156
rect 39117 36119 39175 36125
rect 40034 36116 40040 36128
rect 40092 36116 40098 36168
rect 40236 36165 40264 36196
rect 41049 36193 41061 36196
rect 41095 36193 41107 36227
rect 42702 36224 42708 36236
rect 42663 36196 42708 36224
rect 41049 36187 41107 36193
rect 42702 36184 42708 36196
rect 42760 36184 42766 36236
rect 44174 36224 44180 36236
rect 44135 36196 44180 36224
rect 44174 36184 44180 36196
rect 44232 36184 44238 36236
rect 40221 36159 40279 36165
rect 40221 36125 40233 36159
rect 40267 36125 40279 36159
rect 40862 36156 40868 36168
rect 40823 36128 40868 36156
rect 40221 36119 40279 36125
rect 40862 36116 40868 36128
rect 40920 36116 40926 36168
rect 41506 36156 41512 36168
rect 41467 36128 41512 36156
rect 41506 36116 41512 36128
rect 41564 36116 41570 36168
rect 41693 36159 41751 36165
rect 41693 36125 41705 36159
rect 41739 36156 41751 36159
rect 42058 36156 42064 36168
rect 41739 36128 42064 36156
rect 41739 36125 41751 36128
rect 41693 36119 41751 36125
rect 42058 36116 42064 36128
rect 42116 36116 42122 36168
rect 26108 36060 27292 36088
rect 33137 36091 33195 36097
rect 26108 36048 26114 36060
rect 33137 36057 33149 36091
rect 33183 36088 33195 36091
rect 33318 36088 33324 36100
rect 33183 36060 33324 36088
rect 33183 36057 33195 36060
rect 33137 36051 33195 36057
rect 33318 36048 33324 36060
rect 33376 36048 33382 36100
rect 33686 36048 33692 36100
rect 33744 36088 33750 36100
rect 34146 36088 34152 36100
rect 33744 36060 34152 36088
rect 33744 36048 33750 36060
rect 34146 36048 34152 36060
rect 34204 36048 34210 36100
rect 35894 36048 35900 36100
rect 35952 36097 35958 36100
rect 35952 36088 35964 36097
rect 35952 36060 35997 36088
rect 35952 36051 35964 36060
rect 35952 36048 35958 36051
rect 36722 36048 36728 36100
rect 36780 36088 36786 36100
rect 36878 36091 36936 36097
rect 36878 36088 36890 36091
rect 36780 36060 36890 36088
rect 36780 36048 36786 36060
rect 36878 36057 36890 36060
rect 36924 36057 36936 36091
rect 43990 36088 43996 36100
rect 43951 36060 43996 36088
rect 36878 36051 36936 36057
rect 43990 36048 43996 36060
rect 44048 36048 44054 36100
rect 21600 35992 22508 36020
rect 23661 36023 23719 36029
rect 21600 35980 21606 35992
rect 23661 35989 23673 36023
rect 23707 36020 23719 36023
rect 23842 36020 23848 36032
rect 23707 35992 23848 36020
rect 23707 35989 23719 35992
rect 23661 35983 23719 35989
rect 23842 35980 23848 35992
rect 23900 35980 23906 36032
rect 25590 36020 25596 36032
rect 25551 35992 25596 36020
rect 25590 35980 25596 35992
rect 25648 35980 25654 36032
rect 27430 35980 27436 36032
rect 27488 36020 27494 36032
rect 27801 36023 27859 36029
rect 27801 36020 27813 36023
rect 27488 35992 27813 36020
rect 27488 35980 27494 35992
rect 27801 35989 27813 35992
rect 27847 35989 27859 36023
rect 27801 35983 27859 35989
rect 28074 35980 28080 36032
rect 28132 36020 28138 36032
rect 28353 36023 28411 36029
rect 28353 36020 28365 36023
rect 28132 35992 28365 36020
rect 28132 35980 28138 35992
rect 28353 35989 28365 35992
rect 28399 36020 28411 36023
rect 29546 36020 29552 36032
rect 28399 35992 29552 36020
rect 28399 35989 28411 35992
rect 28353 35983 28411 35989
rect 29546 35980 29552 35992
rect 29604 35980 29610 36032
rect 33949 36023 34007 36029
rect 33949 35989 33961 36023
rect 33995 36020 34007 36023
rect 34698 36020 34704 36032
rect 33995 35992 34704 36020
rect 33995 35989 34007 35992
rect 33949 35983 34007 35989
rect 34698 35980 34704 35992
rect 34756 35980 34762 36032
rect 39850 36020 39856 36032
rect 39811 35992 39856 36020
rect 39850 35980 39856 35992
rect 39908 35980 39914 36032
rect 40678 36020 40684 36032
rect 40639 35992 40684 36020
rect 40678 35980 40684 35992
rect 40736 35980 40742 36032
rect 41598 36020 41604 36032
rect 41559 35992 41604 36020
rect 41598 35980 41604 35992
rect 41656 35980 41662 36032
rect 1104 35930 44896 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 44896 35930
rect 1104 35856 44896 35878
rect 19061 35819 19119 35825
rect 19061 35785 19073 35819
rect 19107 35816 19119 35819
rect 20438 35816 20444 35828
rect 19107 35788 20444 35816
rect 19107 35785 19119 35788
rect 19061 35779 19119 35785
rect 20438 35776 20444 35788
rect 20496 35776 20502 35828
rect 21910 35776 21916 35828
rect 21968 35816 21974 35828
rect 22738 35816 22744 35828
rect 21968 35788 22744 35816
rect 21968 35776 21974 35788
rect 22738 35776 22744 35788
rect 22796 35776 22802 35828
rect 23382 35776 23388 35828
rect 23440 35816 23446 35828
rect 23440 35788 24072 35816
rect 23440 35776 23446 35788
rect 21634 35708 21640 35760
rect 21692 35748 21698 35760
rect 22005 35751 22063 35757
rect 22005 35748 22017 35751
rect 21692 35720 22017 35748
rect 21692 35708 21698 35720
rect 22005 35717 22017 35720
rect 22051 35717 22063 35751
rect 22005 35711 22063 35717
rect 22189 35751 22247 35757
rect 22189 35717 22201 35751
rect 22235 35748 22247 35751
rect 23658 35748 23664 35760
rect 22235 35720 23664 35748
rect 22235 35717 22247 35720
rect 22189 35711 22247 35717
rect 23658 35708 23664 35720
rect 23716 35708 23722 35760
rect 23842 35708 23848 35760
rect 23900 35757 23906 35760
rect 23900 35748 23912 35757
rect 24044 35748 24072 35788
rect 31018 35776 31024 35828
rect 31076 35816 31082 35828
rect 31478 35816 31484 35828
rect 31076 35788 31484 35816
rect 31076 35776 31082 35788
rect 31478 35776 31484 35788
rect 31536 35776 31542 35828
rect 39298 35816 39304 35828
rect 31726 35788 39160 35816
rect 39259 35788 39304 35816
rect 31726 35748 31754 35788
rect 23900 35720 23945 35748
rect 24044 35720 31754 35748
rect 33413 35751 33471 35757
rect 23900 35711 23912 35720
rect 33413 35717 33425 35751
rect 33459 35748 33471 35751
rect 34698 35748 34704 35760
rect 33459 35720 34704 35748
rect 33459 35717 33471 35720
rect 33413 35711 33471 35717
rect 23900 35708 23906 35711
rect 34698 35708 34704 35720
rect 34756 35708 34762 35760
rect 36725 35751 36783 35757
rect 36725 35717 36737 35751
rect 36771 35748 36783 35751
rect 37277 35751 37335 35757
rect 37277 35748 37289 35751
rect 36771 35720 37289 35748
rect 36771 35717 36783 35720
rect 36725 35711 36783 35717
rect 37277 35717 37289 35720
rect 37323 35717 37335 35751
rect 37277 35711 37335 35717
rect 18693 35683 18751 35689
rect 18693 35649 18705 35683
rect 18739 35649 18751 35683
rect 18693 35643 18751 35649
rect 20349 35683 20407 35689
rect 20349 35649 20361 35683
rect 20395 35680 20407 35683
rect 20806 35680 20812 35692
rect 20395 35652 20812 35680
rect 20395 35649 20407 35652
rect 20349 35643 20407 35649
rect 18598 35612 18604 35624
rect 18559 35584 18604 35612
rect 18598 35572 18604 35584
rect 18656 35572 18662 35624
rect 18708 35544 18736 35643
rect 20806 35640 20812 35652
rect 20864 35640 20870 35692
rect 24121 35683 24179 35689
rect 24121 35649 24133 35683
rect 24167 35680 24179 35683
rect 24302 35680 24308 35692
rect 24167 35652 24308 35680
rect 24167 35649 24179 35652
rect 24121 35643 24179 35649
rect 24302 35640 24308 35652
rect 24360 35640 24366 35692
rect 25038 35640 25044 35692
rect 25096 35680 25102 35692
rect 25682 35680 25688 35692
rect 25096 35652 25688 35680
rect 25096 35640 25102 35652
rect 25682 35640 25688 35652
rect 25740 35680 25746 35692
rect 26973 35683 27031 35689
rect 26973 35680 26985 35683
rect 25740 35652 26985 35680
rect 25740 35640 25746 35652
rect 26973 35649 26985 35652
rect 27019 35649 27031 35683
rect 26973 35643 27031 35649
rect 27154 35640 27160 35692
rect 27212 35680 27218 35692
rect 27614 35680 27620 35692
rect 27212 35652 27620 35680
rect 27212 35640 27218 35652
rect 27614 35640 27620 35652
rect 27672 35640 27678 35692
rect 27798 35680 27804 35692
rect 27759 35652 27804 35680
rect 27798 35640 27804 35652
rect 27856 35640 27862 35692
rect 31386 35680 31392 35692
rect 31347 35652 31392 35680
rect 31386 35640 31392 35652
rect 31444 35680 31450 35692
rect 32585 35683 32643 35689
rect 32585 35680 32597 35683
rect 31444 35652 32597 35680
rect 31444 35640 31450 35652
rect 32585 35649 32597 35652
rect 32631 35680 32643 35683
rect 33318 35680 33324 35692
rect 32631 35652 33324 35680
rect 32631 35649 32643 35652
rect 32585 35643 32643 35649
rect 33318 35640 33324 35652
rect 33376 35640 33382 35692
rect 33686 35680 33692 35692
rect 33647 35652 33692 35680
rect 33686 35640 33692 35652
rect 33744 35640 33750 35692
rect 34333 35683 34391 35689
rect 34333 35680 34345 35683
rect 33888 35652 34345 35680
rect 20070 35572 20076 35624
rect 20128 35612 20134 35624
rect 20257 35615 20315 35621
rect 20257 35612 20269 35615
rect 20128 35584 20269 35612
rect 20128 35572 20134 35584
rect 20257 35581 20269 35584
rect 20303 35581 20315 35615
rect 20257 35575 20315 35581
rect 20717 35615 20775 35621
rect 20717 35581 20729 35615
rect 20763 35612 20775 35615
rect 20990 35612 20996 35624
rect 20763 35584 20996 35612
rect 20763 35581 20775 35584
rect 20717 35575 20775 35581
rect 20990 35572 20996 35584
rect 21048 35572 21054 35624
rect 33502 35612 33508 35624
rect 33463 35584 33508 35612
rect 33502 35572 33508 35584
rect 33560 35572 33566 35624
rect 21266 35544 21272 35556
rect 18708 35516 21272 35544
rect 21266 35504 21272 35516
rect 21324 35504 21330 35556
rect 32766 35544 32772 35556
rect 32727 35516 32772 35544
rect 32766 35504 32772 35516
rect 32824 35504 32830 35556
rect 33888 35553 33916 35652
rect 34333 35649 34345 35652
rect 34379 35649 34391 35683
rect 34333 35643 34391 35649
rect 34790 35640 34796 35692
rect 34848 35680 34854 35692
rect 35253 35683 35311 35689
rect 35253 35680 35265 35683
rect 34848 35652 35265 35680
rect 34848 35640 34854 35652
rect 35253 35649 35265 35652
rect 35299 35649 35311 35683
rect 35253 35643 35311 35649
rect 36449 35683 36507 35689
rect 36449 35649 36461 35683
rect 36495 35649 36507 35683
rect 36449 35643 36507 35649
rect 36541 35683 36599 35689
rect 36541 35649 36553 35683
rect 36587 35680 36599 35683
rect 37553 35683 37611 35689
rect 37553 35680 37565 35683
rect 36587 35652 37565 35680
rect 36587 35649 36599 35652
rect 36541 35643 36599 35649
rect 37553 35649 37565 35652
rect 37599 35680 37611 35683
rect 38470 35680 38476 35692
rect 37599 35652 38476 35680
rect 37599 35649 37611 35652
rect 37553 35643 37611 35649
rect 34054 35572 34060 35624
rect 34112 35612 34118 35624
rect 34425 35615 34483 35621
rect 34425 35612 34437 35615
rect 34112 35584 34437 35612
rect 34112 35572 34118 35584
rect 34425 35581 34437 35584
rect 34471 35581 34483 35615
rect 34425 35575 34483 35581
rect 33873 35547 33931 35553
rect 33873 35513 33885 35547
rect 33919 35513 33931 35547
rect 33873 35507 33931 35513
rect 35437 35547 35495 35553
rect 35437 35513 35449 35547
rect 35483 35544 35495 35547
rect 35894 35544 35900 35556
rect 35483 35516 35900 35544
rect 35483 35513 35495 35516
rect 35437 35507 35495 35513
rect 35894 35504 35900 35516
rect 35952 35504 35958 35556
rect 22738 35476 22744 35488
rect 22699 35448 22744 35476
rect 22738 35436 22744 35448
rect 22796 35436 22802 35488
rect 27065 35479 27123 35485
rect 27065 35445 27077 35479
rect 27111 35476 27123 35479
rect 27522 35476 27528 35488
rect 27111 35448 27528 35476
rect 27111 35445 27123 35448
rect 27065 35439 27123 35445
rect 27522 35436 27528 35448
rect 27580 35436 27586 35488
rect 27893 35479 27951 35485
rect 27893 35445 27905 35479
rect 27939 35476 27951 35479
rect 28626 35476 28632 35488
rect 27939 35448 28632 35476
rect 27939 35445 27951 35448
rect 27893 35439 27951 35445
rect 28626 35436 28632 35448
rect 28684 35436 28690 35488
rect 32950 35436 32956 35488
rect 33008 35476 33014 35488
rect 33413 35479 33471 35485
rect 33413 35476 33425 35479
rect 33008 35448 33425 35476
rect 33008 35436 33014 35448
rect 33413 35445 33425 35448
rect 33459 35445 33471 35479
rect 34422 35476 34428 35488
rect 34383 35448 34428 35476
rect 33413 35439 33471 35445
rect 34422 35436 34428 35448
rect 34480 35436 34486 35488
rect 34514 35436 34520 35488
rect 34572 35476 34578 35488
rect 34701 35479 34759 35485
rect 34701 35476 34713 35479
rect 34572 35448 34713 35476
rect 34572 35436 34578 35448
rect 34701 35445 34713 35448
rect 34747 35445 34759 35479
rect 36464 35476 36492 35643
rect 38470 35640 38476 35652
rect 38528 35680 38534 35692
rect 38565 35683 38623 35689
rect 38565 35680 38577 35683
rect 38528 35652 38577 35680
rect 38528 35640 38534 35652
rect 38565 35649 38577 35652
rect 38611 35649 38623 35683
rect 38565 35643 38623 35649
rect 38746 35640 38752 35692
rect 38804 35680 38810 35692
rect 38841 35683 38899 35689
rect 38841 35680 38853 35683
rect 38804 35652 38853 35680
rect 38804 35640 38810 35652
rect 38841 35649 38853 35652
rect 38887 35649 38899 35683
rect 39132 35680 39160 35788
rect 39298 35776 39304 35788
rect 39356 35776 39362 35828
rect 40034 35776 40040 35828
rect 40092 35816 40098 35828
rect 40681 35819 40739 35825
rect 40681 35816 40693 35819
rect 40092 35788 40693 35816
rect 40092 35776 40098 35788
rect 40681 35785 40693 35788
rect 40727 35816 40739 35819
rect 40862 35816 40868 35828
rect 40727 35788 40868 35816
rect 40727 35785 40739 35788
rect 40681 35779 40739 35785
rect 40862 35776 40868 35788
rect 40920 35776 40926 35828
rect 41690 35816 41696 35828
rect 41616 35788 41696 35816
rect 39485 35751 39543 35757
rect 39485 35717 39497 35751
rect 39531 35748 39543 35751
rect 40313 35751 40371 35757
rect 40313 35748 40325 35751
rect 39531 35720 40325 35748
rect 39531 35717 39543 35720
rect 39485 35711 39543 35717
rect 40313 35717 40325 35720
rect 40359 35717 40371 35751
rect 40313 35711 40371 35717
rect 40494 35680 40500 35692
rect 39132 35652 39620 35680
rect 40455 35652 40500 35680
rect 38841 35643 38899 35649
rect 37277 35615 37335 35621
rect 37277 35581 37289 35615
rect 37323 35612 37335 35615
rect 37458 35612 37464 35624
rect 37323 35584 37464 35612
rect 37323 35581 37335 35584
rect 37277 35575 37335 35581
rect 37458 35572 37464 35584
rect 37516 35572 37522 35624
rect 36722 35544 36728 35556
rect 36683 35516 36728 35544
rect 36722 35504 36728 35516
rect 36780 35504 36786 35556
rect 37461 35479 37519 35485
rect 37461 35476 37473 35479
rect 36464 35448 37473 35476
rect 34701 35439 34759 35445
rect 37461 35445 37473 35448
rect 37507 35476 37519 35479
rect 37642 35476 37648 35488
rect 37507 35448 37648 35476
rect 37507 35445 37519 35448
rect 37461 35439 37519 35445
rect 37642 35436 37648 35448
rect 37700 35436 37706 35488
rect 39390 35436 39396 35488
rect 39448 35476 39454 35488
rect 39485 35479 39543 35485
rect 39485 35476 39497 35479
rect 39448 35448 39497 35476
rect 39448 35436 39454 35448
rect 39485 35445 39497 35448
rect 39531 35445 39543 35479
rect 39592 35476 39620 35652
rect 40494 35640 40500 35652
rect 40552 35640 40558 35692
rect 41616 35689 41644 35788
rect 41690 35776 41696 35788
rect 41748 35776 41754 35828
rect 41877 35819 41935 35825
rect 41877 35785 41889 35819
rect 41923 35816 41935 35819
rect 42058 35816 42064 35828
rect 41923 35788 42064 35816
rect 41923 35785 41935 35788
rect 41877 35779 41935 35785
rect 42058 35776 42064 35788
rect 42116 35776 42122 35828
rect 43349 35819 43407 35825
rect 43349 35785 43361 35819
rect 43395 35816 43407 35819
rect 43990 35816 43996 35828
rect 43395 35788 43996 35816
rect 43395 35785 43407 35788
rect 43349 35779 43407 35785
rect 43990 35776 43996 35788
rect 44048 35776 44054 35828
rect 40773 35683 40831 35689
rect 40773 35649 40785 35683
rect 40819 35649 40831 35683
rect 40773 35643 40831 35649
rect 41601 35683 41659 35689
rect 41601 35649 41613 35683
rect 41647 35649 41659 35683
rect 41601 35643 41659 35649
rect 41693 35683 41751 35689
rect 41693 35649 41705 35683
rect 41739 35680 41751 35683
rect 41966 35680 41972 35692
rect 41739 35652 41972 35680
rect 41739 35649 41751 35652
rect 41693 35643 41751 35649
rect 39758 35572 39764 35624
rect 39816 35612 39822 35624
rect 40788 35612 40816 35643
rect 39816 35584 40816 35612
rect 39816 35572 39822 35584
rect 39666 35504 39672 35556
rect 39724 35544 39730 35556
rect 39853 35547 39911 35553
rect 39853 35544 39865 35547
rect 39724 35516 39865 35544
rect 39724 35504 39730 35516
rect 39853 35513 39865 35516
rect 39899 35544 39911 35547
rect 41708 35544 41736 35643
rect 41966 35640 41972 35652
rect 42024 35640 42030 35692
rect 43254 35680 43260 35692
rect 43215 35652 43260 35680
rect 43254 35640 43260 35652
rect 43312 35640 43318 35692
rect 39899 35516 41736 35544
rect 39899 35513 39911 35516
rect 39853 35507 39911 35513
rect 43254 35476 43260 35488
rect 39592 35448 43260 35476
rect 39485 35439 39543 35445
rect 43254 35436 43260 35448
rect 43312 35436 43318 35488
rect 44085 35479 44143 35485
rect 44085 35445 44097 35479
rect 44131 35476 44143 35479
rect 44174 35476 44180 35488
rect 44131 35448 44180 35476
rect 44131 35445 44143 35448
rect 44085 35439 44143 35445
rect 44174 35436 44180 35448
rect 44232 35436 44238 35488
rect 1104 35386 44896 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 44896 35386
rect 1104 35312 44896 35334
rect 22189 35275 22247 35281
rect 22189 35241 22201 35275
rect 22235 35272 22247 35275
rect 22278 35272 22284 35284
rect 22235 35244 22284 35272
rect 22235 35241 22247 35244
rect 22189 35235 22247 35241
rect 22278 35232 22284 35244
rect 22336 35272 22342 35284
rect 22646 35272 22652 35284
rect 22336 35244 22652 35272
rect 22336 35232 22342 35244
rect 22646 35232 22652 35244
rect 22704 35232 22710 35284
rect 22830 35232 22836 35284
rect 22888 35272 22894 35284
rect 22925 35275 22983 35281
rect 22925 35272 22937 35275
rect 22888 35244 22937 35272
rect 22888 35232 22894 35244
rect 22925 35241 22937 35244
rect 22971 35241 22983 35275
rect 22925 35235 22983 35241
rect 23109 35275 23167 35281
rect 23109 35241 23121 35275
rect 23155 35272 23167 35275
rect 23474 35272 23480 35284
rect 23155 35244 23480 35272
rect 23155 35241 23167 35244
rect 23109 35235 23167 35241
rect 23474 35232 23480 35244
rect 23532 35232 23538 35284
rect 23658 35272 23664 35284
rect 23619 35244 23664 35272
rect 23658 35232 23664 35244
rect 23716 35232 23722 35284
rect 27801 35275 27859 35281
rect 27801 35241 27813 35275
rect 27847 35272 27859 35275
rect 28074 35272 28080 35284
rect 27847 35244 28080 35272
rect 27847 35241 27859 35244
rect 27801 35235 27859 35241
rect 28074 35232 28080 35244
rect 28132 35272 28138 35284
rect 28442 35272 28448 35284
rect 28132 35244 28448 35272
rect 28132 35232 28138 35244
rect 28442 35232 28448 35244
rect 28500 35232 28506 35284
rect 28721 35275 28779 35281
rect 28721 35241 28733 35275
rect 28767 35272 28779 35275
rect 29178 35272 29184 35284
rect 28767 35244 29184 35272
rect 28767 35241 28779 35244
rect 28721 35235 28779 35241
rect 29178 35232 29184 35244
rect 29236 35232 29242 35284
rect 34054 35272 34060 35284
rect 34015 35244 34060 35272
rect 34054 35232 34060 35244
rect 34112 35232 34118 35284
rect 34422 35232 34428 35284
rect 34480 35272 34486 35284
rect 35986 35272 35992 35284
rect 34480 35244 35894 35272
rect 35947 35244 35992 35272
rect 34480 35232 34486 35244
rect 26418 35164 26424 35216
rect 26476 35204 26482 35216
rect 27985 35207 28043 35213
rect 27985 35204 27997 35207
rect 26476 35176 27997 35204
rect 26476 35164 26482 35176
rect 22738 35136 22744 35148
rect 22112 35108 22744 35136
rect 19978 35068 19984 35080
rect 19939 35040 19984 35068
rect 19978 35028 19984 35040
rect 20036 35028 20042 35080
rect 22112 35077 22140 35108
rect 22738 35096 22744 35108
rect 22796 35096 22802 35148
rect 23014 35096 23020 35148
rect 23072 35136 23078 35148
rect 23072 35108 26188 35136
rect 23072 35096 23078 35108
rect 22097 35071 22155 35077
rect 22097 35037 22109 35071
rect 22143 35037 22155 35071
rect 22097 35031 22155 35037
rect 22646 35028 22652 35080
rect 22704 35068 22710 35080
rect 24765 35071 24823 35077
rect 22704 35040 24716 35068
rect 22704 35028 22710 35040
rect 17218 35000 17224 35012
rect 17179 34972 17224 35000
rect 17218 34960 17224 34972
rect 17276 34960 17282 35012
rect 17402 35000 17408 35012
rect 17363 34972 17408 35000
rect 17402 34960 17408 34972
rect 17460 34960 17466 35012
rect 22741 35003 22799 35009
rect 22741 34969 22753 35003
rect 22787 35000 22799 35003
rect 23106 35000 23112 35012
rect 22787 34972 23112 35000
rect 22787 34969 22799 34972
rect 22741 34963 22799 34969
rect 23106 34960 23112 34972
rect 23164 34960 23170 35012
rect 23753 35003 23811 35009
rect 23753 34969 23765 35003
rect 23799 35000 23811 35003
rect 24486 35000 24492 35012
rect 23799 34972 24492 35000
rect 23799 34969 23811 34972
rect 23753 34963 23811 34969
rect 24486 34960 24492 34972
rect 24544 34960 24550 35012
rect 24688 35000 24716 35040
rect 24765 35037 24777 35071
rect 24811 35068 24823 35071
rect 24854 35068 24860 35080
rect 24811 35040 24860 35068
rect 24811 35037 24823 35040
rect 24765 35031 24823 35037
rect 24854 35028 24860 35040
rect 24912 35028 24918 35080
rect 25590 35068 25596 35080
rect 25551 35040 25596 35068
rect 25590 35028 25596 35040
rect 25648 35028 25654 35080
rect 25958 35068 25964 35080
rect 25919 35040 25964 35068
rect 25958 35028 25964 35040
rect 26016 35028 26022 35080
rect 25130 35000 25136 35012
rect 24688 34972 25136 35000
rect 25130 34960 25136 34972
rect 25188 34960 25194 35012
rect 26160 34944 26188 35108
rect 26528 35077 26556 35176
rect 27985 35173 27997 35176
rect 28031 35173 28043 35207
rect 29549 35207 29607 35213
rect 29549 35204 29561 35207
rect 27985 35167 28043 35173
rect 28966 35176 29561 35204
rect 28966 35148 28994 35176
rect 29549 35173 29561 35176
rect 29595 35173 29607 35207
rect 33226 35204 33232 35216
rect 29549 35167 29607 35173
rect 32324 35176 33232 35204
rect 26786 35136 26792 35148
rect 26747 35108 26792 35136
rect 26786 35096 26792 35108
rect 26844 35096 26850 35148
rect 27706 35136 27712 35148
rect 27667 35108 27712 35136
rect 27706 35096 27712 35108
rect 27764 35136 27770 35148
rect 28902 35136 28908 35148
rect 27764 35108 28908 35136
rect 27764 35096 27770 35108
rect 28902 35096 28908 35108
rect 28960 35108 28994 35148
rect 30926 35136 30932 35148
rect 30887 35108 30932 35136
rect 28960 35096 28966 35108
rect 30926 35096 30932 35108
rect 30984 35096 30990 35148
rect 32324 35145 32352 35176
rect 33226 35164 33232 35176
rect 33284 35204 33290 35216
rect 33505 35207 33563 35213
rect 33505 35204 33517 35207
rect 33284 35176 33517 35204
rect 33284 35164 33290 35176
rect 33505 35173 33517 35176
rect 33551 35173 33563 35207
rect 35342 35204 35348 35216
rect 35303 35176 35348 35204
rect 33505 35167 33563 35173
rect 35342 35164 35348 35176
rect 35400 35164 35406 35216
rect 35866 35204 35894 35244
rect 35986 35232 35992 35244
rect 36044 35232 36050 35284
rect 39850 35272 39856 35284
rect 37844 35244 39856 35272
rect 37844 35204 37872 35244
rect 39850 35232 39856 35244
rect 39908 35232 39914 35284
rect 41690 35232 41696 35284
rect 41748 35272 41754 35284
rect 41877 35275 41935 35281
rect 41877 35272 41889 35275
rect 41748 35244 41889 35272
rect 41748 35232 41754 35244
rect 41877 35241 41889 35244
rect 41923 35241 41935 35275
rect 41877 35235 41935 35241
rect 38470 35204 38476 35216
rect 35866 35176 37872 35204
rect 38431 35176 38476 35204
rect 38470 35164 38476 35176
rect 38528 35164 38534 35216
rect 39025 35207 39083 35213
rect 39025 35173 39037 35207
rect 39071 35204 39083 35207
rect 39666 35204 39672 35216
rect 39071 35176 39672 35204
rect 39071 35173 39083 35176
rect 39025 35167 39083 35173
rect 39666 35164 39672 35176
rect 39724 35164 39730 35216
rect 32309 35139 32367 35145
rect 32309 35105 32321 35139
rect 32355 35105 32367 35139
rect 32309 35099 32367 35105
rect 32766 35096 32772 35148
rect 32824 35136 32830 35148
rect 36078 35136 36084 35148
rect 32824 35108 36084 35136
rect 32824 35096 32830 35108
rect 36078 35096 36084 35108
rect 36136 35096 36142 35148
rect 38654 35096 38660 35148
rect 38712 35136 38718 35148
rect 39942 35136 39948 35148
rect 38712 35108 39948 35136
rect 38712 35096 38718 35108
rect 39942 35096 39948 35108
rect 40000 35136 40006 35148
rect 40497 35139 40555 35145
rect 40497 35136 40509 35139
rect 40000 35108 40509 35136
rect 40000 35096 40006 35108
rect 40497 35105 40509 35108
rect 40543 35105 40555 35139
rect 42702 35136 42708 35148
rect 42663 35108 42708 35136
rect 40497 35099 40555 35105
rect 42702 35096 42708 35108
rect 42760 35096 42766 35148
rect 44174 35136 44180 35148
rect 44135 35108 44180 35136
rect 44174 35096 44180 35108
rect 44232 35096 44238 35148
rect 26513 35071 26571 35077
rect 26513 35037 26525 35071
rect 26559 35037 26571 35071
rect 26513 35031 26571 35037
rect 26697 35071 26755 35077
rect 26697 35037 26709 35071
rect 26743 35068 26755 35071
rect 27614 35068 27620 35080
rect 26743 35040 27620 35068
rect 26743 35037 26755 35040
rect 26697 35031 26755 35037
rect 27614 35028 27620 35040
rect 27672 35028 27678 35080
rect 27801 35071 27859 35077
rect 27801 35037 27813 35071
rect 27847 35068 27859 35071
rect 28258 35068 28264 35080
rect 27847 35040 28264 35068
rect 27847 35037 27859 35040
rect 27801 35031 27859 35037
rect 28258 35028 28264 35040
rect 28316 35028 28322 35080
rect 29822 35068 29828 35080
rect 28552 35040 29828 35068
rect 26878 34960 26884 35012
rect 26936 35000 26942 35012
rect 28552 35009 28580 35040
rect 29822 35028 29828 35040
rect 29880 35028 29886 35080
rect 32490 35068 32496 35080
rect 32451 35040 32496 35068
rect 32490 35028 32496 35040
rect 32548 35028 32554 35080
rect 32585 35071 32643 35077
rect 32585 35037 32597 35071
rect 32631 35068 32643 35071
rect 33134 35068 33140 35080
rect 32631 35040 33140 35068
rect 32631 35037 32643 35040
rect 32585 35031 32643 35037
rect 33134 35028 33140 35040
rect 33192 35068 33198 35080
rect 33965 35071 34023 35077
rect 33965 35068 33977 35071
rect 33192 35040 33977 35068
rect 33192 35028 33198 35040
rect 33965 35037 33977 35040
rect 34011 35037 34023 35071
rect 33965 35031 34023 35037
rect 34149 35071 34207 35077
rect 34149 35037 34161 35071
rect 34195 35068 34207 35071
rect 34238 35068 34244 35080
rect 34195 35040 34244 35068
rect 34195 35037 34207 35040
rect 34149 35031 34207 35037
rect 34238 35028 34244 35040
rect 34296 35028 34302 35080
rect 40764 35071 40822 35077
rect 40764 35037 40776 35071
rect 40810 35068 40822 35071
rect 41598 35068 41604 35080
rect 40810 35040 41604 35068
rect 40810 35037 40822 35040
rect 40764 35031 40822 35037
rect 41598 35028 41604 35040
rect 41656 35028 41662 35080
rect 27525 35003 27583 35009
rect 27525 35000 27537 35003
rect 26936 34972 27537 35000
rect 26936 34960 26942 34972
rect 27525 34969 27537 34972
rect 27571 34969 27583 35003
rect 27525 34963 27583 34969
rect 28537 35003 28595 35009
rect 28537 34969 28549 35003
rect 28583 34969 28595 35003
rect 28537 34963 28595 34969
rect 28753 35003 28811 35009
rect 28753 34969 28765 35003
rect 28799 35000 28811 35003
rect 29638 35000 29644 35012
rect 28799 34972 29644 35000
rect 28799 34969 28811 34972
rect 28753 34963 28811 34969
rect 17586 34932 17592 34944
rect 17547 34904 17592 34932
rect 17586 34892 17592 34904
rect 17644 34892 17650 34944
rect 19426 34892 19432 34944
rect 19484 34932 19490 34944
rect 19797 34935 19855 34941
rect 19797 34932 19809 34935
rect 19484 34904 19809 34932
rect 19484 34892 19490 34904
rect 19797 34901 19809 34904
rect 19843 34901 19855 34935
rect 19797 34895 19855 34901
rect 22951 34935 23009 34941
rect 22951 34901 22963 34935
rect 22997 34932 23009 34935
rect 23842 34932 23848 34944
rect 22997 34904 23848 34932
rect 22997 34901 23009 34904
rect 22951 34895 23009 34901
rect 23842 34892 23848 34904
rect 23900 34892 23906 34944
rect 24946 34932 24952 34944
rect 24907 34904 24952 34932
rect 24946 34892 24952 34904
rect 25004 34892 25010 34944
rect 26142 34892 26148 34944
rect 26200 34932 26206 34944
rect 28552 34932 28580 34963
rect 29638 34960 29644 34972
rect 29696 34960 29702 35012
rect 30374 34960 30380 35012
rect 30432 35000 30438 35012
rect 30662 35003 30720 35009
rect 30662 35000 30674 35003
rect 30432 34972 30674 35000
rect 30432 34960 30438 34972
rect 30662 34969 30674 34972
rect 30708 34969 30720 35003
rect 33318 35000 33324 35012
rect 33279 34972 33324 35000
rect 30662 34963 30720 34969
rect 33318 34960 33324 34972
rect 33376 35000 33382 35012
rect 35161 35003 35219 35009
rect 35161 35000 35173 35003
rect 33376 34972 35173 35000
rect 33376 34960 33382 34972
rect 35161 34969 35173 34972
rect 35207 34969 35219 35003
rect 35161 34963 35219 34969
rect 35894 34960 35900 35012
rect 35952 35000 35958 35012
rect 35952 34972 35997 35000
rect 35952 34960 35958 34972
rect 38562 34960 38568 35012
rect 38620 35000 38626 35012
rect 38749 35003 38807 35009
rect 38749 35000 38761 35003
rect 38620 34972 38761 35000
rect 38620 34960 38626 34972
rect 38749 34969 38761 34972
rect 38795 34969 38807 35003
rect 38749 34963 38807 34969
rect 38841 35003 38899 35009
rect 38841 34969 38853 35003
rect 38887 35000 38899 35003
rect 40678 35000 40684 35012
rect 38887 34972 40684 35000
rect 38887 34969 38899 34972
rect 38841 34963 38899 34969
rect 40678 34960 40684 34972
rect 40736 34960 40742 35012
rect 43622 34960 43628 35012
rect 43680 35000 43686 35012
rect 43993 35003 44051 35009
rect 43993 35000 44005 35003
rect 43680 34972 44005 35000
rect 43680 34960 43686 34972
rect 43993 34969 44005 34972
rect 44039 34969 44051 35003
rect 43993 34963 44051 34969
rect 26200 34904 28580 34932
rect 28905 34935 28963 34941
rect 26200 34892 26206 34904
rect 28905 34901 28917 34935
rect 28951 34932 28963 34935
rect 29454 34932 29460 34944
rect 28951 34904 29460 34932
rect 28951 34901 28963 34904
rect 28905 34895 28963 34901
rect 29454 34892 29460 34904
rect 29512 34892 29518 34944
rect 32306 34932 32312 34944
rect 32267 34904 32312 34932
rect 32306 34892 32312 34904
rect 32364 34892 32370 34944
rect 38657 34935 38715 34941
rect 38657 34901 38669 34935
rect 38703 34932 38715 34935
rect 38930 34932 38936 34944
rect 38703 34904 38936 34932
rect 38703 34901 38715 34904
rect 38657 34895 38715 34901
rect 38930 34892 38936 34904
rect 38988 34892 38994 34944
rect 1104 34842 44896 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 44896 34842
rect 1104 34768 44896 34790
rect 16117 34731 16175 34737
rect 16117 34697 16129 34731
rect 16163 34697 16175 34731
rect 16117 34691 16175 34697
rect 16132 34660 16160 34691
rect 17402 34688 17408 34740
rect 17460 34728 17466 34740
rect 18049 34731 18107 34737
rect 18049 34728 18061 34731
rect 17460 34700 18061 34728
rect 17460 34688 17466 34700
rect 18049 34697 18061 34700
rect 18095 34697 18107 34731
rect 18049 34691 18107 34697
rect 19889 34731 19947 34737
rect 19889 34697 19901 34731
rect 19935 34728 19947 34731
rect 19978 34728 19984 34740
rect 19935 34700 19984 34728
rect 19935 34697 19947 34700
rect 19889 34691 19947 34697
rect 19978 34688 19984 34700
rect 20036 34688 20042 34740
rect 22646 34728 22652 34740
rect 20088 34700 22652 34728
rect 16914 34663 16972 34669
rect 16914 34660 16926 34663
rect 16132 34632 16926 34660
rect 16914 34629 16926 34632
rect 16960 34629 16972 34663
rect 20088 34660 20116 34700
rect 22646 34688 22652 34700
rect 22704 34688 22710 34740
rect 22830 34728 22836 34740
rect 22791 34700 22836 34728
rect 22830 34688 22836 34700
rect 22888 34688 22894 34740
rect 23014 34688 23020 34740
rect 23072 34728 23078 34740
rect 23842 34728 23848 34740
rect 23072 34700 23244 34728
rect 23803 34700 23848 34728
rect 23072 34688 23078 34700
rect 16914 34623 16972 34629
rect 19536 34632 20116 34660
rect 15933 34595 15991 34601
rect 15933 34561 15945 34595
rect 15979 34592 15991 34595
rect 18509 34595 18567 34601
rect 18509 34592 18521 34595
rect 15979 34564 18521 34592
rect 15979 34561 15991 34564
rect 15933 34555 15991 34561
rect 18509 34561 18521 34564
rect 18555 34561 18567 34595
rect 18690 34592 18696 34604
rect 18651 34564 18696 34592
rect 18509 34555 18567 34561
rect 18690 34552 18696 34564
rect 18748 34552 18754 34604
rect 19536 34601 19564 34632
rect 20714 34620 20720 34672
rect 20772 34660 20778 34672
rect 21085 34663 21143 34669
rect 21085 34660 21097 34663
rect 20772 34632 21097 34660
rect 20772 34620 20778 34632
rect 21085 34629 21097 34632
rect 21131 34629 21143 34663
rect 21266 34660 21272 34672
rect 21227 34632 21272 34660
rect 21085 34623 21143 34629
rect 21266 34620 21272 34632
rect 21324 34620 21330 34672
rect 22186 34660 22192 34672
rect 22147 34632 22192 34660
rect 22186 34620 22192 34632
rect 22244 34620 22250 34672
rect 22738 34620 22744 34672
rect 22796 34660 22802 34672
rect 23109 34663 23167 34669
rect 23109 34660 23121 34663
rect 22796 34632 23121 34660
rect 22796 34620 22802 34632
rect 23109 34629 23121 34632
rect 23155 34629 23167 34663
rect 23216 34660 23244 34700
rect 23842 34688 23848 34700
rect 23900 34688 23906 34740
rect 25866 34688 25872 34740
rect 25924 34728 25930 34740
rect 26053 34731 26111 34737
rect 26053 34728 26065 34731
rect 25924 34700 26065 34728
rect 25924 34688 25930 34700
rect 26053 34697 26065 34700
rect 26099 34728 26111 34731
rect 27154 34728 27160 34740
rect 26099 34700 27160 34728
rect 26099 34697 26111 34700
rect 26053 34691 26111 34697
rect 27154 34688 27160 34700
rect 27212 34688 27218 34740
rect 27614 34688 27620 34740
rect 27672 34728 27678 34740
rect 29178 34728 29184 34740
rect 27672 34700 29040 34728
rect 29139 34700 29184 34728
rect 27672 34688 27678 34700
rect 24946 34669 24952 34672
rect 24940 34660 24952 34669
rect 23216 34632 24808 34660
rect 24907 34632 24952 34660
rect 23109 34623 23167 34629
rect 18877 34595 18935 34601
rect 18877 34561 18889 34595
rect 18923 34592 18935 34595
rect 19521 34595 19579 34601
rect 19521 34592 19533 34595
rect 18923 34564 19533 34592
rect 18923 34561 18935 34564
rect 18877 34555 18935 34561
rect 19521 34561 19533 34564
rect 19567 34561 19579 34595
rect 19702 34592 19708 34604
rect 19663 34564 19708 34592
rect 19521 34555 19579 34561
rect 19702 34552 19708 34564
rect 19760 34552 19766 34604
rect 22830 34552 22836 34604
rect 22888 34592 22894 34604
rect 23014 34592 23020 34604
rect 22888 34564 23020 34592
rect 22888 34552 22894 34564
rect 23014 34552 23020 34564
rect 23072 34552 23078 34604
rect 23198 34552 23204 34604
rect 23256 34592 23262 34604
rect 23382 34592 23388 34604
rect 23256 34564 23301 34592
rect 23343 34564 23388 34592
rect 23256 34552 23262 34564
rect 23382 34552 23388 34564
rect 23440 34552 23446 34604
rect 23845 34595 23903 34601
rect 23845 34561 23857 34595
rect 23891 34561 23903 34595
rect 24026 34592 24032 34604
rect 23987 34564 24032 34592
rect 23845 34555 23903 34561
rect 15378 34484 15384 34536
rect 15436 34524 15442 34536
rect 15838 34524 15844 34536
rect 15436 34496 15844 34524
rect 15436 34484 15442 34496
rect 15838 34484 15844 34496
rect 15896 34524 15902 34536
rect 16669 34527 16727 34533
rect 16669 34524 16681 34527
rect 15896 34496 16681 34524
rect 15896 34484 15902 34496
rect 16669 34493 16681 34496
rect 16715 34493 16727 34527
rect 16669 34487 16727 34493
rect 22373 34527 22431 34533
rect 22373 34493 22385 34527
rect 22419 34524 22431 34527
rect 23216 34524 23244 34552
rect 23860 34524 23888 34555
rect 24026 34552 24032 34564
rect 24084 34552 24090 34604
rect 24302 34552 24308 34604
rect 24360 34592 24366 34604
rect 24673 34595 24731 34601
rect 24673 34592 24685 34595
rect 24360 34564 24685 34592
rect 24360 34552 24366 34564
rect 24673 34561 24685 34564
rect 24719 34561 24731 34595
rect 24780 34592 24808 34632
rect 24940 34623 24952 34632
rect 24946 34620 24952 34623
rect 25004 34620 25010 34672
rect 28902 34660 28908 34672
rect 28000 34632 28764 34660
rect 28863 34632 28908 34660
rect 28000 34604 28028 34632
rect 25774 34592 25780 34604
rect 24780 34564 25780 34592
rect 24673 34555 24731 34561
rect 25774 34552 25780 34564
rect 25832 34552 25838 34604
rect 27341 34595 27399 34601
rect 27341 34561 27353 34595
rect 27387 34592 27399 34595
rect 27430 34592 27436 34604
rect 27387 34564 27436 34592
rect 27387 34561 27399 34564
rect 27341 34555 27399 34561
rect 27430 34552 27436 34564
rect 27488 34552 27494 34604
rect 27617 34595 27675 34601
rect 27617 34561 27629 34595
rect 27663 34592 27675 34595
rect 27982 34592 27988 34604
rect 27663 34564 27988 34592
rect 27663 34561 27675 34564
rect 27617 34555 27675 34561
rect 27982 34552 27988 34564
rect 28040 34552 28046 34604
rect 28626 34592 28632 34604
rect 28587 34564 28632 34592
rect 28626 34552 28632 34564
rect 28684 34552 28690 34604
rect 28736 34592 28764 34632
rect 28902 34620 28908 34632
rect 28960 34620 28966 34672
rect 29012 34660 29040 34700
rect 29178 34688 29184 34700
rect 29236 34688 29242 34740
rect 29638 34728 29644 34740
rect 29599 34700 29644 34728
rect 29638 34688 29644 34700
rect 29696 34688 29702 34740
rect 30745 34731 30803 34737
rect 30745 34697 30757 34731
rect 30791 34728 30803 34731
rect 31386 34728 31392 34740
rect 30791 34700 31392 34728
rect 30791 34697 30803 34700
rect 30745 34691 30803 34697
rect 31386 34688 31392 34700
rect 31444 34688 31450 34740
rect 32582 34688 32588 34740
rect 32640 34728 32646 34740
rect 32877 34731 32935 34737
rect 32877 34728 32889 34731
rect 32640 34700 32889 34728
rect 32640 34688 32646 34700
rect 32877 34697 32889 34700
rect 32923 34728 32935 34731
rect 33042 34728 33048 34740
rect 32923 34700 33048 34728
rect 32923 34697 32935 34700
rect 32877 34691 32935 34697
rect 33042 34688 33048 34700
rect 33100 34688 33106 34740
rect 38194 34688 38200 34740
rect 38252 34728 38258 34740
rect 38470 34728 38476 34740
rect 38252 34700 38476 34728
rect 38252 34688 38258 34700
rect 38470 34688 38476 34700
rect 38528 34728 38534 34740
rect 38749 34731 38807 34737
rect 38749 34728 38761 34731
rect 38528 34700 38761 34728
rect 38528 34688 38534 34700
rect 38749 34697 38761 34700
rect 38795 34697 38807 34731
rect 38749 34691 38807 34697
rect 41233 34731 41291 34737
rect 41233 34697 41245 34731
rect 41279 34728 41291 34731
rect 41506 34728 41512 34740
rect 41279 34700 41512 34728
rect 41279 34697 41291 34700
rect 41233 34691 41291 34697
rect 41506 34688 41512 34700
rect 41564 34688 41570 34740
rect 43622 34728 43628 34740
rect 43583 34700 43628 34728
rect 43622 34688 43628 34700
rect 43680 34688 43686 34740
rect 32677 34663 32735 34669
rect 29012 34632 30604 34660
rect 28813 34595 28871 34601
rect 28813 34592 28825 34595
rect 28736 34564 28825 34592
rect 28813 34561 28825 34564
rect 28859 34561 28871 34595
rect 28813 34555 28871 34561
rect 28994 34552 29000 34604
rect 29052 34592 29058 34604
rect 29638 34592 29644 34604
rect 29052 34564 29097 34592
rect 29599 34564 29644 34592
rect 29052 34552 29058 34564
rect 29638 34552 29644 34564
rect 29696 34552 29702 34604
rect 29825 34595 29883 34601
rect 29825 34561 29837 34595
rect 29871 34561 29883 34595
rect 30466 34592 30472 34604
rect 30427 34564 30472 34592
rect 29825 34555 29883 34561
rect 29840 34524 29868 34555
rect 30466 34552 30472 34564
rect 30524 34552 30530 34604
rect 30576 34601 30604 34632
rect 32677 34629 32689 34663
rect 32723 34660 32735 34663
rect 32766 34660 32772 34672
rect 32723 34632 32772 34660
rect 32723 34629 32735 34632
rect 32677 34623 32735 34629
rect 32766 34620 32772 34632
rect 32824 34620 32830 34672
rect 30561 34595 30619 34601
rect 30561 34561 30573 34595
rect 30607 34592 30619 34595
rect 34514 34592 34520 34604
rect 30607 34564 34520 34592
rect 30607 34561 30619 34564
rect 30561 34555 30619 34561
rect 34514 34552 34520 34564
rect 34572 34552 34578 34604
rect 37366 34592 37372 34604
rect 37279 34564 37372 34592
rect 37366 34552 37372 34564
rect 37424 34592 37430 34604
rect 38562 34592 38568 34604
rect 37424 34564 38568 34592
rect 37424 34552 37430 34564
rect 38562 34552 38568 34564
rect 38620 34552 38626 34604
rect 38657 34595 38715 34601
rect 38657 34561 38669 34595
rect 38703 34561 38715 34595
rect 38930 34592 38936 34604
rect 38891 34564 38936 34592
rect 38657 34555 38715 34561
rect 37642 34524 37648 34536
rect 22419 34496 23244 34524
rect 23400 34496 23888 34524
rect 27724 34496 29868 34524
rect 37603 34496 37648 34524
rect 22419 34493 22431 34496
rect 22373 34487 22431 34493
rect 22278 34416 22284 34468
rect 22336 34456 22342 34468
rect 23400 34456 23428 34496
rect 22336 34428 23428 34456
rect 22336 34416 22342 34428
rect 27522 34416 27528 34468
rect 27580 34456 27586 34468
rect 27724 34456 27752 34496
rect 37642 34484 37648 34496
rect 37700 34524 37706 34536
rect 38378 34524 38384 34536
rect 37700 34496 38384 34524
rect 37700 34484 37706 34496
rect 38378 34484 38384 34496
rect 38436 34524 38442 34536
rect 38672 34524 38700 34555
rect 38930 34552 38936 34564
rect 38988 34552 38994 34604
rect 39758 34552 39764 34604
rect 39816 34592 39822 34604
rect 39945 34595 40003 34601
rect 39945 34592 39957 34595
rect 39816 34564 39957 34592
rect 39816 34552 39822 34564
rect 39945 34561 39957 34564
rect 39991 34561 40003 34595
rect 40126 34592 40132 34604
rect 40087 34564 40132 34592
rect 39945 34555 40003 34561
rect 40126 34552 40132 34564
rect 40184 34552 40190 34604
rect 41509 34595 41567 34601
rect 41509 34561 41521 34595
rect 41555 34592 41567 34595
rect 41690 34592 41696 34604
rect 41555 34564 41696 34592
rect 41555 34561 41567 34564
rect 41509 34555 41567 34561
rect 41690 34552 41696 34564
rect 41748 34552 41754 34604
rect 43533 34595 43591 34601
rect 43533 34561 43545 34595
rect 43579 34592 43591 34595
rect 43622 34592 43628 34604
rect 43579 34564 43628 34592
rect 43579 34561 43591 34564
rect 43533 34555 43591 34561
rect 43622 34552 43628 34564
rect 43680 34552 43686 34604
rect 38436 34496 38700 34524
rect 39853 34527 39911 34533
rect 38436 34484 38442 34496
rect 39853 34493 39865 34527
rect 39899 34524 39911 34527
rect 40034 34524 40040 34536
rect 39899 34496 40040 34524
rect 39899 34493 39911 34496
rect 39853 34487 39911 34493
rect 40034 34484 40040 34496
rect 40092 34484 40098 34536
rect 41230 34524 41236 34536
rect 41191 34496 41236 34524
rect 41230 34484 41236 34496
rect 41288 34484 41294 34536
rect 33134 34456 33140 34468
rect 27580 34428 27752 34456
rect 32876 34428 33140 34456
rect 27580 34416 27586 34428
rect 20901 34391 20959 34397
rect 20901 34357 20913 34391
rect 20947 34388 20959 34391
rect 20990 34388 20996 34400
rect 20947 34360 20996 34388
rect 20947 34357 20959 34360
rect 20901 34351 20959 34357
rect 20990 34348 20996 34360
rect 21048 34348 21054 34400
rect 32876 34397 32904 34428
rect 33134 34416 33140 34428
rect 33192 34416 33198 34468
rect 41417 34459 41475 34465
rect 41417 34425 41429 34459
rect 41463 34456 41475 34459
rect 41966 34456 41972 34468
rect 41463 34428 41972 34456
rect 41463 34425 41475 34428
rect 41417 34419 41475 34425
rect 41966 34416 41972 34428
rect 42024 34416 42030 34468
rect 32861 34391 32919 34397
rect 32861 34357 32873 34391
rect 32907 34357 32919 34391
rect 33042 34388 33048 34400
rect 33003 34360 33048 34388
rect 32861 34351 32919 34357
rect 33042 34348 33048 34360
rect 33100 34348 33106 34400
rect 38746 34348 38752 34400
rect 38804 34388 38810 34400
rect 39117 34391 39175 34397
rect 39117 34388 39129 34391
rect 38804 34360 39129 34388
rect 38804 34348 38810 34360
rect 39117 34357 39129 34360
rect 39163 34357 39175 34391
rect 39117 34351 39175 34357
rect 40218 34348 40224 34400
rect 40276 34388 40282 34400
rect 40313 34391 40371 34397
rect 40313 34388 40325 34391
rect 40276 34360 40325 34388
rect 40276 34348 40282 34360
rect 40313 34357 40325 34360
rect 40359 34357 40371 34391
rect 40313 34351 40371 34357
rect 42334 34348 42340 34400
rect 42392 34388 42398 34400
rect 42889 34391 42947 34397
rect 42889 34388 42901 34391
rect 42392 34360 42901 34388
rect 42392 34348 42398 34360
rect 42889 34357 42901 34360
rect 42935 34357 42947 34391
rect 42889 34351 42947 34357
rect 1104 34298 44896 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 44896 34298
rect 1104 34224 44896 34246
rect 16761 34187 16819 34193
rect 16761 34153 16773 34187
rect 16807 34184 16819 34187
rect 16942 34184 16948 34196
rect 16807 34156 16948 34184
rect 16807 34153 16819 34156
rect 16761 34147 16819 34153
rect 16942 34144 16948 34156
rect 17000 34184 17006 34196
rect 17218 34184 17224 34196
rect 17000 34156 17224 34184
rect 17000 34144 17006 34156
rect 17218 34144 17224 34156
rect 17276 34144 17282 34196
rect 19702 34144 19708 34196
rect 19760 34184 19766 34196
rect 19797 34187 19855 34193
rect 19797 34184 19809 34187
rect 19760 34156 19809 34184
rect 19760 34144 19766 34156
rect 19797 34153 19809 34156
rect 19843 34153 19855 34187
rect 22830 34184 22836 34196
rect 19797 34147 19855 34153
rect 20272 34156 22836 34184
rect 15378 34048 15384 34060
rect 15339 34020 15384 34048
rect 15378 34008 15384 34020
rect 15436 34008 15442 34060
rect 17402 34008 17408 34060
rect 17460 34048 17466 34060
rect 17497 34051 17555 34057
rect 17497 34048 17509 34051
rect 17460 34020 17509 34048
rect 17460 34008 17466 34020
rect 17497 34017 17509 34020
rect 17543 34017 17555 34051
rect 17497 34011 17555 34017
rect 20272 33992 20300 34156
rect 22830 34144 22836 34156
rect 22888 34144 22894 34196
rect 22925 34187 22983 34193
rect 22925 34153 22937 34187
rect 22971 34184 22983 34187
rect 23382 34184 23388 34196
rect 22971 34156 23388 34184
rect 22971 34153 22983 34156
rect 22925 34147 22983 34153
rect 23382 34144 23388 34156
rect 23440 34144 23446 34196
rect 24854 34184 24860 34196
rect 24815 34156 24860 34184
rect 24854 34144 24860 34156
rect 24912 34144 24918 34196
rect 26053 34187 26111 34193
rect 26053 34153 26065 34187
rect 26099 34184 26111 34187
rect 26878 34184 26884 34196
rect 26099 34156 26884 34184
rect 26099 34153 26111 34156
rect 26053 34147 26111 34153
rect 26878 34144 26884 34156
rect 26936 34144 26942 34196
rect 27617 34187 27675 34193
rect 27617 34153 27629 34187
rect 27663 34184 27675 34187
rect 27798 34184 27804 34196
rect 27663 34156 27804 34184
rect 27663 34153 27675 34156
rect 27617 34147 27675 34153
rect 27798 34144 27804 34156
rect 27856 34144 27862 34196
rect 28350 34184 28356 34196
rect 28311 34156 28356 34184
rect 28350 34144 28356 34156
rect 28408 34144 28414 34196
rect 29733 34187 29791 34193
rect 29733 34153 29745 34187
rect 29779 34184 29791 34187
rect 30374 34184 30380 34196
rect 29779 34156 30380 34184
rect 29779 34153 29791 34156
rect 29733 34147 29791 34153
rect 30374 34144 30380 34156
rect 30432 34144 30438 34196
rect 30926 34184 30932 34196
rect 30576 34156 30932 34184
rect 20806 34076 20812 34128
rect 20864 34116 20870 34128
rect 20993 34119 21051 34125
rect 20993 34116 21005 34119
rect 20864 34088 21005 34116
rect 20864 34076 20870 34088
rect 20993 34085 21005 34088
rect 21039 34085 21051 34119
rect 22370 34116 22376 34128
rect 20993 34079 21051 34085
rect 21376 34088 22376 34116
rect 20441 34051 20499 34057
rect 20441 34017 20453 34051
rect 20487 34048 20499 34051
rect 20714 34048 20720 34060
rect 20487 34020 20720 34048
rect 20487 34017 20499 34020
rect 20441 34011 20499 34017
rect 20714 34008 20720 34020
rect 20772 34008 20778 34060
rect 17773 33983 17831 33989
rect 17773 33949 17785 33983
rect 17819 33980 17831 33983
rect 17862 33980 17868 33992
rect 17819 33952 17868 33980
rect 17819 33949 17831 33952
rect 17773 33943 17831 33949
rect 17862 33940 17868 33952
rect 17920 33940 17926 33992
rect 19978 33980 19984 33992
rect 19939 33952 19984 33980
rect 19978 33940 19984 33952
rect 20036 33940 20042 33992
rect 20165 33983 20223 33989
rect 20165 33949 20177 33983
rect 20211 33949 20223 33983
rect 20165 33943 20223 33949
rect 15648 33915 15706 33921
rect 15648 33881 15660 33915
rect 15694 33912 15706 33915
rect 16206 33912 16212 33924
rect 15694 33884 16212 33912
rect 15694 33881 15706 33884
rect 15648 33875 15706 33881
rect 16206 33872 16212 33884
rect 16264 33872 16270 33924
rect 20073 33915 20131 33921
rect 20073 33881 20085 33915
rect 20119 33881 20131 33915
rect 20180 33912 20208 33943
rect 20254 33940 20260 33992
rect 20312 33989 20318 33992
rect 20312 33983 20341 33989
rect 20329 33980 20341 33983
rect 21376 33980 21404 34088
rect 22370 34076 22376 34088
rect 22428 34116 22434 34128
rect 23290 34116 23296 34128
rect 22428 34088 23296 34116
rect 22428 34076 22434 34088
rect 23290 34076 23296 34088
rect 23348 34076 23354 34128
rect 21453 34051 21511 34057
rect 21453 34017 21465 34051
rect 21499 34048 21511 34051
rect 24026 34048 24032 34060
rect 21499 34020 22232 34048
rect 21499 34017 21511 34020
rect 21453 34011 21511 34017
rect 21545 33983 21603 33989
rect 21545 33980 21557 33983
rect 20329 33952 20405 33980
rect 21376 33952 21557 33980
rect 20329 33949 20341 33952
rect 20312 33943 20341 33949
rect 21545 33949 21557 33952
rect 21591 33949 21603 33983
rect 22094 33980 22100 33992
rect 21545 33943 21603 33949
rect 21652 33952 22100 33980
rect 20312 33940 20318 33943
rect 20990 33912 20996 33924
rect 20180 33884 20996 33912
rect 20073 33875 20131 33881
rect 12158 33804 12164 33856
rect 12216 33844 12222 33856
rect 18874 33844 18880 33856
rect 12216 33816 18880 33844
rect 12216 33804 12222 33816
rect 18874 33804 18880 33816
rect 18932 33804 18938 33856
rect 20088 33844 20116 33875
rect 20990 33872 20996 33884
rect 21048 33872 21054 33924
rect 21652 33844 21680 33952
rect 22094 33940 22100 33952
rect 22152 33940 22158 33992
rect 22204 33989 22232 34020
rect 22388 34020 24032 34048
rect 22388 33992 22416 34020
rect 24026 34008 24032 34020
rect 24084 34008 24090 34060
rect 26513 34051 26571 34057
rect 26513 34048 26525 34051
rect 25056 34020 26525 34048
rect 22189 33983 22247 33989
rect 22189 33949 22201 33983
rect 22235 33980 22247 33983
rect 22278 33980 22284 33992
rect 22235 33952 22284 33980
rect 22235 33949 22247 33952
rect 22189 33943 22247 33949
rect 22278 33940 22284 33952
rect 22336 33940 22342 33992
rect 22370 33940 22376 33992
rect 22428 33980 22434 33992
rect 25056 33989 25084 34020
rect 26513 34017 26525 34020
rect 26559 34017 26571 34051
rect 29638 34048 29644 34060
rect 26513 34011 26571 34017
rect 26712 34020 27568 34048
rect 22833 33983 22891 33989
rect 22428 33952 22521 33980
rect 22428 33940 22434 33952
rect 22833 33949 22845 33983
rect 22879 33949 22891 33983
rect 22833 33943 22891 33949
rect 25041 33983 25099 33989
rect 25041 33949 25053 33983
rect 25087 33949 25099 33983
rect 25041 33943 25099 33949
rect 21729 33915 21787 33921
rect 21729 33881 21741 33915
rect 21775 33912 21787 33915
rect 21818 33912 21824 33924
rect 21775 33884 21824 33912
rect 21775 33881 21787 33884
rect 21729 33875 21787 33881
rect 21818 33872 21824 33884
rect 21876 33872 21882 33924
rect 22848 33912 22876 33943
rect 25130 33940 25136 33992
rect 25188 33980 25194 33992
rect 25498 33980 25504 33992
rect 25188 33952 25504 33980
rect 25188 33940 25194 33952
rect 25498 33940 25504 33952
rect 25556 33940 25562 33992
rect 25682 33980 25688 33992
rect 25643 33952 25688 33980
rect 25682 33940 25688 33952
rect 25740 33940 25746 33992
rect 25866 33980 25872 33992
rect 25827 33952 25872 33980
rect 25866 33940 25872 33952
rect 25924 33940 25930 33992
rect 26712 33989 26740 34020
rect 27540 33992 27568 34020
rect 27816 34020 29644 34048
rect 26697 33983 26755 33989
rect 26697 33949 26709 33983
rect 26743 33949 26755 33983
rect 26878 33980 26884 33992
rect 26839 33952 26884 33980
rect 26697 33943 26755 33949
rect 26878 33940 26884 33952
rect 26936 33940 26942 33992
rect 27154 33980 27160 33992
rect 27115 33952 27160 33980
rect 27154 33940 27160 33952
rect 27212 33940 27218 33992
rect 27522 33940 27528 33992
rect 27580 33980 27586 33992
rect 27816 33989 27844 34020
rect 29638 34008 29644 34020
rect 29696 34008 29702 34060
rect 30576 34057 30604 34156
rect 30926 34144 30932 34156
rect 30984 34184 30990 34196
rect 31662 34184 31668 34196
rect 30984 34156 31668 34184
rect 30984 34144 30990 34156
rect 31662 34144 31668 34156
rect 31720 34144 31726 34196
rect 32401 34187 32459 34193
rect 32401 34153 32413 34187
rect 32447 34184 32459 34187
rect 32490 34184 32496 34196
rect 32447 34156 32496 34184
rect 32447 34153 32459 34156
rect 32401 34147 32459 34153
rect 32490 34144 32496 34156
rect 32548 34144 32554 34196
rect 36633 34187 36691 34193
rect 36633 34153 36645 34187
rect 36679 34184 36691 34187
rect 37366 34184 37372 34196
rect 36679 34156 37372 34184
rect 36679 34153 36691 34156
rect 36633 34147 36691 34153
rect 37366 34144 37372 34156
rect 37424 34144 37430 34196
rect 38749 34187 38807 34193
rect 38749 34153 38761 34187
rect 38795 34153 38807 34187
rect 41230 34184 41236 34196
rect 38749 34147 38807 34153
rect 38856 34156 41236 34184
rect 31938 34116 31944 34128
rect 31851 34088 31944 34116
rect 31938 34076 31944 34088
rect 31996 34116 32002 34128
rect 32950 34116 32956 34128
rect 31996 34088 32956 34116
rect 31996 34076 32002 34088
rect 32950 34076 32956 34088
rect 33008 34116 33014 34128
rect 33505 34119 33563 34125
rect 33505 34116 33517 34119
rect 33008 34088 33517 34116
rect 33008 34076 33014 34088
rect 33505 34085 33517 34088
rect 33551 34085 33563 34119
rect 33505 34079 33563 34085
rect 34330 34076 34336 34128
rect 34388 34116 34394 34128
rect 34388 34088 35894 34116
rect 34388 34076 34394 34088
rect 30561 34051 30619 34057
rect 30561 34017 30573 34051
rect 30607 34017 30619 34051
rect 30561 34011 30619 34017
rect 32769 34051 32827 34057
rect 32769 34017 32781 34051
rect 32815 34048 32827 34051
rect 32968 34048 32996 34076
rect 35342 34048 35348 34060
rect 32815 34020 32996 34048
rect 35303 34020 35348 34048
rect 32815 34017 32827 34020
rect 32769 34011 32827 34017
rect 35342 34008 35348 34020
rect 35400 34008 35406 34060
rect 35866 34048 35894 34088
rect 36078 34076 36084 34128
rect 36136 34116 36142 34128
rect 38562 34116 38568 34128
rect 36136 34088 38568 34116
rect 36136 34076 36142 34088
rect 38562 34076 38568 34088
rect 38620 34116 38626 34128
rect 38764 34116 38792 34147
rect 38620 34088 38792 34116
rect 38620 34076 38626 34088
rect 37369 34051 37427 34057
rect 37369 34048 37381 34051
rect 35866 34020 37381 34048
rect 37369 34017 37381 34020
rect 37415 34048 37427 34051
rect 38856 34048 38884 34156
rect 41230 34144 41236 34156
rect 41288 34144 41294 34196
rect 39942 34048 39948 34060
rect 37415 34020 38884 34048
rect 39903 34020 39948 34048
rect 37415 34017 37427 34020
rect 37369 34011 37427 34017
rect 39942 34008 39948 34020
rect 40000 34008 40006 34060
rect 42334 34048 42340 34060
rect 42295 34020 42340 34048
rect 42334 34008 42340 34020
rect 42392 34008 42398 34060
rect 44082 34048 44088 34060
rect 44043 34020 44088 34048
rect 44082 34008 44088 34020
rect 44140 34008 44146 34060
rect 27617 33983 27675 33989
rect 27617 33980 27629 33983
rect 27580 33952 27629 33980
rect 27580 33940 27586 33952
rect 27617 33949 27629 33952
rect 27663 33949 27675 33983
rect 27617 33943 27675 33949
rect 27801 33983 27859 33989
rect 27801 33949 27813 33983
rect 27847 33949 27859 33983
rect 28258 33980 28264 33992
rect 28219 33952 28264 33980
rect 27801 33943 27859 33949
rect 28258 33940 28264 33952
rect 28316 33940 28322 33992
rect 29454 33940 29460 33992
rect 29512 33980 29518 33992
rect 29549 33983 29607 33989
rect 29549 33980 29561 33983
rect 29512 33952 29561 33980
rect 29512 33940 29518 33952
rect 29549 33949 29561 33952
rect 29595 33949 29607 33983
rect 29549 33943 29607 33949
rect 32122 33940 32128 33992
rect 32180 33980 32186 33992
rect 32582 33980 32588 33992
rect 32180 33952 32588 33980
rect 32180 33940 32186 33952
rect 32582 33940 32588 33952
rect 32640 33940 32646 33992
rect 33134 33940 33140 33992
rect 33192 33980 33198 33992
rect 33410 33980 33416 33992
rect 33192 33952 33416 33980
rect 33192 33940 33198 33952
rect 33410 33940 33416 33952
rect 33468 33980 33474 33992
rect 33689 33983 33747 33989
rect 33689 33980 33701 33983
rect 33468 33952 33701 33980
rect 33468 33940 33474 33952
rect 33689 33949 33701 33952
rect 33735 33949 33747 33983
rect 33689 33943 33747 33949
rect 34238 33940 34244 33992
rect 34296 33980 34302 33992
rect 34701 33983 34759 33989
rect 34701 33980 34713 33983
rect 34296 33952 34713 33980
rect 34296 33940 34302 33952
rect 34701 33949 34713 33952
rect 34747 33949 34759 33983
rect 34701 33943 34759 33949
rect 34885 33983 34943 33989
rect 34885 33949 34897 33983
rect 34931 33980 34943 33983
rect 35434 33980 35440 33992
rect 34931 33952 35440 33980
rect 34931 33949 34943 33952
rect 34885 33943 34943 33949
rect 35434 33940 35440 33952
rect 35492 33980 35498 33992
rect 35529 33983 35587 33989
rect 35529 33980 35541 33983
rect 35492 33952 35541 33980
rect 35492 33940 35498 33952
rect 35529 33949 35541 33952
rect 35575 33949 35587 33983
rect 35529 33943 35587 33949
rect 35621 33983 35679 33989
rect 35621 33949 35633 33983
rect 35667 33980 35679 33983
rect 36081 33983 36139 33989
rect 36081 33980 36093 33983
rect 35667 33952 36093 33980
rect 35667 33949 35679 33952
rect 35621 33943 35679 33949
rect 36081 33949 36093 33952
rect 36127 33980 36139 33983
rect 36906 33980 36912 33992
rect 36127 33952 36912 33980
rect 36127 33949 36139 33952
rect 36081 33943 36139 33949
rect 36906 33940 36912 33952
rect 36964 33940 36970 33992
rect 37093 33983 37151 33989
rect 37093 33949 37105 33983
rect 37139 33949 37151 33983
rect 37093 33943 37151 33949
rect 22296 33884 22876 33912
rect 26789 33915 26847 33921
rect 20088 33816 21680 33844
rect 22186 33804 22192 33856
rect 22244 33844 22250 33856
rect 22296 33853 22324 33884
rect 26789 33881 26801 33915
rect 26835 33881 26847 33915
rect 26970 33912 26976 33924
rect 26929 33884 26976 33912
rect 26789 33875 26847 33881
rect 22281 33847 22339 33853
rect 22281 33844 22293 33847
rect 22244 33816 22293 33844
rect 22244 33804 22250 33816
rect 22281 33813 22293 33816
rect 22327 33813 22339 33847
rect 26804 33844 26832 33875
rect 26970 33872 26976 33884
rect 27028 33921 27034 33924
rect 27028 33915 27077 33921
rect 27028 33881 27031 33915
rect 27065 33912 27077 33915
rect 28994 33912 29000 33924
rect 27065 33884 29000 33912
rect 27065 33881 27077 33884
rect 27028 33875 27077 33881
rect 27028 33872 27034 33875
rect 28994 33872 29000 33884
rect 29052 33872 29058 33924
rect 30828 33915 30886 33921
rect 30828 33881 30840 33915
rect 30874 33912 30886 33915
rect 31478 33912 31484 33924
rect 30874 33884 31484 33912
rect 30874 33881 30886 33884
rect 30828 33875 30886 33881
rect 31478 33872 31484 33884
rect 31536 33872 31542 33924
rect 27430 33844 27436 33856
rect 26804 33816 27436 33844
rect 22281 33807 22339 33813
rect 27430 33804 27436 33816
rect 27488 33804 27494 33856
rect 32600 33844 32628 33940
rect 33781 33915 33839 33921
rect 33781 33881 33793 33915
rect 33827 33912 33839 33915
rect 33962 33912 33968 33924
rect 33827 33884 33968 33912
rect 33827 33881 33839 33884
rect 33781 33875 33839 33881
rect 33962 33872 33968 33884
rect 34020 33872 34026 33924
rect 36170 33872 36176 33924
rect 36228 33912 36234 33924
rect 36449 33915 36507 33921
rect 36449 33912 36461 33915
rect 36228 33884 36461 33912
rect 36228 33872 36234 33884
rect 36449 33881 36461 33884
rect 36495 33881 36507 33915
rect 36449 33875 36507 33881
rect 33873 33847 33931 33853
rect 33873 33844 33885 33847
rect 32600 33816 33885 33844
rect 33873 33813 33885 33816
rect 33919 33813 33931 33847
rect 34054 33844 34060 33856
rect 34015 33816 34060 33844
rect 33873 33807 33931 33813
rect 34054 33804 34060 33816
rect 34112 33804 34118 33856
rect 34790 33844 34796 33856
rect 34751 33816 34796 33844
rect 34790 33804 34796 33816
rect 34848 33804 34854 33856
rect 35345 33847 35403 33853
rect 35345 33813 35357 33847
rect 35391 33844 35403 33847
rect 35618 33844 35624 33856
rect 35391 33816 35624 33844
rect 35391 33813 35403 33816
rect 35345 33807 35403 33813
rect 35618 33804 35624 33816
rect 35676 33804 35682 33856
rect 36262 33844 36268 33856
rect 36223 33816 36268 33844
rect 36262 33804 36268 33816
rect 36320 33804 36326 33856
rect 36354 33804 36360 33856
rect 36412 33844 36418 33856
rect 37108 33844 37136 33943
rect 37182 33940 37188 33992
rect 37240 33980 37246 33992
rect 38381 33983 38439 33989
rect 37240 33952 37285 33980
rect 37240 33940 37246 33952
rect 38381 33949 38393 33983
rect 38427 33980 38439 33983
rect 38838 33980 38844 33992
rect 38427 33952 38844 33980
rect 38427 33949 38439 33952
rect 38381 33943 38439 33949
rect 38838 33940 38844 33952
rect 38896 33940 38902 33992
rect 40218 33989 40224 33992
rect 40212 33980 40224 33989
rect 40179 33952 40224 33980
rect 40212 33943 40224 33952
rect 40218 33940 40224 33943
rect 40276 33940 40282 33992
rect 38746 33912 38752 33924
rect 38707 33884 38752 33912
rect 38746 33872 38752 33884
rect 38804 33872 38810 33924
rect 42521 33915 42579 33921
rect 42521 33881 42533 33915
rect 42567 33912 42579 33915
rect 43530 33912 43536 33924
rect 42567 33884 43536 33912
rect 42567 33881 42579 33884
rect 42521 33875 42579 33881
rect 43530 33872 43536 33884
rect 43588 33872 43594 33924
rect 36412 33816 37136 33844
rect 36412 33804 36418 33816
rect 37274 33804 37280 33856
rect 37332 33844 37338 33856
rect 37369 33847 37427 33853
rect 37369 33844 37381 33847
rect 37332 33816 37381 33844
rect 37332 33804 37338 33816
rect 37369 33813 37381 33816
rect 37415 33813 37427 33847
rect 37369 33807 37427 33813
rect 38933 33847 38991 33853
rect 38933 33813 38945 33847
rect 38979 33844 38991 33847
rect 39114 33844 39120 33856
rect 38979 33816 39120 33844
rect 38979 33813 38991 33816
rect 38933 33807 38991 33813
rect 39114 33804 39120 33816
rect 39172 33804 39178 33856
rect 40034 33804 40040 33856
rect 40092 33844 40098 33856
rect 41325 33847 41383 33853
rect 41325 33844 41337 33847
rect 40092 33816 41337 33844
rect 40092 33804 40098 33816
rect 41325 33813 41337 33816
rect 41371 33813 41383 33847
rect 41325 33807 41383 33813
rect 1104 33754 44896 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 44896 33754
rect 1104 33680 44896 33702
rect 18598 33640 18604 33652
rect 15948 33612 18604 33640
rect 15948 33513 15976 33612
rect 18598 33600 18604 33612
rect 18656 33600 18662 33652
rect 18690 33600 18696 33652
rect 18748 33640 18754 33652
rect 18785 33643 18843 33649
rect 18785 33640 18797 33643
rect 18748 33612 18797 33640
rect 18748 33600 18754 33612
rect 18785 33609 18797 33612
rect 18831 33609 18843 33643
rect 18785 33603 18843 33609
rect 18874 33600 18880 33652
rect 18932 33640 18938 33652
rect 35986 33640 35992 33652
rect 18932 33612 35992 33640
rect 18932 33600 18938 33612
rect 35986 33600 35992 33612
rect 36044 33600 36050 33652
rect 36262 33600 36268 33652
rect 36320 33640 36326 33652
rect 37550 33640 37556 33652
rect 36320 33612 37556 33640
rect 36320 33600 36326 33612
rect 37550 33600 37556 33612
rect 37608 33600 37614 33652
rect 38378 33600 38384 33652
rect 38436 33649 38442 33652
rect 38436 33643 38455 33649
rect 38443 33609 38455 33643
rect 38436 33603 38455 33609
rect 38565 33643 38623 33649
rect 38565 33609 38577 33643
rect 38611 33609 38623 33643
rect 38565 33603 38623 33609
rect 39761 33643 39819 33649
rect 39761 33609 39773 33643
rect 39807 33640 39819 33643
rect 40126 33640 40132 33652
rect 39807 33612 40132 33640
rect 39807 33609 39819 33612
rect 39761 33603 39819 33609
rect 38436 33600 38442 33603
rect 18417 33575 18475 33581
rect 18417 33541 18429 33575
rect 18463 33572 18475 33575
rect 19334 33572 19340 33584
rect 18463 33544 19340 33572
rect 18463 33541 18475 33544
rect 18417 33535 18475 33541
rect 19334 33532 19340 33544
rect 19392 33532 19398 33584
rect 19426 33532 19432 33584
rect 19484 33581 19490 33584
rect 19484 33575 19548 33581
rect 19484 33541 19502 33575
rect 19536 33541 19548 33575
rect 19484 33535 19548 33541
rect 19484 33532 19490 33535
rect 19978 33532 19984 33584
rect 20036 33572 20042 33584
rect 21177 33575 21235 33581
rect 21177 33572 21189 33575
rect 20036 33544 21189 33572
rect 20036 33532 20042 33544
rect 21177 33541 21189 33544
rect 21223 33572 21235 33575
rect 22370 33572 22376 33584
rect 21223 33544 22376 33572
rect 21223 33541 21235 33544
rect 21177 33535 21235 33541
rect 22370 33532 22376 33544
rect 22428 33532 22434 33584
rect 23290 33532 23296 33584
rect 23348 33572 23354 33584
rect 23569 33575 23627 33581
rect 23569 33572 23581 33575
rect 23348 33544 23581 33572
rect 23348 33532 23354 33544
rect 23569 33541 23581 33544
rect 23615 33541 23627 33575
rect 24486 33572 24492 33584
rect 24447 33544 24492 33572
rect 23569 33535 23627 33541
rect 24486 33532 24492 33544
rect 24544 33532 24550 33584
rect 24673 33575 24731 33581
rect 24673 33541 24685 33575
rect 24719 33572 24731 33575
rect 29641 33575 29699 33581
rect 29641 33572 29653 33575
rect 24719 33544 29653 33572
rect 24719 33541 24731 33544
rect 24673 33535 24731 33541
rect 29641 33541 29653 33544
rect 29687 33541 29699 33575
rect 31478 33572 31484 33584
rect 31439 33544 31484 33572
rect 29641 33535 29699 33541
rect 15933 33507 15991 33513
rect 15933 33473 15945 33507
rect 15979 33473 15991 33507
rect 15933 33467 15991 33473
rect 16117 33507 16175 33513
rect 16117 33473 16129 33507
rect 16163 33504 16175 33507
rect 16942 33504 16948 33516
rect 16163 33476 16528 33504
rect 16903 33476 16948 33504
rect 16163 33473 16175 33476
rect 16117 33467 16175 33473
rect 16500 33380 16528 33476
rect 16942 33464 16948 33476
rect 17000 33464 17006 33516
rect 17586 33464 17592 33516
rect 17644 33504 17650 33516
rect 17770 33504 17776 33516
rect 17644 33476 17776 33504
rect 17644 33464 17650 33476
rect 17770 33464 17776 33476
rect 17828 33504 17834 33516
rect 18233 33507 18291 33513
rect 18233 33504 18245 33507
rect 17828 33476 18245 33504
rect 17828 33464 17834 33476
rect 18233 33473 18245 33476
rect 18279 33473 18291 33507
rect 18233 33467 18291 33473
rect 18509 33507 18567 33513
rect 18509 33473 18521 33507
rect 18555 33473 18567 33507
rect 18509 33467 18567 33473
rect 18601 33507 18659 33513
rect 18601 33473 18613 33507
rect 18647 33504 18659 33507
rect 20254 33504 20260 33516
rect 18647 33476 20260 33504
rect 18647 33473 18659 33476
rect 18601 33467 18659 33473
rect 17221 33439 17279 33445
rect 17221 33405 17233 33439
rect 17267 33405 17279 33439
rect 17221 33399 17279 33405
rect 16482 33328 16488 33380
rect 16540 33368 16546 33380
rect 17236 33368 17264 33399
rect 17862 33396 17868 33448
rect 17920 33436 17926 33448
rect 18524 33436 18552 33467
rect 20254 33464 20260 33476
rect 20312 33464 20318 33516
rect 20714 33464 20720 33516
rect 20772 33504 20778 33516
rect 21085 33507 21143 33513
rect 21085 33504 21097 33507
rect 20772 33476 21097 33504
rect 20772 33464 20778 33476
rect 21085 33473 21097 33476
rect 21131 33473 21143 33507
rect 21266 33504 21272 33516
rect 21227 33476 21272 33504
rect 21085 33467 21143 33473
rect 21266 33464 21272 33476
rect 21324 33464 21330 33516
rect 22462 33504 22468 33516
rect 22066 33476 22468 33504
rect 19242 33436 19248 33448
rect 17920 33408 18552 33436
rect 19203 33408 19248 33436
rect 17920 33396 17926 33408
rect 19242 33396 19248 33408
rect 19300 33396 19306 33448
rect 20806 33396 20812 33448
rect 20864 33436 20870 33448
rect 22066 33436 22094 33476
rect 22462 33464 22468 33476
rect 22520 33504 22526 33516
rect 22833 33507 22891 33513
rect 22833 33504 22845 33507
rect 22520 33476 22845 33504
rect 22520 33464 22526 33476
rect 22833 33473 22845 33476
rect 22879 33473 22891 33507
rect 22833 33467 22891 33473
rect 22925 33507 22983 33513
rect 22925 33473 22937 33507
rect 22971 33504 22983 33507
rect 23658 33504 23664 33516
rect 22971 33476 23664 33504
rect 22971 33473 22983 33476
rect 22925 33467 22983 33473
rect 23658 33464 23664 33476
rect 23716 33464 23722 33516
rect 25958 33504 25964 33516
rect 25919 33476 25964 33504
rect 25958 33464 25964 33476
rect 26016 33464 26022 33516
rect 26973 33507 27031 33513
rect 26973 33473 26985 33507
rect 27019 33473 27031 33507
rect 27154 33504 27160 33516
rect 27115 33476 27160 33504
rect 26973 33467 27031 33473
rect 20864 33408 22094 33436
rect 20864 33396 20870 33408
rect 22186 33396 22192 33448
rect 22244 33436 22250 33448
rect 22649 33439 22707 33445
rect 22649 33436 22661 33439
rect 22244 33408 22661 33436
rect 22244 33396 22250 33408
rect 22649 33405 22661 33408
rect 22695 33405 22707 33439
rect 22649 33399 22707 33405
rect 22738 33396 22744 33448
rect 22796 33436 22802 33448
rect 23198 33436 23204 33448
rect 22796 33408 23204 33436
rect 22796 33396 22802 33408
rect 23198 33396 23204 33408
rect 23256 33396 23262 33448
rect 25682 33396 25688 33448
rect 25740 33436 25746 33448
rect 26050 33436 26056 33448
rect 25740 33408 26056 33436
rect 25740 33396 25746 33408
rect 26050 33396 26056 33408
rect 26108 33436 26114 33448
rect 26988 33436 27016 33467
rect 27154 33464 27160 33476
rect 27212 33464 27218 33516
rect 27798 33464 27804 33516
rect 27856 33504 27862 33516
rect 27893 33507 27951 33513
rect 27893 33504 27905 33507
rect 27856 33476 27905 33504
rect 27856 33464 27862 33476
rect 27893 33473 27905 33476
rect 27939 33473 27951 33507
rect 28074 33504 28080 33516
rect 28035 33476 28080 33504
rect 27893 33467 27951 33473
rect 28074 33464 28080 33476
rect 28132 33464 28138 33516
rect 29454 33504 29460 33516
rect 29415 33476 29460 33504
rect 29454 33464 29460 33476
rect 29512 33464 29518 33516
rect 27982 33436 27988 33448
rect 26108 33408 27016 33436
rect 27943 33408 27988 33436
rect 26108 33396 26114 33408
rect 27982 33396 27988 33408
rect 28040 33396 28046 33448
rect 28169 33439 28227 33445
rect 28169 33405 28181 33439
rect 28215 33436 28227 33439
rect 28258 33436 28264 33448
rect 28215 33408 28264 33436
rect 28215 33405 28227 33408
rect 28169 33399 28227 33405
rect 28258 33396 28264 33408
rect 28316 33436 28322 33448
rect 28626 33436 28632 33448
rect 28316 33408 28632 33436
rect 28316 33396 28322 33408
rect 28626 33396 28632 33408
rect 28684 33396 28690 33448
rect 17954 33368 17960 33380
rect 16540 33340 17960 33368
rect 16540 33328 16546 33340
rect 17954 33328 17960 33340
rect 18012 33328 18018 33380
rect 20625 33371 20683 33377
rect 20625 33337 20637 33371
rect 20671 33368 20683 33371
rect 20714 33368 20720 33380
rect 20671 33340 20720 33368
rect 20671 33337 20683 33340
rect 20625 33331 20683 33337
rect 20714 33328 20720 33340
rect 20772 33328 20778 33380
rect 21818 33328 21824 33380
rect 21876 33368 21882 33380
rect 24762 33368 24768 33380
rect 21876 33340 24768 33368
rect 21876 33328 21882 33340
rect 24762 33328 24768 33340
rect 24820 33328 24826 33380
rect 25774 33368 25780 33380
rect 25687 33340 25780 33368
rect 25774 33328 25780 33340
rect 25832 33368 25838 33380
rect 26970 33368 26976 33380
rect 25832 33340 26976 33368
rect 25832 33328 25838 33340
rect 26970 33328 26976 33340
rect 27028 33328 27034 33380
rect 29656 33368 29684 33535
rect 31478 33532 31484 33544
rect 31536 33532 31542 33584
rect 32490 33572 32496 33584
rect 31588 33544 32496 33572
rect 31588 33513 31616 33544
rect 32490 33532 32496 33544
rect 32548 33532 32554 33584
rect 34238 33572 34244 33584
rect 34199 33544 34244 33572
rect 34238 33532 34244 33544
rect 34296 33532 34302 33584
rect 35434 33532 35440 33584
rect 35492 33572 35498 33584
rect 36449 33575 36507 33581
rect 35492 33544 36400 33572
rect 35492 33532 35498 33544
rect 31389 33507 31447 33513
rect 31389 33473 31401 33507
rect 31435 33473 31447 33507
rect 31389 33467 31447 33473
rect 31573 33507 31631 33513
rect 31573 33473 31585 33507
rect 31619 33473 31631 33507
rect 31573 33467 31631 33473
rect 31404 33436 31432 33467
rect 31662 33464 31668 33516
rect 31720 33504 31726 33516
rect 32125 33507 32183 33513
rect 32125 33504 32137 33507
rect 31720 33476 32137 33504
rect 31720 33464 31726 33476
rect 32125 33473 32137 33476
rect 32171 33473 32183 33507
rect 32125 33467 32183 33473
rect 32392 33507 32450 33513
rect 32392 33473 32404 33507
rect 32438 33504 32450 33507
rect 32674 33504 32680 33516
rect 32438 33476 32680 33504
rect 32438 33473 32450 33476
rect 32392 33467 32450 33473
rect 32674 33464 32680 33476
rect 32732 33464 32738 33516
rect 33962 33504 33968 33516
rect 33923 33476 33968 33504
rect 33962 33464 33968 33476
rect 34020 33464 34026 33516
rect 34054 33464 34060 33516
rect 34112 33504 34118 33516
rect 35621 33507 35679 33513
rect 35621 33504 35633 33507
rect 34112 33476 35633 33504
rect 34112 33464 34118 33476
rect 35621 33473 35633 33476
rect 35667 33504 35679 33507
rect 36170 33504 36176 33516
rect 35667 33476 36176 33504
rect 35667 33473 35679 33476
rect 35621 33467 35679 33473
rect 36170 33464 36176 33476
rect 36228 33464 36234 33516
rect 36372 33504 36400 33544
rect 36449 33541 36461 33575
rect 36495 33572 36507 33575
rect 37737 33575 37795 33581
rect 37737 33572 37749 33575
rect 36495 33544 37749 33572
rect 36495 33541 36507 33544
rect 36449 33535 36507 33541
rect 37737 33541 37749 33544
rect 37783 33541 37795 33575
rect 38194 33572 38200 33584
rect 38155 33544 38200 33572
rect 37737 33535 37795 33541
rect 38194 33532 38200 33544
rect 38252 33532 38258 33584
rect 38580 33572 38608 33603
rect 40126 33600 40132 33612
rect 40184 33600 40190 33652
rect 43530 33640 43536 33652
rect 43491 33612 43536 33640
rect 43530 33600 43536 33612
rect 43588 33600 43594 33652
rect 38838 33572 38844 33584
rect 38580 33544 38844 33572
rect 38838 33532 38844 33544
rect 38896 33572 38902 33584
rect 39853 33575 39911 33581
rect 38896 33544 39804 33572
rect 38896 33532 38902 33544
rect 39776 33516 39804 33544
rect 39853 33541 39865 33575
rect 39899 33572 39911 33575
rect 40034 33572 40040 33584
rect 39899 33544 40040 33572
rect 39899 33541 39911 33544
rect 39853 33535 39911 33541
rect 40034 33532 40040 33544
rect 40092 33532 40098 33584
rect 37277 33507 37335 33513
rect 37277 33504 37289 33507
rect 36372 33476 37289 33504
rect 37277 33473 37289 33476
rect 37323 33473 37335 33507
rect 37277 33467 37335 33473
rect 37369 33507 37427 33513
rect 37369 33473 37381 33507
rect 37415 33473 37427 33507
rect 37550 33504 37556 33516
rect 37511 33476 37556 33504
rect 37369 33467 37427 33473
rect 32030 33436 32036 33448
rect 31404 33408 32036 33436
rect 32030 33396 32036 33408
rect 32088 33396 32094 33448
rect 33134 33396 33140 33448
rect 33192 33436 33198 33448
rect 34241 33439 34299 33445
rect 33192 33408 34100 33436
rect 33192 33396 33198 33408
rect 29656 33340 31754 33368
rect 16025 33303 16083 33309
rect 16025 33269 16037 33303
rect 16071 33300 16083 33303
rect 16666 33300 16672 33312
rect 16071 33272 16672 33300
rect 16071 33269 16083 33272
rect 16025 33263 16083 33269
rect 16666 33260 16672 33272
rect 16724 33260 16730 33312
rect 18598 33260 18604 33312
rect 18656 33300 18662 33312
rect 21358 33300 21364 33312
rect 18656 33272 21364 33300
rect 18656 33260 18662 33272
rect 21358 33260 21364 33272
rect 21416 33260 21422 33312
rect 22370 33260 22376 33312
rect 22428 33300 22434 33312
rect 22465 33303 22523 33309
rect 22465 33300 22477 33303
rect 22428 33272 22477 33300
rect 22428 33260 22434 33272
rect 22465 33269 22477 33272
rect 22511 33269 22523 33303
rect 27062 33300 27068 33312
rect 27023 33272 27068 33300
rect 22465 33263 22523 33269
rect 27062 33260 27068 33272
rect 27120 33260 27126 33312
rect 27709 33303 27767 33309
rect 27709 33269 27721 33303
rect 27755 33300 27767 33303
rect 27890 33300 27896 33312
rect 27755 33272 27896 33300
rect 27755 33269 27767 33272
rect 27709 33263 27767 33269
rect 27890 33260 27896 33272
rect 27948 33260 27954 33312
rect 31726 33300 31754 33340
rect 33410 33328 33416 33380
rect 33468 33368 33474 33380
rect 34072 33377 34100 33408
rect 34241 33405 34253 33439
rect 34287 33436 34299 33439
rect 34330 33436 34336 33448
rect 34287 33408 34336 33436
rect 34287 33405 34299 33408
rect 34241 33399 34299 33405
rect 33505 33371 33563 33377
rect 33505 33368 33517 33371
rect 33468 33340 33517 33368
rect 33468 33328 33474 33340
rect 33505 33337 33517 33340
rect 33551 33337 33563 33371
rect 33505 33331 33563 33337
rect 34057 33371 34115 33377
rect 34057 33337 34069 33371
rect 34103 33337 34115 33371
rect 34057 33331 34115 33337
rect 33134 33300 33140 33312
rect 31726 33272 33140 33300
rect 33134 33260 33140 33272
rect 33192 33260 33198 33312
rect 33226 33260 33232 33312
rect 33284 33300 33290 33312
rect 34256 33300 34284 33399
rect 34330 33396 34336 33408
rect 34388 33396 34394 33448
rect 35345 33439 35403 33445
rect 35345 33405 35357 33439
rect 35391 33436 35403 33439
rect 35434 33436 35440 33448
rect 35391 33408 35440 33436
rect 35391 33405 35403 33408
rect 35345 33399 35403 33405
rect 35434 33396 35440 33408
rect 35492 33396 35498 33448
rect 36081 33439 36139 33445
rect 36081 33405 36093 33439
rect 36127 33436 36139 33439
rect 36446 33436 36452 33448
rect 36127 33408 36452 33436
rect 36127 33405 36139 33408
rect 36081 33399 36139 33405
rect 36446 33396 36452 33408
rect 36504 33436 36510 33448
rect 37182 33436 37188 33448
rect 36504 33408 37188 33436
rect 36504 33396 36510 33408
rect 37182 33396 37188 33408
rect 37240 33396 37246 33448
rect 35986 33328 35992 33380
rect 36044 33368 36050 33380
rect 36044 33340 36860 33368
rect 36044 33328 36050 33340
rect 33284 33272 34284 33300
rect 33284 33260 33290 33272
rect 36078 33260 36084 33312
rect 36136 33300 36142 33312
rect 36449 33303 36507 33309
rect 36449 33300 36461 33303
rect 36136 33272 36461 33300
rect 36136 33260 36142 33272
rect 36449 33269 36461 33272
rect 36495 33269 36507 33303
rect 36630 33300 36636 33312
rect 36591 33272 36636 33300
rect 36449 33263 36507 33269
rect 36630 33260 36636 33272
rect 36688 33260 36694 33312
rect 36832 33300 36860 33340
rect 36906 33328 36912 33380
rect 36964 33368 36970 33380
rect 37384 33368 37412 33467
rect 37550 33464 37556 33476
rect 37608 33464 37614 33516
rect 38562 33464 38568 33516
rect 38620 33504 38626 33516
rect 39485 33507 39543 33513
rect 39485 33504 39497 33507
rect 38620 33476 39497 33504
rect 38620 33464 38626 33476
rect 39485 33473 39497 33476
rect 39531 33473 39543 33507
rect 39485 33467 39543 33473
rect 39758 33464 39764 33516
rect 39816 33504 39822 33516
rect 39945 33507 40003 33513
rect 39945 33504 39957 33507
rect 39816 33476 39957 33504
rect 39816 33464 39822 33476
rect 39945 33473 39957 33476
rect 39991 33473 40003 33507
rect 42981 33507 43039 33513
rect 42981 33504 42993 33507
rect 39945 33467 40003 33473
rect 41386 33476 42993 33504
rect 41386 33436 41414 33476
rect 42981 33473 42993 33476
rect 43027 33504 43039 33507
rect 43070 33504 43076 33516
rect 43027 33476 43076 33504
rect 43027 33473 43039 33476
rect 42981 33467 43039 33473
rect 43070 33464 43076 33476
rect 43128 33464 43134 33516
rect 43438 33504 43444 33516
rect 43399 33476 43444 33504
rect 43438 33464 43444 33476
rect 43496 33464 43502 33516
rect 36964 33340 37412 33368
rect 37476 33408 41414 33436
rect 36964 33328 36970 33340
rect 37476 33300 37504 33408
rect 38930 33368 38936 33380
rect 38396 33340 38936 33368
rect 38396 33309 38424 33340
rect 38930 33328 38936 33340
rect 38988 33328 38994 33380
rect 36832 33272 37504 33300
rect 38381 33303 38439 33309
rect 38381 33269 38393 33303
rect 38427 33269 38439 33303
rect 42886 33300 42892 33312
rect 42847 33272 42892 33300
rect 38381 33263 38439 33269
rect 42886 33260 42892 33272
rect 42944 33260 42950 33312
rect 1104 33210 44896 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 44896 33210
rect 1104 33136 44896 33158
rect 16206 33096 16212 33108
rect 16167 33068 16212 33096
rect 16206 33056 16212 33068
rect 16264 33056 16270 33108
rect 19334 33056 19340 33108
rect 19392 33096 19398 33108
rect 19429 33099 19487 33105
rect 19429 33096 19441 33099
rect 19392 33068 19441 33096
rect 19392 33056 19398 33068
rect 19429 33065 19441 33068
rect 19475 33065 19487 33099
rect 19429 33059 19487 33065
rect 23658 33056 23664 33108
rect 23716 33096 23722 33108
rect 23845 33099 23903 33105
rect 23845 33096 23857 33099
rect 23716 33068 23857 33096
rect 23716 33056 23722 33068
rect 23845 33065 23857 33068
rect 23891 33065 23903 33099
rect 26050 33096 26056 33108
rect 26011 33068 26056 33096
rect 23845 33059 23903 33065
rect 26050 33056 26056 33068
rect 26108 33056 26114 33108
rect 32030 33056 32036 33108
rect 32088 33096 32094 33108
rect 32125 33099 32183 33105
rect 32125 33096 32137 33099
rect 32088 33068 32137 33096
rect 32088 33056 32094 33068
rect 32125 33065 32137 33068
rect 32171 33065 32183 33099
rect 32674 33096 32680 33108
rect 32635 33068 32680 33096
rect 32125 33059 32183 33065
rect 32674 33056 32680 33068
rect 32732 33056 32738 33108
rect 34698 33056 34704 33108
rect 34756 33096 34762 33108
rect 35253 33099 35311 33105
rect 35253 33096 35265 33099
rect 34756 33068 35265 33096
rect 34756 33056 34762 33068
rect 35253 33065 35265 33068
rect 35299 33065 35311 33099
rect 35253 33059 35311 33065
rect 35529 33099 35587 33105
rect 35529 33065 35541 33099
rect 35575 33096 35587 33099
rect 36262 33096 36268 33108
rect 35575 33068 36268 33096
rect 35575 33065 35587 33068
rect 35529 33059 35587 33065
rect 36262 33056 36268 33068
rect 36320 33056 36326 33108
rect 36446 33096 36452 33108
rect 36407 33068 36452 33096
rect 36446 33056 36452 33068
rect 36504 33056 36510 33108
rect 36633 33099 36691 33105
rect 36633 33065 36645 33099
rect 36679 33096 36691 33099
rect 37550 33096 37556 33108
rect 36679 33068 37556 33096
rect 36679 33065 36691 33068
rect 36633 33059 36691 33065
rect 37550 33056 37556 33068
rect 37608 33056 37614 33108
rect 13906 32988 13912 33040
rect 13964 33028 13970 33040
rect 19242 33028 19248 33040
rect 13964 33000 19248 33028
rect 13964 32988 13970 33000
rect 19242 32988 19248 33000
rect 19300 32988 19306 33040
rect 27246 33028 27252 33040
rect 27207 33000 27252 33028
rect 27246 32988 27252 33000
rect 27304 32988 27310 33040
rect 27614 32988 27620 33040
rect 27672 33028 27678 33040
rect 28074 33028 28080 33040
rect 27672 33000 28080 33028
rect 27672 32988 27678 33000
rect 28074 32988 28080 33000
rect 28132 32988 28138 33040
rect 33962 32988 33968 33040
rect 34020 33028 34026 33040
rect 34149 33031 34207 33037
rect 34020 33000 34100 33028
rect 34020 32988 34026 33000
rect 15657 32963 15715 32969
rect 15657 32929 15669 32963
rect 15703 32960 15715 32963
rect 16390 32960 16396 32972
rect 15703 32932 16396 32960
rect 15703 32929 15715 32932
rect 15657 32923 15715 32929
rect 16390 32920 16396 32932
rect 16448 32960 16454 32972
rect 17862 32960 17868 32972
rect 16448 32932 16620 32960
rect 17823 32932 17868 32960
rect 16448 32920 16454 32932
rect 15746 32892 15752 32904
rect 15707 32864 15752 32892
rect 15746 32852 15752 32864
rect 15804 32852 15810 32904
rect 16482 32892 16488 32904
rect 16443 32864 16488 32892
rect 16482 32852 16488 32864
rect 16540 32852 16546 32904
rect 16592 32901 16620 32932
rect 17862 32920 17868 32932
rect 17920 32920 17926 32972
rect 17954 32920 17960 32972
rect 18012 32960 18018 32972
rect 18506 32960 18512 32972
rect 18012 32932 18512 32960
rect 18012 32920 18018 32932
rect 16577 32895 16635 32901
rect 16577 32861 16589 32895
rect 16623 32861 16635 32895
rect 16577 32855 16635 32861
rect 16666 32852 16672 32904
rect 16724 32892 16730 32904
rect 18064 32901 18092 32932
rect 18506 32920 18512 32932
rect 18564 32920 18570 32972
rect 27798 32960 27804 32972
rect 26804 32932 27804 32960
rect 16853 32895 16911 32901
rect 16724 32864 16769 32892
rect 16724 32852 16730 32864
rect 16853 32861 16865 32895
rect 16899 32861 16911 32895
rect 16853 32855 16911 32861
rect 18049 32895 18107 32901
rect 18049 32861 18061 32895
rect 18095 32861 18107 32895
rect 18049 32855 18107 32861
rect 16868 32756 16896 32855
rect 18414 32852 18420 32904
rect 18472 32892 18478 32904
rect 19245 32895 19303 32901
rect 19245 32892 19257 32895
rect 18472 32864 19257 32892
rect 18472 32852 18478 32864
rect 19245 32861 19257 32864
rect 19291 32861 19303 32895
rect 19245 32855 19303 32861
rect 19429 32895 19487 32901
rect 19429 32861 19441 32895
rect 19475 32861 19487 32895
rect 19429 32855 19487 32861
rect 18233 32827 18291 32833
rect 18233 32793 18245 32827
rect 18279 32824 18291 32827
rect 19150 32824 19156 32836
rect 18279 32796 19156 32824
rect 18279 32793 18291 32796
rect 18233 32787 18291 32793
rect 19150 32784 19156 32796
rect 19208 32824 19214 32836
rect 19444 32824 19472 32855
rect 21174 32852 21180 32904
rect 21232 32892 21238 32904
rect 22465 32895 22523 32901
rect 22465 32892 22477 32895
rect 21232 32864 22477 32892
rect 21232 32852 21238 32864
rect 22465 32861 22477 32864
rect 22511 32861 22523 32895
rect 22465 32855 22523 32861
rect 24673 32895 24731 32901
rect 24673 32861 24685 32895
rect 24719 32892 24731 32895
rect 25682 32892 25688 32904
rect 24719 32864 25688 32892
rect 24719 32861 24731 32864
rect 24673 32855 24731 32861
rect 25682 32852 25688 32864
rect 25740 32852 25746 32904
rect 26804 32901 26832 32932
rect 27798 32920 27804 32932
rect 27856 32920 27862 32972
rect 32033 32963 32091 32969
rect 32033 32929 32045 32963
rect 32079 32960 32091 32963
rect 32122 32960 32128 32972
rect 32079 32932 32128 32960
rect 32079 32929 32091 32932
rect 32033 32923 32091 32929
rect 32122 32920 32128 32932
rect 32180 32920 32186 32972
rect 32217 32963 32275 32969
rect 32217 32929 32229 32963
rect 32263 32960 32275 32963
rect 33226 32960 33232 32972
rect 32263 32932 33232 32960
rect 32263 32929 32275 32932
rect 32217 32923 32275 32929
rect 33226 32920 33232 32932
rect 33284 32920 33290 32972
rect 34072 32960 34100 33000
rect 34149 32997 34161 33031
rect 34195 33028 34207 33031
rect 35342 33028 35348 33040
rect 34195 33000 35348 33028
rect 34195 32997 34207 33000
rect 34149 32991 34207 32997
rect 35342 32988 35348 33000
rect 35400 33028 35406 33040
rect 35894 33028 35900 33040
rect 35400 33000 35900 33028
rect 35400 32988 35406 33000
rect 35894 32988 35900 33000
rect 35952 32988 35958 33040
rect 36354 32988 36360 33040
rect 36412 33028 36418 33040
rect 37277 33031 37335 33037
rect 37277 33028 37289 33031
rect 36412 33000 37289 33028
rect 36412 32988 36418 33000
rect 37277 32997 37289 33000
rect 37323 32997 37335 33031
rect 37277 32991 37335 32997
rect 38654 32960 38660 32972
rect 34072 32932 35848 32960
rect 38615 32932 38660 32960
rect 26789 32895 26847 32901
rect 26789 32861 26801 32895
rect 26835 32861 26847 32895
rect 26789 32855 26847 32861
rect 27065 32895 27123 32901
rect 27065 32861 27077 32895
rect 27111 32892 27123 32895
rect 27614 32892 27620 32904
rect 27111 32864 27620 32892
rect 27111 32861 27123 32864
rect 27065 32855 27123 32861
rect 27614 32852 27620 32864
rect 27672 32852 27678 32904
rect 27706 32852 27712 32904
rect 27764 32892 27770 32904
rect 27890 32892 27896 32904
rect 27764 32864 27809 32892
rect 27851 32864 27896 32892
rect 27764 32852 27770 32864
rect 27890 32852 27896 32864
rect 27948 32852 27954 32904
rect 27985 32895 28043 32901
rect 27985 32861 27997 32895
rect 28031 32861 28043 32895
rect 27985 32855 28043 32861
rect 28077 32895 28135 32901
rect 28077 32861 28089 32895
rect 28123 32892 28135 32895
rect 28350 32892 28356 32904
rect 28123 32864 28356 32892
rect 28123 32861 28135 32864
rect 28077 32855 28135 32861
rect 19208 32796 19472 32824
rect 22732 32827 22790 32833
rect 19208 32784 19214 32796
rect 22732 32793 22744 32827
rect 22778 32824 22790 32827
rect 22830 32824 22836 32836
rect 22778 32796 22836 32824
rect 22778 32793 22790 32796
rect 22732 32787 22790 32793
rect 22830 32784 22836 32796
rect 22888 32784 22894 32836
rect 24946 32833 24952 32836
rect 24940 32787 24952 32833
rect 25004 32824 25010 32836
rect 25004 32796 25040 32824
rect 24946 32784 24952 32787
rect 25004 32784 25010 32796
rect 27338 32784 27344 32836
rect 27396 32824 27402 32836
rect 28000 32824 28028 32855
rect 28350 32852 28356 32864
rect 28408 32852 28414 32904
rect 31938 32892 31944 32904
rect 31899 32864 31944 32892
rect 31938 32852 31944 32864
rect 31996 32852 32002 32904
rect 32306 32852 32312 32904
rect 32364 32892 32370 32904
rect 32677 32895 32735 32901
rect 32677 32892 32689 32895
rect 32364 32864 32689 32892
rect 32364 32852 32370 32864
rect 32677 32861 32689 32864
rect 32723 32861 32735 32895
rect 32677 32855 32735 32861
rect 32861 32895 32919 32901
rect 32861 32861 32873 32895
rect 32907 32892 32919 32895
rect 33042 32892 33048 32904
rect 32907 32864 33048 32892
rect 32907 32861 32919 32864
rect 32861 32855 32919 32861
rect 33042 32852 33048 32864
rect 33100 32852 33106 32904
rect 33134 32852 33140 32904
rect 33192 32892 33198 32904
rect 33965 32895 34023 32901
rect 33965 32892 33977 32895
rect 33192 32864 33977 32892
rect 33192 32852 33198 32864
rect 33965 32861 33977 32864
rect 34011 32861 34023 32895
rect 33965 32855 34023 32861
rect 35437 32895 35495 32901
rect 35437 32861 35449 32895
rect 35483 32892 35495 32895
rect 35710 32892 35716 32904
rect 35483 32864 35716 32892
rect 35483 32861 35495 32864
rect 35437 32855 35495 32861
rect 35710 32852 35716 32864
rect 35768 32852 35774 32904
rect 35820 32901 35848 32932
rect 38654 32920 38660 32932
rect 38712 32920 38718 32972
rect 42521 32963 42579 32969
rect 42521 32929 42533 32963
rect 42567 32960 42579 32963
rect 42886 32960 42892 32972
rect 42567 32932 42892 32960
rect 42567 32929 42579 32932
rect 42521 32923 42579 32929
rect 42886 32920 42892 32932
rect 42944 32920 42950 32972
rect 44082 32960 44088 32972
rect 44043 32932 44088 32960
rect 44082 32920 44088 32932
rect 44140 32920 44146 32972
rect 35805 32895 35863 32901
rect 35805 32861 35817 32895
rect 35851 32861 35863 32895
rect 35805 32855 35863 32861
rect 35897 32895 35955 32901
rect 35897 32861 35909 32895
rect 35943 32892 35955 32895
rect 36354 32892 36360 32904
rect 35943 32864 36360 32892
rect 35943 32861 35955 32864
rect 35897 32855 35955 32861
rect 36354 32852 36360 32864
rect 36412 32852 36418 32904
rect 39114 32892 39120 32904
rect 39075 32864 39120 32892
rect 39114 32852 39120 32864
rect 39172 32852 39178 32904
rect 42334 32892 42340 32904
rect 42295 32864 42340 32892
rect 42334 32852 42340 32864
rect 42392 32852 42398 32904
rect 30926 32824 30932 32836
rect 27396 32796 28028 32824
rect 28092 32796 30932 32824
rect 27396 32784 27402 32796
rect 19426 32756 19432 32768
rect 16868 32728 19432 32756
rect 19426 32716 19432 32728
rect 19484 32716 19490 32768
rect 21358 32716 21364 32768
rect 21416 32756 21422 32768
rect 23842 32756 23848 32768
rect 21416 32728 23848 32756
rect 21416 32716 21422 32728
rect 23842 32716 23848 32728
rect 23900 32716 23906 32768
rect 26878 32756 26884 32768
rect 26839 32728 26884 32756
rect 26878 32716 26884 32728
rect 26936 32716 26942 32768
rect 27706 32716 27712 32768
rect 27764 32756 27770 32768
rect 28092 32756 28120 32796
rect 30926 32784 30932 32796
rect 30984 32784 30990 32836
rect 35526 32784 35532 32836
rect 35584 32824 35590 32836
rect 36601 32827 36659 32833
rect 36601 32824 36613 32827
rect 35584 32796 36613 32824
rect 35584 32784 35590 32796
rect 36601 32793 36613 32796
rect 36647 32793 36659 32827
rect 36601 32787 36659 32793
rect 36817 32827 36875 32833
rect 36817 32793 36829 32827
rect 36863 32824 36875 32827
rect 36906 32824 36912 32836
rect 36863 32796 36912 32824
rect 36863 32793 36875 32796
rect 36817 32787 36875 32793
rect 36906 32784 36912 32796
rect 36964 32784 36970 32836
rect 37366 32784 37372 32836
rect 37424 32824 37430 32836
rect 38390 32827 38448 32833
rect 38390 32824 38402 32827
rect 37424 32796 38402 32824
rect 37424 32784 37430 32796
rect 38390 32793 38402 32796
rect 38436 32793 38448 32827
rect 38390 32787 38448 32793
rect 28350 32756 28356 32768
rect 27764 32728 28120 32756
rect 28311 32728 28356 32756
rect 27764 32716 27770 32728
rect 28350 32716 28356 32728
rect 28408 32716 28414 32768
rect 39301 32759 39359 32765
rect 39301 32725 39313 32759
rect 39347 32756 39359 32759
rect 39942 32756 39948 32768
rect 39347 32728 39948 32756
rect 39347 32725 39359 32728
rect 39301 32719 39359 32725
rect 39942 32716 39948 32728
rect 40000 32716 40006 32768
rect 1104 32666 44896 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 44896 32666
rect 1104 32592 44896 32614
rect 16758 32552 16764 32564
rect 16224 32524 16764 32552
rect 16224 32484 16252 32524
rect 16758 32512 16764 32524
rect 16816 32512 16822 32564
rect 17880 32524 20760 32552
rect 16132 32456 16252 32484
rect 15562 32416 15568 32428
rect 15523 32388 15568 32416
rect 15562 32376 15568 32388
rect 15620 32376 15626 32428
rect 15930 32416 15936 32428
rect 15891 32388 15936 32416
rect 15930 32376 15936 32388
rect 15988 32376 15994 32428
rect 16132 32425 16160 32456
rect 16390 32444 16396 32496
rect 16448 32484 16454 32496
rect 17880 32493 17908 32524
rect 17865 32487 17923 32493
rect 17865 32484 17877 32487
rect 16448 32456 17877 32484
rect 16448 32444 16454 32456
rect 17865 32453 17877 32456
rect 17911 32453 17923 32487
rect 19426 32484 19432 32496
rect 17865 32447 17923 32453
rect 18984 32456 19432 32484
rect 16117 32419 16175 32425
rect 16117 32385 16129 32419
rect 16163 32385 16175 32419
rect 16117 32379 16175 32385
rect 16206 32376 16212 32428
rect 16264 32416 16270 32428
rect 16853 32419 16911 32425
rect 16853 32416 16865 32419
rect 16264 32388 16865 32416
rect 16264 32376 16270 32388
rect 16853 32385 16865 32388
rect 16899 32416 16911 32419
rect 16899 32388 18092 32416
rect 16899 32385 16911 32388
rect 16853 32379 16911 32385
rect 15749 32351 15807 32357
rect 15749 32317 15761 32351
rect 15795 32317 15807 32351
rect 15749 32311 15807 32317
rect 15841 32351 15899 32357
rect 15841 32317 15853 32351
rect 15887 32348 15899 32351
rect 16022 32348 16028 32360
rect 15887 32320 16028 32348
rect 15887 32317 15899 32320
rect 15841 32311 15899 32317
rect 15764 32280 15792 32311
rect 16022 32308 16028 32320
rect 16080 32348 16086 32360
rect 16390 32348 16396 32360
rect 16080 32320 16396 32348
rect 16080 32308 16086 32320
rect 16390 32308 16396 32320
rect 16448 32308 16454 32360
rect 16482 32308 16488 32360
rect 16540 32348 16546 32360
rect 17037 32351 17095 32357
rect 17037 32348 17049 32351
rect 16540 32320 17049 32348
rect 16540 32308 16546 32320
rect 17037 32317 17049 32320
rect 17083 32317 17095 32351
rect 17037 32311 17095 32317
rect 17957 32351 18015 32357
rect 17957 32317 17969 32351
rect 18003 32317 18015 32351
rect 18064 32348 18092 32388
rect 18138 32376 18144 32428
rect 18196 32416 18202 32428
rect 18233 32419 18291 32425
rect 18233 32416 18245 32419
rect 18196 32388 18245 32416
rect 18196 32376 18202 32388
rect 18233 32385 18245 32388
rect 18279 32416 18291 32419
rect 18414 32416 18420 32428
rect 18279 32388 18420 32416
rect 18279 32385 18291 32388
rect 18233 32379 18291 32385
rect 18414 32376 18420 32388
rect 18472 32376 18478 32428
rect 18984 32425 19012 32456
rect 19426 32444 19432 32456
rect 19484 32484 19490 32496
rect 20622 32484 20628 32496
rect 19484 32456 20628 32484
rect 19484 32444 19490 32456
rect 20622 32444 20628 32456
rect 20680 32444 20686 32496
rect 18969 32419 19027 32425
rect 18969 32385 18981 32419
rect 19015 32385 19027 32419
rect 19153 32419 19211 32425
rect 19153 32417 19165 32419
rect 18969 32379 19027 32385
rect 19076 32389 19165 32417
rect 18322 32348 18328 32360
rect 18064 32320 18328 32348
rect 17957 32311 18015 32317
rect 16669 32283 16727 32289
rect 16669 32280 16681 32283
rect 15764 32252 16681 32280
rect 16669 32249 16681 32252
rect 16715 32249 16727 32283
rect 16669 32243 16727 32249
rect 14366 32172 14372 32224
rect 14424 32212 14430 32224
rect 15381 32215 15439 32221
rect 15381 32212 15393 32215
rect 14424 32184 15393 32212
rect 14424 32172 14430 32184
rect 15381 32181 15393 32184
rect 15427 32181 15439 32215
rect 15381 32175 15439 32181
rect 16206 32172 16212 32224
rect 16264 32212 16270 32224
rect 16758 32212 16764 32224
rect 16264 32184 16764 32212
rect 16264 32172 16270 32184
rect 16758 32172 16764 32184
rect 16816 32172 16822 32224
rect 17972 32212 18000 32311
rect 18322 32308 18328 32320
rect 18380 32308 18386 32360
rect 19076 32348 19104 32389
rect 19153 32385 19165 32389
rect 19199 32385 19211 32419
rect 19153 32379 19211 32385
rect 19245 32419 19303 32425
rect 19245 32385 19257 32419
rect 19291 32385 19303 32419
rect 19245 32379 19303 32385
rect 19337 32419 19395 32425
rect 19337 32385 19349 32419
rect 19383 32385 19395 32419
rect 19337 32379 19395 32385
rect 18524 32320 19104 32348
rect 18524 32289 18552 32320
rect 18509 32283 18567 32289
rect 18509 32249 18521 32283
rect 18555 32249 18567 32283
rect 18509 32243 18567 32249
rect 19150 32240 19156 32292
rect 19208 32280 19214 32292
rect 19260 32280 19288 32379
rect 19208 32252 19288 32280
rect 19208 32240 19214 32252
rect 18966 32212 18972 32224
rect 17972 32184 18972 32212
rect 18966 32172 18972 32184
rect 19024 32212 19030 32224
rect 19352 32212 19380 32379
rect 20732 32348 20760 32524
rect 21266 32512 21272 32564
rect 21324 32512 21330 32564
rect 22830 32552 22836 32564
rect 22791 32524 22836 32552
rect 22830 32512 22836 32524
rect 22888 32512 22894 32564
rect 24946 32552 24952 32564
rect 24907 32524 24952 32552
rect 24946 32512 24952 32524
rect 25004 32512 25010 32564
rect 26878 32552 26884 32564
rect 25332 32524 26884 32552
rect 21284 32484 21312 32512
rect 21100 32456 21312 32484
rect 21100 32425 21128 32456
rect 22738 32444 22744 32496
rect 22796 32484 22802 32496
rect 23661 32487 23719 32493
rect 23661 32484 23673 32487
rect 22796 32456 23673 32484
rect 22796 32444 22802 32456
rect 23661 32453 23673 32456
rect 23707 32453 23719 32487
rect 23661 32447 23719 32453
rect 24397 32487 24455 32493
rect 24397 32453 24409 32487
rect 24443 32484 24455 32487
rect 24486 32484 24492 32496
rect 24443 32456 24492 32484
rect 24443 32453 24455 32456
rect 24397 32447 24455 32453
rect 24486 32444 24492 32456
rect 24544 32444 24550 32496
rect 25332 32431 25360 32524
rect 26878 32512 26884 32524
rect 26936 32552 26942 32564
rect 27341 32555 27399 32561
rect 27341 32552 27353 32555
rect 26936 32524 27353 32552
rect 26936 32512 26942 32524
rect 27341 32521 27353 32524
rect 27387 32552 27399 32555
rect 27982 32552 27988 32564
rect 27387 32524 27988 32552
rect 27387 32521 27399 32524
rect 27341 32515 27399 32521
rect 27982 32512 27988 32524
rect 28040 32512 28046 32564
rect 28626 32552 28632 32564
rect 28587 32524 28632 32552
rect 28626 32512 28632 32524
rect 28684 32512 28690 32564
rect 33413 32555 33471 32561
rect 33413 32521 33425 32555
rect 33459 32552 33471 32555
rect 33962 32552 33968 32564
rect 33459 32524 33968 32552
rect 33459 32521 33471 32524
rect 33413 32515 33471 32521
rect 33962 32512 33968 32524
rect 34020 32512 34026 32564
rect 35437 32555 35495 32561
rect 35437 32521 35449 32555
rect 35483 32552 35495 32555
rect 36173 32555 36231 32561
rect 36173 32552 36185 32555
rect 35483 32524 36185 32552
rect 35483 32521 35495 32524
rect 35437 32515 35495 32521
rect 36173 32521 36185 32524
rect 36219 32552 36231 32555
rect 36906 32552 36912 32564
rect 36219 32524 36912 32552
rect 36219 32521 36231 32524
rect 36173 32515 36231 32521
rect 36906 32512 36912 32524
rect 36964 32512 36970 32564
rect 37366 32552 37372 32564
rect 37327 32524 37372 32552
rect 37366 32512 37372 32524
rect 37424 32512 37430 32564
rect 38841 32555 38899 32561
rect 38841 32521 38853 32555
rect 38887 32552 38899 32555
rect 38930 32552 38936 32564
rect 38887 32524 38936 32552
rect 38887 32521 38899 32524
rect 38841 32515 38899 32521
rect 38930 32512 38936 32524
rect 38988 32512 38994 32564
rect 27062 32484 27068 32496
rect 25424 32456 27068 32484
rect 21085 32419 21143 32425
rect 21085 32385 21097 32419
rect 21131 32385 21143 32419
rect 21085 32379 21143 32385
rect 21269 32419 21327 32425
rect 21269 32385 21281 32419
rect 21315 32416 21327 32419
rect 21358 32416 21364 32428
rect 21315 32388 21364 32416
rect 21315 32385 21327 32388
rect 21269 32379 21327 32385
rect 21358 32376 21364 32388
rect 21416 32376 21422 32428
rect 22189 32419 22247 32425
rect 22189 32385 22201 32419
rect 22235 32385 22247 32419
rect 22370 32416 22376 32428
rect 22331 32388 22376 32416
rect 22189 32379 22247 32385
rect 22204 32348 22232 32379
rect 22370 32376 22376 32388
rect 22428 32376 22434 32428
rect 22465 32419 22523 32425
rect 22465 32385 22477 32419
rect 22511 32385 22523 32419
rect 22465 32379 22523 32385
rect 22557 32419 22615 32425
rect 22557 32385 22569 32419
rect 22603 32416 22615 32419
rect 23198 32416 23204 32428
rect 22603 32388 23204 32416
rect 22603 32385 22615 32388
rect 22557 32379 22615 32385
rect 22278 32348 22284 32360
rect 20732 32320 22094 32348
rect 22204 32320 22284 32348
rect 22066 32280 22094 32320
rect 22278 32308 22284 32320
rect 22336 32308 22342 32360
rect 22480 32348 22508 32379
rect 23198 32376 23204 32388
rect 23256 32376 23262 32428
rect 23477 32419 23535 32425
rect 23477 32416 23489 32419
rect 23400 32388 23489 32416
rect 23290 32348 23296 32360
rect 22480 32320 23296 32348
rect 23290 32308 23296 32320
rect 23348 32308 23354 32360
rect 23400 32348 23428 32388
rect 23477 32385 23489 32388
rect 23523 32385 23535 32419
rect 23477 32379 23535 32385
rect 23753 32419 23811 32425
rect 23753 32385 23765 32419
rect 23799 32416 23811 32419
rect 24670 32416 24676 32428
rect 23799 32388 24676 32416
rect 23799 32385 23811 32388
rect 23753 32379 23811 32385
rect 24670 32376 24676 32388
rect 24728 32376 24734 32428
rect 25314 32425 25372 32431
rect 25424 32428 25452 32456
rect 27062 32444 27068 32456
rect 27120 32444 27126 32496
rect 27706 32484 27712 32496
rect 27264 32456 27712 32484
rect 25225 32419 25283 32425
rect 25225 32385 25237 32419
rect 25271 32385 25283 32419
rect 25314 32391 25326 32425
rect 25360 32391 25372 32425
rect 25314 32385 25372 32391
rect 25409 32422 25467 32428
rect 25409 32388 25421 32422
rect 25455 32388 25467 32422
rect 25225 32379 25283 32385
rect 25409 32382 25467 32388
rect 25593 32419 25651 32425
rect 25593 32385 25605 32419
rect 25639 32416 25651 32419
rect 26237 32419 26295 32425
rect 25639 32388 26188 32416
rect 25639 32385 25651 32388
rect 25593 32379 25651 32385
rect 25130 32348 25136 32360
rect 23400 32320 25136 32348
rect 23400 32280 23428 32320
rect 25130 32308 25136 32320
rect 25188 32308 25194 32360
rect 25240 32348 25268 32379
rect 26050 32348 26056 32360
rect 25240 32320 26056 32348
rect 26050 32308 26056 32320
rect 26108 32308 26114 32360
rect 26160 32348 26188 32388
rect 26237 32385 26249 32419
rect 26283 32416 26295 32419
rect 26326 32416 26332 32428
rect 26283 32388 26332 32416
rect 26283 32385 26295 32388
rect 26237 32379 26295 32385
rect 26326 32376 26332 32388
rect 26384 32376 26390 32428
rect 26878 32376 26884 32428
rect 26936 32416 26942 32428
rect 27157 32419 27215 32425
rect 27157 32416 27169 32419
rect 26936 32388 27169 32416
rect 26936 32376 26942 32388
rect 27157 32385 27169 32388
rect 27203 32385 27215 32419
rect 27157 32379 27215 32385
rect 27264 32348 27292 32456
rect 27706 32444 27712 32456
rect 27764 32444 27770 32496
rect 28350 32444 28356 32496
rect 28408 32484 28414 32496
rect 29742 32487 29800 32493
rect 29742 32484 29754 32487
rect 28408 32456 29754 32484
rect 28408 32444 28414 32456
rect 29742 32453 29754 32456
rect 29788 32453 29800 32487
rect 29742 32447 29800 32453
rect 34548 32487 34606 32493
rect 34548 32453 34560 32487
rect 34594 32484 34606 32487
rect 34790 32484 34796 32496
rect 34594 32456 34796 32484
rect 34594 32453 34606 32456
rect 34548 32447 34606 32453
rect 34790 32444 34796 32456
rect 34848 32444 34854 32496
rect 35253 32487 35311 32493
rect 35253 32453 35265 32487
rect 35299 32484 35311 32487
rect 35618 32484 35624 32496
rect 35299 32456 35624 32484
rect 35299 32453 35311 32456
rect 35253 32447 35311 32453
rect 35618 32444 35624 32456
rect 35676 32444 35682 32496
rect 36078 32444 36084 32496
rect 36136 32484 36142 32496
rect 36136 32456 40264 32484
rect 36136 32444 36142 32456
rect 27433 32419 27491 32425
rect 27433 32385 27445 32419
rect 27479 32385 27491 32419
rect 27433 32379 27491 32385
rect 26160 32320 27292 32348
rect 27448 32348 27476 32379
rect 27798 32376 27804 32428
rect 27856 32416 27862 32428
rect 27893 32419 27951 32425
rect 27893 32416 27905 32419
rect 27856 32388 27905 32416
rect 27856 32376 27862 32388
rect 27893 32385 27905 32388
rect 27939 32385 27951 32419
rect 28074 32416 28080 32428
rect 28035 32388 28080 32416
rect 27893 32379 27951 32385
rect 28074 32376 28080 32388
rect 28132 32376 28138 32428
rect 30650 32416 30656 32428
rect 30611 32388 30656 32416
rect 30650 32376 30656 32388
rect 30708 32376 30714 32428
rect 35526 32416 35532 32428
rect 35487 32388 35532 32416
rect 35526 32376 35532 32388
rect 35584 32376 35590 32428
rect 35710 32376 35716 32428
rect 35768 32416 35774 32428
rect 35989 32419 36047 32425
rect 35989 32416 36001 32419
rect 35768 32388 36001 32416
rect 35768 32376 35774 32388
rect 35989 32385 36001 32388
rect 36035 32385 36047 32419
rect 37274 32416 37280 32428
rect 37235 32388 37280 32416
rect 35989 32379 36047 32385
rect 37274 32376 37280 32388
rect 37332 32376 37338 32428
rect 37461 32419 37519 32425
rect 37461 32385 37473 32419
rect 37507 32416 37519 32419
rect 38378 32416 38384 32428
rect 37507 32388 38384 32416
rect 37507 32385 37519 32388
rect 37461 32379 37519 32385
rect 38378 32376 38384 32388
rect 38436 32376 38442 32428
rect 39942 32376 39948 32428
rect 40000 32425 40006 32428
rect 40236 32425 40264 32456
rect 40000 32416 40012 32425
rect 40221 32419 40279 32425
rect 40000 32388 40045 32416
rect 40000 32379 40012 32388
rect 40221 32385 40233 32419
rect 40267 32385 40279 32419
rect 40221 32379 40279 32385
rect 40000 32376 40006 32379
rect 42334 32376 42340 32428
rect 42392 32416 42398 32428
rect 43625 32419 43683 32425
rect 43625 32416 43637 32419
rect 42392 32388 43637 32416
rect 42392 32376 42398 32388
rect 43625 32385 43637 32388
rect 43671 32385 43683 32419
rect 43625 32379 43683 32385
rect 27985 32351 28043 32357
rect 27985 32348 27997 32351
rect 27448 32320 27997 32348
rect 24210 32280 24216 32292
rect 22066 32252 23428 32280
rect 24171 32252 24216 32280
rect 24210 32240 24216 32252
rect 24268 32240 24274 32292
rect 19024 32184 19380 32212
rect 19613 32215 19671 32221
rect 19024 32172 19030 32184
rect 19613 32181 19625 32215
rect 19659 32212 19671 32215
rect 20346 32212 20352 32224
rect 19659 32184 20352 32212
rect 19659 32181 19671 32184
rect 19613 32175 19671 32181
rect 20346 32172 20352 32184
rect 20404 32172 20410 32224
rect 20714 32172 20720 32224
rect 20772 32212 20778 32224
rect 21177 32215 21235 32221
rect 21177 32212 21189 32215
rect 20772 32184 21189 32212
rect 20772 32172 20778 32184
rect 21177 32181 21189 32184
rect 21223 32181 21235 32215
rect 21177 32175 21235 32181
rect 22094 32172 22100 32224
rect 22152 32212 22158 32224
rect 22278 32212 22284 32224
rect 22152 32184 22284 32212
rect 22152 32172 22158 32184
rect 22278 32172 22284 32184
rect 22336 32212 22342 32224
rect 26160 32212 26188 32320
rect 27985 32317 27997 32320
rect 28031 32317 28043 32351
rect 27985 32311 28043 32317
rect 30009 32351 30067 32357
rect 30009 32317 30021 32351
rect 30055 32348 30067 32351
rect 31754 32348 31760 32360
rect 30055 32320 31760 32348
rect 30055 32317 30067 32320
rect 30009 32311 30067 32317
rect 31754 32308 31760 32320
rect 31812 32308 31818 32360
rect 34790 32348 34796 32360
rect 34751 32320 34796 32348
rect 34790 32308 34796 32320
rect 34848 32308 34854 32360
rect 26970 32280 26976 32292
rect 26883 32252 26976 32280
rect 26970 32240 26976 32252
rect 27028 32280 27034 32292
rect 27338 32280 27344 32292
rect 27028 32252 27344 32280
rect 27028 32240 27034 32252
rect 27338 32240 27344 32252
rect 27396 32240 27402 32292
rect 30466 32280 30472 32292
rect 30427 32252 30472 32280
rect 30466 32240 30472 32252
rect 30524 32240 30530 32292
rect 26418 32212 26424 32224
rect 22336 32184 26188 32212
rect 26379 32184 26424 32212
rect 22336 32172 22342 32184
rect 26418 32172 26424 32184
rect 26476 32172 26482 32224
rect 35253 32215 35311 32221
rect 35253 32181 35265 32215
rect 35299 32212 35311 32215
rect 35434 32212 35440 32224
rect 35299 32184 35440 32212
rect 35299 32181 35311 32184
rect 35253 32175 35311 32181
rect 35434 32172 35440 32184
rect 35492 32172 35498 32224
rect 1104 32122 44896 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 44896 32122
rect 1104 32048 44896 32070
rect 16666 32008 16672 32020
rect 15488 31980 16672 32008
rect 15488 31949 15516 31980
rect 16666 31968 16672 31980
rect 16724 31968 16730 32020
rect 17862 31968 17868 32020
rect 17920 32008 17926 32020
rect 18509 32011 18567 32017
rect 18509 32008 18521 32011
rect 17920 31980 18521 32008
rect 17920 31968 17926 31980
rect 18509 31977 18521 31980
rect 18555 31977 18567 32011
rect 18509 31971 18567 31977
rect 22649 32011 22707 32017
rect 22649 31977 22661 32011
rect 22695 32008 22707 32011
rect 23293 32011 23351 32017
rect 23293 32008 23305 32011
rect 22695 31980 23305 32008
rect 22695 31977 22707 31980
rect 22649 31971 22707 31977
rect 23293 31977 23305 31980
rect 23339 31977 23351 32011
rect 24670 32008 24676 32020
rect 23293 31971 23351 31977
rect 23400 31980 24348 32008
rect 24631 31980 24676 32008
rect 15473 31943 15531 31949
rect 15473 31909 15485 31943
rect 15519 31909 15531 31943
rect 15473 31903 15531 31909
rect 15562 31900 15568 31952
rect 15620 31940 15626 31952
rect 18322 31940 18328 31952
rect 15620 31912 16344 31940
rect 18283 31912 18328 31940
rect 15620 31900 15626 31912
rect 16114 31832 16120 31884
rect 16172 31872 16178 31884
rect 16316 31881 16344 31912
rect 18322 31900 18328 31912
rect 18380 31900 18386 31952
rect 22186 31900 22192 31952
rect 22244 31940 22250 31952
rect 23400 31940 23428 31980
rect 22244 31912 23428 31940
rect 22244 31900 22250 31912
rect 16301 31875 16359 31881
rect 16172 31844 16217 31872
rect 16172 31832 16178 31844
rect 16301 31841 16313 31875
rect 16347 31841 16359 31875
rect 24210 31872 24216 31884
rect 16301 31835 16359 31841
rect 22066 31844 24216 31872
rect 13906 31764 13912 31816
rect 13964 31804 13970 31816
rect 14093 31807 14151 31813
rect 14093 31804 14105 31807
rect 13964 31776 14105 31804
rect 13964 31764 13970 31776
rect 14093 31773 14105 31776
rect 14139 31773 14151 31807
rect 14093 31767 14151 31773
rect 16209 31807 16267 31813
rect 16209 31773 16221 31807
rect 16255 31804 16267 31807
rect 16393 31807 16451 31813
rect 16255 31776 16289 31804
rect 16255 31773 16267 31776
rect 16209 31767 16267 31773
rect 16393 31773 16405 31807
rect 16439 31804 16451 31807
rect 16482 31804 16488 31816
rect 16439 31776 16488 31804
rect 16439 31773 16451 31776
rect 16393 31767 16451 31773
rect 14366 31745 14372 31748
rect 14360 31699 14372 31745
rect 14424 31736 14430 31748
rect 16224 31736 16252 31767
rect 16482 31764 16488 31776
rect 16540 31804 16546 31816
rect 17037 31807 17095 31813
rect 17037 31804 17049 31807
rect 16540 31776 17049 31804
rect 16540 31764 16546 31776
rect 17037 31773 17049 31776
rect 17083 31773 17095 31807
rect 17037 31767 17095 31773
rect 17313 31807 17371 31813
rect 17313 31773 17325 31807
rect 17359 31804 17371 31807
rect 17589 31807 17647 31813
rect 17359 31776 17393 31804
rect 17359 31773 17371 31776
rect 17313 31767 17371 31773
rect 17589 31773 17601 31807
rect 17635 31804 17647 31807
rect 17770 31804 17776 31816
rect 17635 31776 17669 31804
rect 17731 31776 17776 31804
rect 17635 31773 17647 31776
rect 17589 31767 17647 31773
rect 16574 31736 16580 31748
rect 14424 31708 14460 31736
rect 16224 31708 16580 31736
rect 14366 31696 14372 31699
rect 14424 31696 14430 31708
rect 16574 31696 16580 31708
rect 16632 31696 16638 31748
rect 16666 31696 16672 31748
rect 16724 31736 16730 31748
rect 17328 31736 17356 31767
rect 16724 31708 17356 31736
rect 17604 31736 17632 31767
rect 17770 31764 17776 31776
rect 17828 31764 17834 31816
rect 19242 31764 19248 31816
rect 19300 31804 19306 31816
rect 20625 31807 20683 31813
rect 20625 31804 20637 31807
rect 19300 31776 20637 31804
rect 19300 31764 19306 31776
rect 20625 31773 20637 31776
rect 20671 31804 20683 31807
rect 21174 31804 21180 31816
rect 20671 31776 21180 31804
rect 20671 31773 20683 31776
rect 20625 31767 20683 31773
rect 21174 31764 21180 31776
rect 21232 31764 21238 31816
rect 21361 31807 21419 31813
rect 21361 31773 21373 31807
rect 21407 31804 21419 31807
rect 22066 31804 22094 31844
rect 24210 31832 24216 31844
rect 24268 31832 24274 31884
rect 24320 31872 24348 31980
rect 24670 31968 24676 31980
rect 24728 31968 24734 32020
rect 25130 31968 25136 32020
rect 25188 32008 25194 32020
rect 25869 32011 25927 32017
rect 25869 32008 25881 32011
rect 25188 31980 25881 32008
rect 25188 31968 25194 31980
rect 25869 31977 25881 31980
rect 25915 32008 25927 32011
rect 26878 32008 26884 32020
rect 25915 31980 26884 32008
rect 25915 31977 25927 31980
rect 25869 31971 25927 31977
rect 26878 31968 26884 31980
rect 26936 31968 26942 32020
rect 28166 31968 28172 32020
rect 28224 32008 28230 32020
rect 28629 32011 28687 32017
rect 28629 32008 28641 32011
rect 28224 31980 28641 32008
rect 28224 31968 28230 31980
rect 28629 31977 28641 31980
rect 28675 31977 28687 32011
rect 28629 31971 28687 31977
rect 35710 31968 35716 32020
rect 35768 32008 35774 32020
rect 36173 32011 36231 32017
rect 36173 32008 36185 32011
rect 35768 31980 36185 32008
rect 35768 31968 35774 31980
rect 36173 31977 36185 31980
rect 36219 31977 36231 32011
rect 36173 31971 36231 31977
rect 29825 31943 29883 31949
rect 29825 31909 29837 31943
rect 29871 31940 29883 31943
rect 30374 31940 30380 31952
rect 29871 31912 30380 31940
rect 29871 31909 29883 31912
rect 29825 31903 29883 31909
rect 30374 31900 30380 31912
rect 30432 31940 30438 31952
rect 30650 31940 30656 31952
rect 30432 31912 30656 31940
rect 30432 31900 30438 31912
rect 30650 31900 30656 31912
rect 30708 31900 30714 31952
rect 24320 31844 24808 31872
rect 21407 31776 22094 31804
rect 21407 31773 21419 31776
rect 21361 31767 21419 31773
rect 22186 31764 22192 31816
rect 22244 31804 22250 31816
rect 22462 31804 22468 31816
rect 22244 31776 22289 31804
rect 22423 31776 22468 31804
rect 22244 31764 22250 31776
rect 22462 31764 22468 31776
rect 22520 31764 22526 31816
rect 23382 31764 23388 31816
rect 23440 31804 23446 31816
rect 24780 31813 24808 31844
rect 25682 31832 25688 31884
rect 25740 31872 25746 31884
rect 27249 31875 27307 31881
rect 27249 31872 27261 31875
rect 25740 31844 27261 31872
rect 25740 31832 25746 31844
rect 27249 31841 27261 31844
rect 27295 31841 27307 31875
rect 32122 31872 32128 31884
rect 27249 31835 27307 31841
rect 31588 31844 32128 31872
rect 24581 31807 24639 31813
rect 24581 31804 24593 31807
rect 23440 31776 24593 31804
rect 23440 31764 23446 31776
rect 24581 31773 24593 31776
rect 24627 31773 24639 31807
rect 24581 31767 24639 31773
rect 24765 31807 24823 31813
rect 24765 31773 24777 31807
rect 24811 31773 24823 31807
rect 24765 31767 24823 31773
rect 25038 31764 25044 31816
rect 25096 31804 25102 31816
rect 25096 31776 25636 31804
rect 25096 31764 25102 31776
rect 18693 31739 18751 31745
rect 17604 31708 18644 31736
rect 16724 31696 16730 31708
rect 15930 31668 15936 31680
rect 15891 31640 15936 31668
rect 15930 31628 15936 31640
rect 15988 31628 15994 31680
rect 17494 31628 17500 31680
rect 17552 31668 17558 31680
rect 18506 31677 18512 31680
rect 17589 31671 17647 31677
rect 17589 31668 17601 31671
rect 17552 31640 17601 31668
rect 17552 31628 17558 31640
rect 17589 31637 17601 31640
rect 17635 31637 17647 31671
rect 17589 31631 17647 31637
rect 18493 31671 18512 31677
rect 18493 31637 18505 31671
rect 18493 31631 18512 31637
rect 18506 31628 18512 31631
rect 18564 31628 18570 31680
rect 18616 31668 18644 31708
rect 18693 31705 18705 31739
rect 18739 31736 18751 31739
rect 18966 31736 18972 31748
rect 18739 31708 18972 31736
rect 18739 31705 18751 31708
rect 18693 31699 18751 31705
rect 18966 31696 18972 31708
rect 19024 31696 19030 31748
rect 20346 31736 20352 31748
rect 20404 31745 20410 31748
rect 20316 31708 20352 31736
rect 20346 31696 20352 31708
rect 20404 31699 20416 31745
rect 22281 31739 22339 31745
rect 22281 31705 22293 31739
rect 22327 31736 22339 31739
rect 22738 31736 22744 31748
rect 22327 31708 22744 31736
rect 22327 31705 22339 31708
rect 22281 31699 22339 31705
rect 20404 31696 20410 31699
rect 22738 31696 22744 31708
rect 22796 31696 22802 31748
rect 23290 31745 23296 31748
rect 23272 31739 23296 31745
rect 23272 31705 23284 31739
rect 23272 31699 23296 31705
rect 23290 31696 23296 31699
rect 23348 31696 23354 31748
rect 23477 31739 23535 31745
rect 23477 31705 23489 31739
rect 23523 31705 23535 31739
rect 25608 31736 25636 31776
rect 26418 31764 26424 31816
rect 26476 31804 26482 31816
rect 27505 31807 27563 31813
rect 27505 31804 27517 31807
rect 26476 31776 27517 31804
rect 26476 31764 26482 31776
rect 27505 31773 27517 31776
rect 27551 31773 27563 31807
rect 29638 31804 29644 31816
rect 29551 31776 29644 31804
rect 27505 31767 27563 31773
rect 29638 31764 29644 31776
rect 29696 31804 29702 31816
rect 30282 31804 30288 31816
rect 29696 31776 30288 31804
rect 29696 31764 29702 31776
rect 30282 31764 30288 31776
rect 30340 31764 30346 31816
rect 31409 31807 31467 31813
rect 31409 31773 31421 31807
rect 31455 31804 31467 31807
rect 31588 31804 31616 31844
rect 32122 31832 32128 31844
rect 32180 31832 32186 31884
rect 31455 31776 31616 31804
rect 31665 31807 31723 31813
rect 31455 31773 31467 31776
rect 31409 31767 31467 31773
rect 31665 31773 31677 31807
rect 31711 31804 31723 31807
rect 31754 31804 31760 31816
rect 31711 31776 31760 31804
rect 31711 31773 31723 31776
rect 31665 31767 31723 31773
rect 31754 31764 31760 31776
rect 31812 31804 31818 31816
rect 32766 31804 32772 31816
rect 31812 31776 32772 31804
rect 31812 31764 31818 31776
rect 32766 31764 32772 31776
rect 32824 31804 32830 31816
rect 34790 31804 34796 31816
rect 32824 31776 34796 31804
rect 32824 31764 32830 31776
rect 34790 31764 34796 31776
rect 34848 31764 34854 31816
rect 35060 31807 35118 31813
rect 35060 31773 35072 31807
rect 35106 31804 35118 31807
rect 35434 31804 35440 31816
rect 35106 31776 35440 31804
rect 35106 31773 35118 31776
rect 35060 31767 35118 31773
rect 35434 31764 35440 31776
rect 35492 31764 35498 31816
rect 36630 31764 36636 31816
rect 36688 31804 36694 31816
rect 36817 31807 36875 31813
rect 36817 31804 36829 31807
rect 36688 31776 36829 31804
rect 36688 31764 36694 31776
rect 36817 31773 36829 31776
rect 36863 31773 36875 31807
rect 36817 31767 36875 31773
rect 25958 31736 25964 31748
rect 25608 31708 25964 31736
rect 23477 31699 23535 31705
rect 19150 31668 19156 31680
rect 18616 31640 19156 31668
rect 19150 31628 19156 31640
rect 19208 31668 19214 31680
rect 19245 31671 19303 31677
rect 19245 31668 19257 31671
rect 19208 31640 19257 31668
rect 19208 31628 19214 31640
rect 19245 31637 19257 31640
rect 19291 31637 19303 31671
rect 23106 31668 23112 31680
rect 23067 31640 23112 31668
rect 19245 31631 19303 31637
rect 23106 31628 23112 31640
rect 23164 31628 23170 31680
rect 23492 31668 23520 31699
rect 25958 31696 25964 31708
rect 26016 31696 26022 31748
rect 26142 31696 26148 31748
rect 26200 31736 26206 31748
rect 30466 31736 30472 31748
rect 26200 31708 30472 31736
rect 26200 31696 26206 31708
rect 30466 31696 30472 31708
rect 30524 31696 30530 31748
rect 26160 31668 26188 31696
rect 23492 31640 26188 31668
rect 30285 31671 30343 31677
rect 30285 31637 30297 31671
rect 30331 31668 30343 31671
rect 30834 31668 30840 31680
rect 30331 31640 30840 31668
rect 30331 31637 30343 31640
rect 30285 31631 30343 31637
rect 30834 31628 30840 31640
rect 30892 31628 30898 31680
rect 36630 31668 36636 31680
rect 36591 31640 36636 31668
rect 36630 31628 36636 31640
rect 36688 31628 36694 31680
rect 1104 31578 44896 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 44896 31578
rect 1104 31504 44896 31526
rect 15562 31424 15568 31476
rect 15620 31464 15626 31476
rect 16025 31467 16083 31473
rect 16025 31464 16037 31467
rect 15620 31436 16037 31464
rect 15620 31424 15626 31436
rect 16025 31433 16037 31436
rect 16071 31433 16083 31467
rect 16025 31427 16083 31433
rect 16040 31396 16068 31427
rect 18598 31424 18604 31476
rect 18656 31464 18662 31476
rect 18656 31436 22094 31464
rect 18656 31424 18662 31436
rect 16040 31368 16988 31396
rect 14176 31331 14234 31337
rect 14176 31297 14188 31331
rect 14222 31328 14234 31331
rect 15470 31328 15476 31340
rect 14222 31300 15476 31328
rect 14222 31297 14234 31300
rect 14176 31291 14234 31297
rect 15470 31288 15476 31300
rect 15528 31288 15534 31340
rect 15746 31288 15752 31340
rect 15804 31328 15810 31340
rect 15841 31331 15899 31337
rect 15841 31328 15853 31331
rect 15804 31300 15853 31328
rect 15804 31288 15810 31300
rect 15841 31297 15853 31300
rect 15887 31297 15899 31331
rect 15841 31291 15899 31297
rect 13906 31260 13912 31272
rect 13867 31232 13912 31260
rect 13906 31220 13912 31232
rect 13964 31220 13970 31272
rect 15856 31260 15884 31291
rect 16114 31288 16120 31340
rect 16172 31328 16178 31340
rect 16666 31328 16672 31340
rect 16172 31300 16217 31328
rect 16627 31300 16672 31328
rect 16172 31288 16178 31300
rect 16666 31288 16672 31300
rect 16724 31288 16730 31340
rect 16960 31337 16988 31368
rect 19242 31356 19248 31408
rect 19300 31396 19306 31408
rect 22066 31396 22094 31436
rect 22278 31424 22284 31476
rect 22336 31464 22342 31476
rect 23382 31464 23388 31476
rect 22336 31436 23388 31464
rect 22336 31424 22342 31436
rect 23382 31424 23388 31436
rect 23440 31424 23446 31476
rect 25222 31464 25228 31476
rect 24136 31436 25228 31464
rect 24136 31396 24164 31436
rect 25222 31424 25228 31436
rect 25280 31424 25286 31476
rect 26970 31424 26976 31476
rect 27028 31464 27034 31476
rect 27223 31467 27281 31473
rect 27223 31464 27235 31467
rect 27028 31436 27235 31464
rect 27028 31424 27034 31436
rect 27223 31433 27235 31436
rect 27269 31433 27281 31467
rect 27223 31427 27281 31433
rect 31573 31467 31631 31473
rect 31573 31433 31585 31467
rect 31619 31464 31631 31467
rect 32122 31464 32128 31476
rect 31619 31436 31754 31464
rect 32083 31436 32128 31464
rect 31619 31433 31631 31436
rect 31573 31427 31631 31433
rect 19300 31368 19932 31396
rect 22066 31368 24164 31396
rect 19300 31356 19306 31368
rect 19904 31337 19932 31368
rect 24210 31356 24216 31408
rect 24268 31396 24274 31408
rect 24581 31399 24639 31405
rect 24581 31396 24593 31399
rect 24268 31368 24593 31396
rect 24268 31356 24274 31368
rect 24581 31365 24593 31368
rect 24627 31365 24639 31399
rect 24581 31359 24639 31365
rect 25774 31356 25780 31408
rect 25832 31396 25838 31408
rect 27433 31399 27491 31405
rect 27433 31396 27445 31399
rect 25832 31368 27445 31396
rect 25832 31356 25838 31368
rect 27433 31365 27445 31368
rect 27479 31396 27491 31399
rect 28166 31396 28172 31408
rect 27479 31368 28172 31396
rect 27479 31365 27491 31368
rect 27433 31359 27491 31365
rect 28166 31356 28172 31368
rect 28224 31396 28230 31408
rect 31205 31399 31263 31405
rect 28224 31368 30236 31396
rect 28224 31356 28230 31368
rect 20162 31337 20168 31340
rect 16945 31331 17003 31337
rect 16945 31297 16957 31331
rect 16991 31297 17003 31331
rect 16945 31291 17003 31297
rect 19889 31331 19947 31337
rect 19889 31297 19901 31331
rect 19935 31297 19947 31331
rect 19889 31291 19947 31297
rect 20156 31291 20168 31337
rect 20220 31328 20226 31340
rect 22278 31337 22284 31340
rect 20220 31300 20256 31328
rect 20162 31288 20168 31291
rect 20220 31288 20226 31300
rect 22272 31291 22284 31337
rect 22336 31328 22342 31340
rect 25593 31331 25651 31337
rect 22336 31300 22372 31328
rect 22278 31288 22284 31291
rect 22336 31288 22342 31300
rect 25593 31297 25605 31331
rect 25639 31328 25651 31331
rect 25866 31328 25872 31340
rect 25639 31300 25872 31328
rect 25639 31297 25651 31300
rect 25593 31291 25651 31297
rect 25866 31288 25872 31300
rect 25924 31288 25930 31340
rect 26326 31328 26332 31340
rect 26287 31300 26332 31328
rect 26326 31288 26332 31300
rect 26384 31288 26390 31340
rect 28261 31331 28319 31337
rect 28261 31297 28273 31331
rect 28307 31328 28319 31331
rect 28442 31328 28448 31340
rect 28307 31300 28448 31328
rect 28307 31297 28319 31300
rect 28261 31291 28319 31297
rect 28442 31288 28448 31300
rect 28500 31288 28506 31340
rect 30208 31337 30236 31368
rect 31205 31365 31217 31399
rect 31251 31365 31263 31399
rect 31205 31359 31263 31365
rect 30193 31331 30251 31337
rect 30193 31297 30205 31331
rect 30239 31328 30251 31331
rect 31220 31328 31248 31359
rect 31294 31356 31300 31408
rect 31352 31396 31358 31408
rect 31405 31399 31463 31405
rect 31405 31396 31417 31399
rect 31352 31368 31417 31396
rect 31352 31356 31358 31368
rect 31405 31365 31417 31368
rect 31451 31365 31463 31399
rect 31405 31359 31463 31365
rect 30239 31300 31248 31328
rect 31726 31328 31754 31436
rect 32122 31424 32128 31436
rect 32180 31424 32186 31476
rect 35161 31399 35219 31405
rect 35161 31365 35173 31399
rect 35207 31396 35219 31399
rect 35342 31396 35348 31408
rect 35207 31368 35348 31396
rect 35207 31365 35219 31368
rect 35161 31359 35219 31365
rect 35342 31356 35348 31368
rect 35400 31356 35406 31408
rect 32309 31331 32367 31337
rect 32309 31328 32321 31331
rect 31726 31300 32321 31328
rect 30239 31297 30251 31300
rect 30193 31291 30251 31297
rect 32309 31297 32321 31300
rect 32355 31297 32367 31331
rect 32309 31291 32367 31297
rect 16390 31260 16396 31272
rect 15856 31232 16396 31260
rect 16390 31220 16396 31232
rect 16448 31220 16454 31272
rect 18966 31260 18972 31272
rect 18927 31232 18972 31260
rect 18966 31220 18972 31232
rect 19024 31220 19030 31272
rect 19150 31220 19156 31272
rect 19208 31260 19214 31272
rect 19245 31263 19303 31269
rect 19245 31260 19257 31263
rect 19208 31232 19257 31260
rect 19208 31220 19214 31232
rect 19245 31229 19257 31232
rect 19291 31229 19303 31263
rect 19245 31223 19303 31229
rect 21174 31220 21180 31272
rect 21232 31260 21238 31272
rect 21818 31260 21824 31272
rect 21232 31232 21824 31260
rect 21232 31220 21238 31232
rect 21818 31220 21824 31232
rect 21876 31260 21882 31272
rect 22005 31263 22063 31269
rect 22005 31260 22017 31263
rect 21876 31232 22017 31260
rect 21876 31220 21882 31232
rect 22005 31229 22017 31232
rect 22051 31229 22063 31263
rect 25884 31260 25912 31288
rect 29638 31260 29644 31272
rect 25884 31232 29644 31260
rect 22005 31223 22063 31229
rect 29638 31220 29644 31232
rect 29696 31220 29702 31272
rect 29917 31263 29975 31269
rect 29917 31229 29929 31263
rect 29963 31260 29975 31263
rect 30374 31260 30380 31272
rect 29963 31232 30380 31260
rect 29963 31229 29975 31232
rect 29917 31223 29975 31229
rect 30374 31220 30380 31232
rect 30432 31260 30438 31272
rect 30742 31260 30748 31272
rect 30432 31232 30748 31260
rect 30432 31220 30438 31232
rect 30742 31220 30748 31232
rect 30800 31220 30806 31272
rect 15838 31192 15844 31204
rect 15799 31164 15844 31192
rect 15838 31152 15844 31164
rect 15896 31152 15902 31204
rect 24765 31195 24823 31201
rect 24765 31161 24777 31195
rect 24811 31192 24823 31195
rect 25682 31192 25688 31204
rect 24811 31164 25688 31192
rect 24811 31161 24823 31164
rect 24765 31155 24823 31161
rect 25682 31152 25688 31164
rect 25740 31152 25746 31204
rect 26418 31152 26424 31204
rect 26476 31192 26482 31204
rect 27065 31195 27123 31201
rect 27065 31192 27077 31195
rect 26476 31164 27077 31192
rect 26476 31152 26482 31164
rect 27065 31161 27077 31164
rect 27111 31161 27123 31195
rect 27065 31155 27123 31161
rect 34790 31152 34796 31204
rect 34848 31192 34854 31204
rect 34977 31195 35035 31201
rect 34977 31192 34989 31195
rect 34848 31164 34989 31192
rect 34848 31152 34854 31164
rect 34977 31161 34989 31164
rect 35023 31161 35035 31195
rect 34977 31155 35035 31161
rect 15289 31127 15347 31133
rect 15289 31093 15301 31127
rect 15335 31124 15347 31127
rect 16482 31124 16488 31136
rect 15335 31096 16488 31124
rect 15335 31093 15347 31096
rect 15289 31087 15347 31093
rect 16482 31084 16488 31096
rect 16540 31084 16546 31136
rect 21266 31124 21272 31136
rect 21227 31096 21272 31124
rect 21266 31084 21272 31096
rect 21324 31084 21330 31136
rect 25314 31124 25320 31136
rect 25275 31096 25320 31124
rect 25314 31084 25320 31096
rect 25372 31084 25378 31136
rect 25958 31084 25964 31136
rect 26016 31124 26022 31136
rect 26145 31127 26203 31133
rect 26145 31124 26157 31127
rect 26016 31096 26157 31124
rect 26016 31084 26022 31096
rect 26145 31093 26157 31096
rect 26191 31093 26203 31127
rect 27246 31124 27252 31136
rect 27207 31096 27252 31124
rect 26145 31087 26203 31093
rect 27246 31084 27252 31096
rect 27304 31084 27310 31136
rect 28074 31124 28080 31136
rect 28035 31096 28080 31124
rect 28074 31084 28080 31096
rect 28132 31084 28138 31136
rect 31110 31084 31116 31136
rect 31168 31124 31174 31136
rect 31389 31127 31447 31133
rect 31389 31124 31401 31127
rect 31168 31096 31401 31124
rect 31168 31084 31174 31096
rect 31389 31093 31401 31096
rect 31435 31093 31447 31127
rect 31389 31087 31447 31093
rect 1104 31034 44896 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 44896 31034
rect 1104 30960 44896 30982
rect 15470 30920 15476 30932
rect 15431 30892 15476 30920
rect 15470 30880 15476 30892
rect 15528 30880 15534 30932
rect 16666 30920 16672 30932
rect 15672 30892 16672 30920
rect 1762 30716 1768 30728
rect 1723 30688 1768 30716
rect 1762 30676 1768 30688
rect 1820 30676 1826 30728
rect 15672 30725 15700 30892
rect 16666 30880 16672 30892
rect 16724 30880 16730 30932
rect 17681 30923 17739 30929
rect 17681 30889 17693 30923
rect 17727 30920 17739 30923
rect 18138 30920 18144 30932
rect 17727 30892 18144 30920
rect 17727 30889 17739 30892
rect 17681 30883 17739 30889
rect 15838 30852 15844 30864
rect 15799 30824 15844 30852
rect 15838 30812 15844 30824
rect 15896 30812 15902 30864
rect 16390 30812 16396 30864
rect 16448 30852 16454 30864
rect 17696 30852 17724 30883
rect 18138 30880 18144 30892
rect 18196 30880 18202 30932
rect 20162 30880 20168 30932
rect 20220 30920 20226 30932
rect 20257 30923 20315 30929
rect 20257 30920 20269 30923
rect 20220 30892 20269 30920
rect 20220 30880 20226 30892
rect 20257 30889 20269 30892
rect 20303 30889 20315 30923
rect 20257 30883 20315 30889
rect 22278 30880 22284 30932
rect 22336 30920 22342 30932
rect 22373 30923 22431 30929
rect 22373 30920 22385 30923
rect 22336 30892 22385 30920
rect 22336 30880 22342 30892
rect 22373 30889 22385 30892
rect 22419 30889 22431 30923
rect 23750 30920 23756 30932
rect 23711 30892 23756 30920
rect 22373 30883 22431 30889
rect 23750 30880 23756 30892
rect 23808 30880 23814 30932
rect 25222 30880 25228 30932
rect 25280 30920 25286 30932
rect 25501 30923 25559 30929
rect 25501 30920 25513 30923
rect 25280 30892 25513 30920
rect 25280 30880 25286 30892
rect 25501 30889 25513 30892
rect 25547 30889 25559 30923
rect 28258 30920 28264 30932
rect 28219 30892 28264 30920
rect 25501 30883 25559 30889
rect 28258 30880 28264 30892
rect 28316 30880 28322 30932
rect 28442 30920 28448 30932
rect 28403 30892 28448 30920
rect 28442 30880 28448 30892
rect 28500 30880 28506 30932
rect 31110 30920 31116 30932
rect 31071 30892 31116 30920
rect 31110 30880 31116 30892
rect 31168 30880 31174 30932
rect 37369 30923 37427 30929
rect 37369 30889 37381 30923
rect 37415 30920 37427 30923
rect 37550 30920 37556 30932
rect 37415 30892 37556 30920
rect 37415 30889 37427 30892
rect 37369 30883 37427 30889
rect 37550 30880 37556 30892
rect 37608 30880 37614 30932
rect 18598 30852 18604 30864
rect 16448 30824 17724 30852
rect 17788 30824 18604 30852
rect 16448 30812 16454 30824
rect 15749 30787 15807 30793
rect 15749 30753 15761 30787
rect 15795 30784 15807 30787
rect 16022 30784 16028 30796
rect 15795 30756 16028 30784
rect 15795 30753 15807 30756
rect 15749 30747 15807 30753
rect 16022 30744 16028 30756
rect 16080 30744 16086 30796
rect 16850 30784 16856 30796
rect 16132 30756 16856 30784
rect 15657 30719 15715 30725
rect 15657 30685 15669 30719
rect 15703 30685 15715 30719
rect 15657 30679 15715 30685
rect 15930 30676 15936 30728
rect 15988 30716 15994 30728
rect 16132 30725 16160 30756
rect 16850 30744 16856 30756
rect 16908 30784 16914 30796
rect 17788 30784 17816 30824
rect 18598 30812 18604 30824
rect 18656 30812 18662 30864
rect 21266 30852 21272 30864
rect 20548 30824 21272 30852
rect 17954 30784 17960 30796
rect 16908 30756 17816 30784
rect 17915 30756 17960 30784
rect 16908 30744 16914 30756
rect 17954 30744 17960 30756
rect 18012 30744 18018 30796
rect 18138 30784 18144 30796
rect 18099 30756 18144 30784
rect 18138 30744 18144 30756
rect 18196 30744 18202 30796
rect 16117 30719 16175 30725
rect 15988 30688 16033 30716
rect 15988 30676 15994 30688
rect 16117 30685 16129 30719
rect 16163 30685 16175 30719
rect 16117 30679 16175 30685
rect 16482 30676 16488 30728
rect 16540 30716 16546 30728
rect 16761 30719 16819 30725
rect 16761 30716 16773 30719
rect 16540 30688 16773 30716
rect 16540 30676 16546 30688
rect 16761 30685 16773 30688
rect 16807 30685 16819 30719
rect 16761 30679 16819 30685
rect 17310 30676 17316 30728
rect 17368 30716 17374 30728
rect 17865 30719 17923 30725
rect 17865 30716 17877 30719
rect 17368 30688 17877 30716
rect 17368 30676 17374 30688
rect 17865 30685 17877 30688
rect 17911 30685 17923 30719
rect 17865 30679 17923 30685
rect 18046 30676 18052 30728
rect 18104 30716 18110 30728
rect 18104 30688 18149 30716
rect 18104 30676 18110 30688
rect 18506 30676 18512 30728
rect 18564 30716 18570 30728
rect 20548 30725 20576 30824
rect 21266 30812 21272 30824
rect 21324 30812 21330 30864
rect 22738 30784 22744 30796
rect 20640 30756 22744 30784
rect 20640 30725 20668 30756
rect 22738 30744 22744 30756
rect 22796 30744 22802 30796
rect 23768 30784 23796 30880
rect 23842 30812 23848 30864
rect 23900 30852 23906 30864
rect 26605 30855 26663 30861
rect 26605 30852 26617 30855
rect 23900 30824 26617 30852
rect 23900 30812 23906 30824
rect 24581 30787 24639 30793
rect 24581 30784 24593 30787
rect 23768 30756 24593 30784
rect 24581 30753 24593 30756
rect 24627 30753 24639 30787
rect 24762 30784 24768 30796
rect 24723 30756 24768 30784
rect 24581 30747 24639 30753
rect 24762 30744 24768 30756
rect 24820 30744 24826 30796
rect 19245 30719 19303 30725
rect 19245 30716 19257 30719
rect 18564 30688 19257 30716
rect 18564 30676 18570 30688
rect 19245 30685 19257 30688
rect 19291 30685 19303 30719
rect 19245 30679 19303 30685
rect 20533 30719 20591 30725
rect 20533 30685 20545 30719
rect 20579 30685 20591 30719
rect 20533 30679 20591 30685
rect 20625 30719 20683 30725
rect 20625 30685 20637 30719
rect 20671 30685 20683 30719
rect 20625 30679 20683 30685
rect 20714 30676 20720 30728
rect 20772 30716 20778 30728
rect 20772 30688 20817 30716
rect 20772 30676 20778 30688
rect 20898 30676 20904 30728
rect 20956 30716 20962 30728
rect 22557 30719 22615 30725
rect 20956 30688 21001 30716
rect 20956 30676 20962 30688
rect 22557 30685 22569 30719
rect 22603 30716 22615 30719
rect 23106 30716 23112 30728
rect 22603 30688 23112 30716
rect 22603 30685 22615 30688
rect 22557 30679 22615 30685
rect 23106 30676 23112 30688
rect 23164 30676 23170 30728
rect 24489 30719 24547 30725
rect 24489 30685 24501 30719
rect 24535 30685 24547 30719
rect 24489 30679 24547 30685
rect 24673 30719 24731 30725
rect 24673 30685 24685 30719
rect 24719 30716 24731 30719
rect 24872 30716 24900 30824
rect 26605 30821 26617 30824
rect 26651 30852 26663 30855
rect 27154 30852 27160 30864
rect 26651 30824 27160 30852
rect 26651 30821 26663 30824
rect 26605 30815 26663 30821
rect 27154 30812 27160 30824
rect 27212 30812 27218 30864
rect 30466 30812 30472 30864
rect 30524 30852 30530 30864
rect 30524 30824 31795 30852
rect 30524 30812 30530 30824
rect 27525 30787 27583 30793
rect 27525 30753 27537 30787
rect 27571 30753 27583 30787
rect 27525 30747 27583 30753
rect 25774 30716 25780 30728
rect 24719 30688 24900 30716
rect 25735 30688 25780 30716
rect 24719 30685 24731 30688
rect 24673 30679 24731 30685
rect 8018 30608 8024 30660
rect 8076 30648 8082 30660
rect 23661 30651 23719 30657
rect 23661 30648 23673 30651
rect 8076 30620 23673 30648
rect 8076 30608 8082 30620
rect 23661 30617 23673 30620
rect 23707 30648 23719 30651
rect 24302 30648 24308 30660
rect 23707 30620 24308 30648
rect 23707 30617 23719 30620
rect 23661 30611 23719 30617
rect 24302 30608 24308 30620
rect 24360 30608 24366 30660
rect 24504 30648 24532 30679
rect 25774 30676 25780 30688
rect 25832 30676 25838 30728
rect 27430 30716 27436 30728
rect 27391 30688 27436 30716
rect 27430 30676 27436 30688
rect 27488 30676 27494 30728
rect 25590 30648 25596 30660
rect 24504 30620 25596 30648
rect 25590 30608 25596 30620
rect 25648 30608 25654 30660
rect 26418 30648 26424 30660
rect 26379 30620 26424 30648
rect 26418 30608 26424 30620
rect 26476 30608 26482 30660
rect 19334 30580 19340 30592
rect 19295 30552 19340 30580
rect 19334 30540 19340 30552
rect 19392 30540 19398 30592
rect 24949 30583 25007 30589
rect 24949 30549 24961 30583
rect 24995 30580 25007 30583
rect 25406 30580 25412 30592
rect 24995 30552 25412 30580
rect 24995 30549 25007 30552
rect 24949 30543 25007 30549
rect 25406 30540 25412 30552
rect 25464 30540 25470 30592
rect 27062 30580 27068 30592
rect 27023 30552 27068 30580
rect 27062 30540 27068 30552
rect 27120 30540 27126 30592
rect 27540 30580 27568 30747
rect 30650 30716 30656 30728
rect 30611 30688 30656 30716
rect 30650 30676 30656 30688
rect 30708 30676 30714 30728
rect 30834 30676 30840 30728
rect 30892 30716 30898 30728
rect 30929 30719 30987 30725
rect 30929 30716 30941 30719
rect 30892 30688 30941 30716
rect 30892 30676 30898 30688
rect 30929 30685 30941 30688
rect 30975 30685 30987 30719
rect 30929 30679 30987 30685
rect 31018 30676 31024 30728
rect 31076 30716 31082 30728
rect 31767 30725 31795 30824
rect 31846 30812 31852 30864
rect 31904 30852 31910 30864
rect 31904 30824 31984 30852
rect 31904 30812 31910 30824
rect 31956 30725 31984 30824
rect 31573 30719 31631 30725
rect 31573 30716 31585 30719
rect 31076 30688 31585 30716
rect 31076 30676 31082 30688
rect 31573 30685 31585 30688
rect 31619 30685 31631 30719
rect 31573 30679 31631 30685
rect 31752 30719 31810 30725
rect 31752 30685 31764 30719
rect 31798 30685 31810 30719
rect 31852 30716 31910 30722
rect 31852 30706 31864 30716
rect 31898 30706 31910 30716
rect 31752 30679 31810 30685
rect 28077 30651 28135 30657
rect 28077 30617 28089 30651
rect 28123 30648 28135 30651
rect 28166 30648 28172 30660
rect 28123 30620 28172 30648
rect 28123 30617 28135 30620
rect 28077 30611 28135 30617
rect 28166 30608 28172 30620
rect 28224 30608 28230 30660
rect 30006 30608 30012 30660
rect 30064 30648 30070 30660
rect 30745 30651 30803 30657
rect 30745 30648 30757 30651
rect 30064 30620 30757 30648
rect 30064 30608 30070 30620
rect 30745 30617 30757 30620
rect 30791 30648 30803 30651
rect 31662 30648 31668 30660
rect 30791 30620 31668 30648
rect 30791 30617 30803 30620
rect 30745 30611 30803 30617
rect 31662 30608 31668 30620
rect 31720 30608 31726 30660
rect 31846 30654 31852 30706
rect 31904 30654 31910 30706
rect 31941 30719 31999 30725
rect 31941 30685 31953 30719
rect 31987 30685 31999 30719
rect 32766 30716 32772 30728
rect 32727 30688 32772 30716
rect 31941 30679 31999 30685
rect 32766 30676 32772 30688
rect 32824 30676 32830 30728
rect 35986 30716 35992 30728
rect 35947 30688 35992 30716
rect 35986 30676 35992 30688
rect 36044 30676 36050 30728
rect 36256 30719 36314 30725
rect 36256 30685 36268 30719
rect 36302 30716 36314 30719
rect 36630 30716 36636 30728
rect 36302 30688 36636 30716
rect 36302 30685 36314 30688
rect 36256 30679 36314 30685
rect 36630 30676 36636 30688
rect 36688 30676 36694 30728
rect 32217 30651 32275 30657
rect 32217 30617 32229 30651
rect 32263 30648 32275 30651
rect 33014 30651 33072 30657
rect 33014 30648 33026 30651
rect 32263 30620 33026 30648
rect 32263 30617 32275 30620
rect 32217 30611 32275 30617
rect 33014 30617 33026 30620
rect 33060 30617 33072 30651
rect 43714 30648 43720 30660
rect 43675 30620 43720 30648
rect 33014 30611 33072 30617
rect 43714 30608 43720 30620
rect 43772 30608 43778 30660
rect 44082 30648 44088 30660
rect 44043 30620 44088 30648
rect 44082 30608 44088 30620
rect 44140 30608 44146 30660
rect 28287 30583 28345 30589
rect 28287 30580 28299 30583
rect 27540 30552 28299 30580
rect 28287 30549 28299 30552
rect 28333 30580 28345 30583
rect 28810 30580 28816 30592
rect 28333 30552 28816 30580
rect 28333 30549 28345 30552
rect 28287 30543 28345 30549
rect 28810 30540 28816 30552
rect 28868 30540 28874 30592
rect 30834 30540 30840 30592
rect 30892 30580 30898 30592
rect 33686 30580 33692 30592
rect 30892 30552 33692 30580
rect 30892 30540 30898 30552
rect 33686 30540 33692 30552
rect 33744 30540 33750 30592
rect 33870 30540 33876 30592
rect 33928 30580 33934 30592
rect 34149 30583 34207 30589
rect 34149 30580 34161 30583
rect 33928 30552 34161 30580
rect 33928 30540 33934 30552
rect 34149 30549 34161 30552
rect 34195 30549 34207 30583
rect 34149 30543 34207 30549
rect 1104 30490 44896 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 44896 30490
rect 1104 30416 44896 30438
rect 26326 30376 26332 30388
rect 26287 30348 26332 30376
rect 26326 30336 26332 30348
rect 26384 30336 26390 30388
rect 30466 30376 30472 30388
rect 30427 30348 30472 30376
rect 30466 30336 30472 30348
rect 30524 30336 30530 30388
rect 16666 30268 16672 30320
rect 16724 30308 16730 30320
rect 17586 30308 17592 30320
rect 16724 30280 17592 30308
rect 16724 30268 16730 30280
rect 17586 30268 17592 30280
rect 17644 30308 17650 30320
rect 18141 30311 18199 30317
rect 18141 30308 18153 30311
rect 17644 30280 18153 30308
rect 17644 30268 17650 30280
rect 18141 30277 18153 30280
rect 18187 30277 18199 30311
rect 19334 30308 19340 30320
rect 18141 30271 18199 30277
rect 18432 30280 19340 30308
rect 1762 30240 1768 30252
rect 1723 30212 1768 30240
rect 1762 30200 1768 30212
rect 1820 30200 1826 30252
rect 16758 30200 16764 30252
rect 16816 30240 16822 30252
rect 17037 30243 17095 30249
rect 17037 30240 17049 30243
rect 16816 30212 17049 30240
rect 16816 30200 16822 30212
rect 17037 30209 17049 30212
rect 17083 30209 17095 30243
rect 17037 30203 17095 30209
rect 17129 30243 17187 30249
rect 17129 30209 17141 30243
rect 17175 30209 17187 30243
rect 17129 30203 17187 30209
rect 17313 30243 17371 30249
rect 17313 30209 17325 30243
rect 17359 30240 17371 30243
rect 18044 30243 18102 30249
rect 18044 30240 18056 30243
rect 17359 30212 17908 30240
rect 17359 30209 17371 30212
rect 17313 30203 17371 30209
rect 1949 30175 2007 30181
rect 1949 30141 1961 30175
rect 1995 30172 2007 30175
rect 2222 30172 2228 30184
rect 1995 30144 2228 30172
rect 1995 30141 2007 30144
rect 1949 30135 2007 30141
rect 2222 30132 2228 30144
rect 2280 30132 2286 30184
rect 2774 30172 2780 30184
rect 2735 30144 2780 30172
rect 2774 30132 2780 30144
rect 2832 30132 2838 30184
rect 15838 30132 15844 30184
rect 15896 30172 15902 30184
rect 17144 30172 17172 30203
rect 15896 30144 17172 30172
rect 15896 30132 15902 30144
rect 17310 30104 17316 30116
rect 17271 30076 17316 30104
rect 17310 30064 17316 30076
rect 17368 30064 17374 30116
rect 17880 30113 17908 30212
rect 17972 30212 18056 30240
rect 17865 30107 17923 30113
rect 17865 30073 17877 30107
rect 17911 30073 17923 30107
rect 17865 30067 17923 30073
rect 17678 29996 17684 30048
rect 17736 30036 17742 30048
rect 17972 30036 18000 30212
rect 18044 30209 18056 30212
rect 18090 30209 18102 30243
rect 18230 30240 18236 30252
rect 18191 30212 18236 30240
rect 18044 30203 18102 30209
rect 18230 30200 18236 30212
rect 18288 30200 18294 30252
rect 18432 30249 18460 30280
rect 19334 30268 19340 30280
rect 19392 30268 19398 30320
rect 22094 30268 22100 30320
rect 22152 30308 22158 30320
rect 22465 30311 22523 30317
rect 22465 30308 22477 30311
rect 22152 30280 22477 30308
rect 22152 30268 22158 30280
rect 22465 30277 22477 30280
rect 22511 30277 22523 30311
rect 22465 30271 22523 30277
rect 24136 30280 25452 30308
rect 18416 30243 18474 30249
rect 18416 30209 18428 30243
rect 18462 30209 18474 30243
rect 18416 30203 18474 30209
rect 18509 30243 18567 30249
rect 18509 30209 18521 30243
rect 18555 30240 18567 30243
rect 19242 30240 19248 30252
rect 18555 30212 19248 30240
rect 18555 30209 18567 30212
rect 18509 30203 18567 30209
rect 19242 30200 19248 30212
rect 19300 30200 19306 30252
rect 20438 30200 20444 30252
rect 20496 30240 20502 30252
rect 22281 30243 22339 30249
rect 22281 30240 22293 30243
rect 20496 30212 22293 30240
rect 20496 30200 20502 30212
rect 22281 30209 22293 30212
rect 22327 30209 22339 30243
rect 22281 30203 22339 30209
rect 19058 30132 19064 30184
rect 19116 30172 19122 30184
rect 24136 30172 24164 30280
rect 24302 30240 24308 30252
rect 24263 30212 24308 30240
rect 24302 30200 24308 30212
rect 24360 30200 24366 30252
rect 24489 30243 24547 30249
rect 24489 30209 24501 30243
rect 24535 30240 24547 30243
rect 24762 30240 24768 30252
rect 24535 30212 24768 30240
rect 24535 30209 24547 30212
rect 24489 30203 24547 30209
rect 24762 30200 24768 30212
rect 24820 30200 24826 30252
rect 25133 30243 25191 30249
rect 25133 30209 25145 30243
rect 25179 30240 25191 30243
rect 25222 30240 25228 30252
rect 25179 30212 25228 30240
rect 25179 30209 25191 30212
rect 25133 30203 25191 30209
rect 19116 30144 24164 30172
rect 24213 30175 24271 30181
rect 19116 30132 19122 30144
rect 24213 30141 24225 30175
rect 24259 30141 24271 30175
rect 24213 30135 24271 30141
rect 24397 30175 24455 30181
rect 24397 30141 24409 30175
rect 24443 30172 24455 30175
rect 25148 30172 25176 30203
rect 25222 30200 25228 30212
rect 25280 30200 25286 30252
rect 25424 30240 25452 30280
rect 25774 30268 25780 30320
rect 25832 30308 25838 30320
rect 25961 30311 26019 30317
rect 25961 30308 25973 30311
rect 25832 30280 25973 30308
rect 25832 30268 25838 30280
rect 25961 30277 25973 30280
rect 26007 30277 26019 30311
rect 25961 30271 26019 30277
rect 26177 30311 26235 30317
rect 26177 30277 26189 30311
rect 26223 30308 26235 30311
rect 27062 30308 27068 30320
rect 26223 30280 27068 30308
rect 26223 30277 26235 30280
rect 26177 30271 26235 30277
rect 27062 30268 27068 30280
rect 27120 30268 27126 30320
rect 28074 30317 28080 30320
rect 28068 30308 28080 30317
rect 28035 30280 28080 30308
rect 28068 30271 28080 30280
rect 28074 30268 28080 30271
rect 28132 30268 28138 30320
rect 31573 30311 31631 30317
rect 31573 30277 31585 30311
rect 31619 30308 31631 30311
rect 33014 30311 33072 30317
rect 33014 30308 33026 30311
rect 31619 30280 33026 30308
rect 31619 30277 31631 30280
rect 31573 30271 31631 30277
rect 33014 30277 33026 30280
rect 33060 30277 33072 30311
rect 33014 30271 33072 30277
rect 34790 30268 34796 30320
rect 34848 30308 34854 30320
rect 36173 30311 36231 30317
rect 36173 30308 36185 30311
rect 34848 30280 36185 30308
rect 34848 30268 34854 30280
rect 36173 30277 36185 30280
rect 36219 30277 36231 30311
rect 36173 30271 36231 30277
rect 26510 30240 26516 30252
rect 25424 30212 26516 30240
rect 24443 30144 25176 30172
rect 24443 30141 24455 30144
rect 24397 30135 24455 30141
rect 24228 30104 24256 30135
rect 24854 30104 24860 30116
rect 24228 30076 24860 30104
rect 24854 30064 24860 30076
rect 24912 30064 24918 30116
rect 25317 30107 25375 30113
rect 25317 30073 25329 30107
rect 25363 30104 25375 30107
rect 25424 30104 25452 30212
rect 26510 30200 26516 30212
rect 26568 30200 26574 30252
rect 27157 30243 27215 30249
rect 27157 30209 27169 30243
rect 27203 30240 27215 30243
rect 28994 30240 29000 30252
rect 27203 30212 29000 30240
rect 27203 30209 27215 30212
rect 27157 30203 27215 30209
rect 28994 30200 29000 30212
rect 29052 30200 29058 30252
rect 30006 30240 30012 30252
rect 29967 30212 30012 30240
rect 30006 30200 30012 30212
rect 30064 30200 30070 30252
rect 30469 30243 30527 30249
rect 30469 30209 30481 30243
rect 30515 30240 30527 30243
rect 30650 30240 30656 30252
rect 30515 30212 30656 30240
rect 30515 30209 30527 30212
rect 30469 30203 30527 30209
rect 30650 30200 30656 30212
rect 30708 30200 30714 30252
rect 30926 30240 30932 30252
rect 30887 30212 30932 30240
rect 30926 30200 30932 30212
rect 30984 30200 30990 30252
rect 31113 30243 31171 30249
rect 31113 30209 31125 30243
rect 31159 30209 31171 30243
rect 31113 30203 31171 30209
rect 25682 30132 25688 30184
rect 25740 30172 25746 30184
rect 27801 30175 27859 30181
rect 27801 30172 27813 30175
rect 25740 30144 27813 30172
rect 25740 30132 25746 30144
rect 27801 30141 27813 30144
rect 27847 30141 27859 30175
rect 31128 30172 31156 30203
rect 31202 30200 31208 30252
rect 31260 30240 31266 30252
rect 31343 30243 31401 30249
rect 31260 30212 31305 30240
rect 31260 30200 31266 30212
rect 31343 30209 31355 30243
rect 31389 30240 31401 30243
rect 31478 30240 31484 30252
rect 31389 30212 31484 30240
rect 31389 30209 31401 30212
rect 31343 30203 31401 30209
rect 31478 30200 31484 30212
rect 31536 30200 31542 30252
rect 31846 30200 31852 30252
rect 31904 30240 31910 30252
rect 32125 30243 32183 30249
rect 32125 30240 32137 30243
rect 31904 30212 32137 30240
rect 31904 30200 31910 30212
rect 32125 30209 32137 30212
rect 32171 30209 32183 30243
rect 32306 30240 32312 30252
rect 32267 30212 32312 30240
rect 32125 30203 32183 30209
rect 32306 30200 32312 30212
rect 32364 30200 32370 30252
rect 34514 30200 34520 30252
rect 34572 30240 34578 30252
rect 34885 30243 34943 30249
rect 34885 30240 34897 30243
rect 34572 30212 34897 30240
rect 34572 30200 34578 30212
rect 34885 30209 34897 30212
rect 34931 30209 34943 30243
rect 37458 30240 37464 30252
rect 37419 30212 37464 30240
rect 34885 30203 34943 30209
rect 37458 30200 37464 30212
rect 37516 30200 37522 30252
rect 43346 30240 43352 30252
rect 43307 30212 43352 30240
rect 43346 30200 43352 30212
rect 43404 30200 43410 30252
rect 32766 30172 32772 30184
rect 31128 30144 31754 30172
rect 32727 30144 32772 30172
rect 27801 30135 27859 30141
rect 25363 30076 25452 30104
rect 25363 30073 25375 30076
rect 25317 30067 25375 30073
rect 25590 30064 25596 30116
rect 25648 30104 25654 30116
rect 27065 30107 27123 30113
rect 27065 30104 27077 30107
rect 25648 30076 27077 30104
rect 25648 30064 25654 30076
rect 27065 30073 27077 30076
rect 27111 30073 27123 30107
rect 31726 30104 31754 30144
rect 32766 30132 32772 30144
rect 32824 30132 32830 30184
rect 33870 30132 33876 30184
rect 33928 30172 33934 30184
rect 34609 30175 34667 30181
rect 34609 30172 34621 30175
rect 33928 30144 34621 30172
rect 33928 30132 33934 30144
rect 34609 30141 34621 30144
rect 34655 30141 34667 30175
rect 34609 30135 34667 30141
rect 32217 30107 32275 30113
rect 32217 30104 32229 30107
rect 31726 30076 32229 30104
rect 27065 30067 27123 30073
rect 32217 30073 32229 30076
rect 32263 30073 32275 30107
rect 32217 30067 32275 30073
rect 35986 30064 35992 30116
rect 36044 30104 36050 30116
rect 36357 30107 36415 30113
rect 36357 30104 36369 30107
rect 36044 30076 36369 30104
rect 36044 30064 36050 30076
rect 36357 30073 36369 30076
rect 36403 30104 36415 30107
rect 37182 30104 37188 30116
rect 36403 30076 37188 30104
rect 36403 30073 36415 30076
rect 36357 30067 36415 30073
rect 37182 30064 37188 30076
rect 37240 30064 37246 30116
rect 24670 30036 24676 30048
rect 17736 30008 18000 30036
rect 24631 30008 24676 30036
rect 17736 29996 17742 30008
rect 24670 29996 24676 30008
rect 24728 29996 24734 30048
rect 25406 29996 25412 30048
rect 25464 30036 25470 30048
rect 26050 30036 26056 30048
rect 25464 30008 26056 30036
rect 25464 29996 25470 30008
rect 26050 29996 26056 30008
rect 26108 30036 26114 30048
rect 26145 30039 26203 30045
rect 26145 30036 26157 30039
rect 26108 30008 26157 30036
rect 26108 29996 26114 30008
rect 26145 30005 26157 30008
rect 26191 30005 26203 30039
rect 26145 29999 26203 30005
rect 28902 29996 28908 30048
rect 28960 30036 28966 30048
rect 29181 30039 29239 30045
rect 29181 30036 29193 30039
rect 28960 30008 29193 30036
rect 28960 29996 28966 30008
rect 29181 30005 29193 30008
rect 29227 30005 29239 30039
rect 29181 29999 29239 30005
rect 29546 29996 29552 30048
rect 29604 30036 29610 30048
rect 30147 30039 30205 30045
rect 30147 30036 30159 30039
rect 29604 30008 30159 30036
rect 29604 29996 29610 30008
rect 30147 30005 30159 30008
rect 30193 30005 30205 30039
rect 30147 29999 30205 30005
rect 30285 30039 30343 30045
rect 30285 30005 30297 30039
rect 30331 30036 30343 30039
rect 30466 30036 30472 30048
rect 30331 30008 30472 30036
rect 30331 30005 30343 30008
rect 30285 29999 30343 30005
rect 30466 29996 30472 30008
rect 30524 29996 30530 30048
rect 33962 29996 33968 30048
rect 34020 30036 34026 30048
rect 34149 30039 34207 30045
rect 34149 30036 34161 30039
rect 34020 30008 34161 30036
rect 34020 29996 34026 30008
rect 34149 30005 34161 30008
rect 34195 30005 34207 30039
rect 34149 29999 34207 30005
rect 36814 29996 36820 30048
rect 36872 30036 36878 30048
rect 37277 30039 37335 30045
rect 37277 30036 37289 30039
rect 36872 30008 37289 30036
rect 36872 29996 36878 30008
rect 37277 30005 37289 30008
rect 37323 30005 37335 30039
rect 37277 29999 37335 30005
rect 43441 30039 43499 30045
rect 43441 30005 43453 30039
rect 43487 30036 43499 30039
rect 43990 30036 43996 30048
rect 43487 30008 43996 30036
rect 43487 30005 43499 30008
rect 43441 29999 43499 30005
rect 43990 29996 43996 30008
rect 44048 29996 44054 30048
rect 44174 30036 44180 30048
rect 44135 30008 44180 30036
rect 44174 29996 44180 30008
rect 44232 29996 44238 30048
rect 1104 29946 44896 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 44896 29946
rect 1104 29872 44896 29894
rect 2222 29832 2228 29844
rect 2183 29804 2228 29832
rect 2222 29792 2228 29804
rect 2280 29792 2286 29844
rect 15838 29832 15844 29844
rect 15799 29804 15844 29832
rect 15838 29792 15844 29804
rect 15896 29792 15902 29844
rect 16758 29832 16764 29844
rect 16719 29804 16764 29832
rect 16758 29792 16764 29804
rect 16816 29792 16822 29844
rect 18046 29792 18052 29844
rect 18104 29832 18110 29844
rect 18141 29835 18199 29841
rect 18141 29832 18153 29835
rect 18104 29804 18153 29832
rect 18104 29792 18110 29804
rect 18141 29801 18153 29804
rect 18187 29801 18199 29835
rect 19242 29832 19248 29844
rect 19203 29804 19248 29832
rect 18141 29795 18199 29801
rect 19242 29792 19248 29804
rect 19300 29792 19306 29844
rect 19978 29792 19984 29844
rect 20036 29832 20042 29844
rect 20625 29835 20683 29841
rect 20625 29832 20637 29835
rect 20036 29804 20637 29832
rect 20036 29792 20042 29804
rect 20625 29801 20637 29804
rect 20671 29832 20683 29835
rect 21450 29832 21456 29844
rect 20671 29804 21456 29832
rect 20671 29801 20683 29804
rect 20625 29795 20683 29801
rect 21450 29792 21456 29804
rect 21508 29792 21514 29844
rect 24670 29792 24676 29844
rect 24728 29832 24734 29844
rect 28258 29832 28264 29844
rect 24728 29804 28120 29832
rect 28219 29804 28264 29832
rect 24728 29792 24734 29804
rect 28092 29764 28120 29804
rect 28258 29792 28264 29804
rect 28316 29792 28322 29844
rect 28810 29832 28816 29844
rect 28771 29804 28816 29832
rect 28810 29792 28816 29804
rect 28868 29792 28874 29844
rect 30653 29835 30711 29841
rect 30653 29801 30665 29835
rect 30699 29832 30711 29835
rect 31294 29832 31300 29844
rect 30699 29804 31300 29832
rect 30699 29801 30711 29804
rect 30653 29795 30711 29801
rect 31294 29792 31300 29804
rect 31352 29792 31358 29844
rect 31386 29792 31392 29844
rect 31444 29832 31450 29844
rect 33594 29832 33600 29844
rect 31444 29804 33600 29832
rect 31444 29792 31450 29804
rect 33594 29792 33600 29804
rect 33652 29832 33658 29844
rect 43346 29832 43352 29844
rect 33652 29804 34100 29832
rect 33652 29792 33658 29804
rect 28534 29764 28540 29776
rect 28092 29736 28540 29764
rect 28534 29724 28540 29736
rect 28592 29724 28598 29776
rect 34072 29773 34100 29804
rect 34900 29804 43352 29832
rect 34057 29767 34115 29773
rect 34057 29733 34069 29767
rect 34103 29733 34115 29767
rect 34057 29727 34115 29733
rect 15562 29656 15568 29708
rect 15620 29696 15626 29708
rect 15620 29668 15976 29696
rect 15620 29656 15626 29668
rect 2317 29631 2375 29637
rect 2317 29597 2329 29631
rect 2363 29628 2375 29631
rect 2406 29628 2412 29640
rect 2363 29600 2412 29628
rect 2363 29597 2375 29600
rect 2317 29591 2375 29597
rect 2406 29588 2412 29600
rect 2464 29588 2470 29640
rect 14458 29628 14464 29640
rect 14419 29600 14464 29628
rect 14458 29588 14464 29600
rect 14516 29588 14522 29640
rect 15948 29637 15976 29668
rect 16482 29656 16488 29708
rect 16540 29696 16546 29708
rect 17678 29696 17684 29708
rect 16540 29668 17684 29696
rect 16540 29656 16546 29668
rect 17678 29656 17684 29668
rect 17736 29656 17742 29708
rect 17880 29668 19840 29696
rect 17880 29640 17908 29668
rect 15749 29631 15807 29637
rect 15749 29597 15761 29631
rect 15795 29597 15807 29631
rect 15749 29591 15807 29597
rect 15933 29631 15991 29637
rect 15933 29597 15945 29631
rect 15979 29628 15991 29631
rect 16577 29631 16635 29637
rect 16577 29628 16589 29631
rect 15979 29600 16589 29628
rect 15979 29597 15991 29600
rect 15933 29591 15991 29597
rect 16577 29597 16589 29600
rect 16623 29597 16635 29631
rect 17586 29628 17592 29640
rect 17547 29600 17592 29628
rect 16577 29591 16635 29597
rect 15764 29560 15792 29591
rect 17586 29588 17592 29600
rect 17644 29588 17650 29640
rect 17862 29628 17868 29640
rect 17823 29600 17868 29628
rect 17862 29588 17868 29600
rect 17920 29588 17926 29640
rect 17957 29631 18015 29637
rect 17957 29597 17969 29631
rect 18003 29597 18015 29631
rect 17957 29591 18015 29597
rect 16390 29560 16396 29572
rect 15764 29532 16396 29560
rect 16390 29520 16396 29532
rect 16448 29520 16454 29572
rect 14182 29452 14188 29504
rect 14240 29492 14246 29504
rect 14277 29495 14335 29501
rect 14277 29492 14289 29495
rect 14240 29464 14289 29492
rect 14240 29452 14246 29464
rect 14277 29461 14289 29464
rect 14323 29461 14335 29495
rect 14277 29455 14335 29461
rect 17402 29452 17408 29504
rect 17460 29492 17466 29504
rect 17972 29492 18000 29591
rect 18322 29588 18328 29640
rect 18380 29628 18386 29640
rect 19812 29637 19840 29668
rect 30650 29656 30656 29708
rect 30708 29696 30714 29708
rect 30745 29699 30803 29705
rect 30745 29696 30757 29699
rect 30708 29668 30757 29696
rect 30708 29656 30714 29668
rect 30745 29665 30757 29668
rect 30791 29696 30803 29699
rect 31481 29699 31539 29705
rect 31481 29696 31493 29699
rect 30791 29668 31493 29696
rect 30791 29665 30803 29668
rect 30745 29659 30803 29665
rect 31481 29665 31493 29668
rect 31527 29696 31539 29699
rect 31846 29696 31852 29708
rect 31527 29668 31852 29696
rect 31527 29665 31539 29668
rect 31481 29659 31539 29665
rect 31846 29656 31852 29668
rect 31904 29656 31910 29708
rect 19429 29631 19487 29637
rect 19429 29628 19441 29631
rect 18380 29600 19441 29628
rect 18380 29588 18386 29600
rect 19429 29597 19441 29600
rect 19475 29597 19487 29631
rect 19429 29591 19487 29597
rect 19797 29631 19855 29637
rect 19797 29597 19809 29631
rect 19843 29597 19855 29631
rect 20438 29628 20444 29640
rect 20399 29600 20444 29628
rect 19797 29591 19855 29597
rect 20438 29588 20444 29600
rect 20496 29588 20502 29640
rect 25682 29628 25688 29640
rect 25643 29600 25688 29628
rect 25682 29588 25688 29600
rect 25740 29588 25746 29640
rect 25958 29637 25964 29640
rect 25952 29628 25964 29637
rect 25919 29600 25964 29628
rect 25952 29591 25964 29600
rect 25958 29588 25964 29591
rect 26016 29588 26022 29640
rect 27706 29588 27712 29640
rect 27764 29628 27770 29640
rect 27893 29631 27951 29637
rect 27893 29628 27905 29631
rect 27764 29600 27905 29628
rect 27764 29588 27770 29600
rect 27893 29597 27905 29600
rect 27939 29628 27951 29631
rect 28721 29631 28779 29637
rect 28721 29628 28733 29631
rect 27939 29600 28733 29628
rect 27939 29597 27951 29600
rect 27893 29591 27951 29597
rect 28721 29597 28733 29600
rect 28767 29597 28779 29631
rect 28902 29628 28908 29640
rect 28863 29600 28908 29628
rect 28721 29591 28779 29597
rect 28902 29588 28908 29600
rect 28960 29588 28966 29640
rect 30466 29628 30472 29640
rect 30427 29600 30472 29628
rect 30466 29588 30472 29600
rect 30524 29588 30530 29640
rect 30558 29588 30564 29640
rect 30616 29628 30622 29640
rect 30616 29600 30661 29628
rect 30616 29588 30622 29600
rect 31018 29588 31024 29640
rect 31076 29628 31082 29640
rect 31205 29631 31263 29637
rect 31205 29628 31217 29631
rect 31076 29600 31217 29628
rect 31076 29588 31082 29600
rect 31205 29597 31217 29600
rect 31251 29597 31263 29631
rect 31205 29591 31263 29597
rect 32769 29631 32827 29637
rect 32769 29597 32781 29631
rect 32815 29628 32827 29631
rect 34790 29628 34796 29640
rect 32815 29600 34796 29628
rect 32815 29597 32827 29600
rect 32769 29591 32827 29597
rect 34790 29588 34796 29600
rect 34848 29588 34854 29640
rect 34900 29637 34928 29804
rect 43346 29792 43352 29804
rect 43404 29792 43410 29844
rect 42702 29696 42708 29708
rect 42663 29668 42708 29696
rect 42702 29656 42708 29668
rect 42760 29656 42766 29708
rect 43990 29696 43996 29708
rect 43951 29668 43996 29696
rect 43990 29656 43996 29668
rect 44048 29656 44054 29708
rect 44174 29696 44180 29708
rect 44135 29668 44180 29696
rect 44174 29656 44180 29668
rect 44232 29656 44238 29708
rect 34885 29631 34943 29637
rect 34885 29597 34897 29631
rect 34931 29597 34943 29631
rect 34885 29591 34943 29597
rect 36653 29631 36711 29637
rect 36653 29597 36665 29631
rect 36699 29628 36711 29631
rect 36814 29628 36820 29640
rect 36699 29600 36820 29628
rect 36699 29597 36711 29600
rect 36653 29591 36711 29597
rect 36814 29588 36820 29600
rect 36872 29588 36878 29640
rect 36909 29631 36967 29637
rect 36909 29597 36921 29631
rect 36955 29628 36967 29631
rect 37182 29628 37188 29640
rect 36955 29600 37188 29628
rect 36955 29597 36967 29600
rect 36909 29591 36967 29597
rect 37182 29588 37188 29600
rect 37240 29588 37246 29640
rect 18414 29520 18420 29572
rect 18472 29560 18478 29572
rect 18966 29560 18972 29572
rect 18472 29532 18972 29560
rect 18472 29520 18478 29532
rect 18966 29520 18972 29532
rect 19024 29560 19030 29572
rect 19521 29563 19579 29569
rect 19521 29560 19533 29563
rect 19024 29532 19533 29560
rect 19024 29520 19030 29532
rect 19521 29529 19533 29532
rect 19567 29529 19579 29563
rect 19521 29523 19579 29529
rect 19613 29563 19671 29569
rect 19613 29529 19625 29563
rect 19659 29529 19671 29563
rect 19613 29523 19671 29529
rect 19628 29492 19656 29523
rect 25222 29520 25228 29572
rect 25280 29560 25286 29572
rect 26418 29560 26424 29572
rect 25280 29532 26424 29560
rect 25280 29520 25286 29532
rect 26418 29520 26424 29532
rect 26476 29520 26482 29572
rect 28077 29563 28135 29569
rect 28077 29529 28089 29563
rect 28123 29560 28135 29563
rect 28920 29560 28948 29588
rect 28123 29532 28948 29560
rect 28123 29529 28135 29532
rect 28077 29523 28135 29529
rect 30374 29520 30380 29572
rect 30432 29560 30438 29572
rect 33318 29560 33324 29572
rect 30432 29532 33324 29560
rect 30432 29520 30438 29532
rect 33318 29520 33324 29532
rect 33376 29520 33382 29572
rect 33870 29520 33876 29572
rect 33928 29560 33934 29572
rect 34057 29563 34115 29569
rect 34057 29560 34069 29563
rect 33928 29532 34069 29560
rect 33928 29520 33934 29532
rect 34057 29529 34069 29532
rect 34103 29529 34115 29563
rect 34057 29523 34115 29529
rect 34977 29563 35035 29569
rect 34977 29529 34989 29563
rect 35023 29560 35035 29563
rect 35618 29560 35624 29572
rect 35023 29532 35624 29560
rect 35023 29529 35035 29532
rect 34977 29523 35035 29529
rect 35618 29520 35624 29532
rect 35676 29520 35682 29572
rect 17460 29464 19656 29492
rect 27065 29495 27123 29501
rect 17460 29452 17466 29464
rect 27065 29461 27077 29495
rect 27111 29492 27123 29495
rect 27430 29492 27436 29504
rect 27111 29464 27436 29492
rect 27111 29461 27123 29464
rect 27065 29455 27123 29461
rect 27430 29452 27436 29464
rect 27488 29452 27494 29504
rect 32677 29495 32735 29501
rect 32677 29461 32689 29495
rect 32723 29492 32735 29495
rect 32766 29492 32772 29504
rect 32723 29464 32772 29492
rect 32723 29461 32735 29464
rect 32677 29455 32735 29461
rect 32766 29452 32772 29464
rect 32824 29452 32830 29504
rect 33226 29452 33232 29504
rect 33284 29492 33290 29504
rect 33505 29495 33563 29501
rect 33505 29492 33517 29495
rect 33284 29464 33517 29492
rect 33284 29452 33290 29464
rect 33505 29461 33517 29464
rect 33551 29461 33563 29495
rect 33505 29455 33563 29461
rect 33597 29495 33655 29501
rect 33597 29461 33609 29495
rect 33643 29492 33655 29495
rect 33686 29492 33692 29504
rect 33643 29464 33692 29492
rect 33643 29461 33655 29464
rect 33597 29455 33655 29461
rect 33686 29452 33692 29464
rect 33744 29452 33750 29504
rect 35529 29495 35587 29501
rect 35529 29461 35541 29495
rect 35575 29492 35587 29495
rect 35802 29492 35808 29504
rect 35575 29464 35808 29492
rect 35575 29461 35587 29464
rect 35529 29455 35587 29461
rect 35802 29452 35808 29464
rect 35860 29452 35866 29504
rect 1104 29402 44896 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 44896 29402
rect 1104 29328 44896 29350
rect 13906 29248 13912 29300
rect 13964 29248 13970 29300
rect 17865 29291 17923 29297
rect 17865 29257 17877 29291
rect 17911 29288 17923 29291
rect 17954 29288 17960 29300
rect 17911 29260 17960 29288
rect 17911 29257 17923 29260
rect 17865 29251 17923 29257
rect 17954 29248 17960 29260
rect 18012 29248 18018 29300
rect 18138 29248 18144 29300
rect 18196 29288 18202 29300
rect 18877 29291 18935 29297
rect 18877 29288 18889 29291
rect 18196 29260 18889 29288
rect 18196 29248 18202 29260
rect 18877 29257 18889 29260
rect 18923 29257 18935 29291
rect 18877 29251 18935 29257
rect 18966 29248 18972 29300
rect 19024 29288 19030 29300
rect 19426 29288 19432 29300
rect 19024 29260 19432 29288
rect 19024 29248 19030 29260
rect 19426 29248 19432 29260
rect 19484 29288 19490 29300
rect 29546 29288 29552 29300
rect 19484 29260 25544 29288
rect 29507 29260 29552 29288
rect 19484 29248 19490 29260
rect 13924 29220 13952 29248
rect 14274 29220 14280 29232
rect 13648 29192 14280 29220
rect 13648 29161 13676 29192
rect 14274 29180 14280 29192
rect 14332 29180 14338 29232
rect 19334 29220 19340 29232
rect 18156 29192 19340 29220
rect 13633 29155 13691 29161
rect 13633 29121 13645 29155
rect 13679 29121 13691 29155
rect 13633 29115 13691 29121
rect 13900 29155 13958 29161
rect 13900 29121 13912 29155
rect 13946 29152 13958 29155
rect 14182 29152 14188 29164
rect 13946 29124 14188 29152
rect 13946 29121 13958 29124
rect 13900 29115 13958 29121
rect 14182 29112 14188 29124
rect 14240 29112 14246 29164
rect 17034 29152 17040 29164
rect 16995 29124 17040 29152
rect 17034 29112 17040 29124
rect 17092 29112 17098 29164
rect 18156 29161 18184 29192
rect 19334 29180 19340 29192
rect 19392 29180 19398 29232
rect 21266 29180 21272 29232
rect 21324 29220 21330 29232
rect 24578 29220 24584 29232
rect 21324 29192 24584 29220
rect 21324 29180 21330 29192
rect 24578 29180 24584 29192
rect 24636 29180 24642 29232
rect 25240 29229 25268 29260
rect 25225 29223 25283 29229
rect 25225 29189 25237 29223
rect 25271 29189 25283 29223
rect 25225 29183 25283 29189
rect 25314 29180 25320 29232
rect 25372 29220 25378 29232
rect 25425 29223 25483 29229
rect 25425 29220 25437 29223
rect 25372 29192 25437 29220
rect 25372 29180 25378 29192
rect 25425 29189 25437 29192
rect 25471 29189 25483 29223
rect 25516 29220 25544 29260
rect 29546 29248 29552 29260
rect 29604 29248 29610 29300
rect 30466 29248 30472 29300
rect 30524 29288 30530 29300
rect 30561 29291 30619 29297
rect 30561 29288 30573 29291
rect 30524 29260 30573 29288
rect 30524 29248 30530 29260
rect 30561 29257 30573 29260
rect 30607 29257 30619 29291
rect 30561 29251 30619 29257
rect 31573 29291 31631 29297
rect 31573 29257 31585 29291
rect 31619 29288 31631 29291
rect 32306 29288 32312 29300
rect 31619 29260 32312 29288
rect 31619 29257 31631 29260
rect 31573 29251 31631 29257
rect 32306 29248 32312 29260
rect 32364 29248 32370 29300
rect 43714 29288 43720 29300
rect 35912 29260 43720 29288
rect 35912 29220 35940 29260
rect 43714 29248 43720 29260
rect 43772 29248 43778 29300
rect 25516 29192 35940 29220
rect 25425 29183 25483 29189
rect 35986 29180 35992 29232
rect 36044 29220 36050 29232
rect 36044 29192 36676 29220
rect 36044 29180 36050 29192
rect 18049 29155 18107 29161
rect 18049 29121 18061 29155
rect 18095 29121 18107 29155
rect 18049 29115 18107 29121
rect 18141 29155 18199 29161
rect 18141 29121 18153 29155
rect 18187 29121 18199 29155
rect 18414 29152 18420 29164
rect 18375 29124 18420 29152
rect 18141 29115 18199 29121
rect 17310 29084 17316 29096
rect 17271 29056 17316 29084
rect 17310 29044 17316 29056
rect 17368 29044 17374 29096
rect 18064 29084 18092 29115
rect 18414 29112 18420 29124
rect 18472 29112 18478 29164
rect 18874 29152 18880 29164
rect 18835 29124 18880 29152
rect 18874 29112 18880 29124
rect 18932 29112 18938 29164
rect 19058 29152 19064 29164
rect 19019 29124 19064 29152
rect 19058 29112 19064 29124
rect 19116 29112 19122 29164
rect 20257 29155 20315 29161
rect 20257 29121 20269 29155
rect 20303 29152 20315 29155
rect 20438 29152 20444 29164
rect 20303 29124 20444 29152
rect 20303 29121 20315 29124
rect 20257 29115 20315 29121
rect 20438 29112 20444 29124
rect 20496 29112 20502 29164
rect 21726 29112 21732 29164
rect 21784 29152 21790 29164
rect 22077 29155 22135 29161
rect 22077 29152 22089 29155
rect 21784 29124 22089 29152
rect 21784 29112 21790 29124
rect 22077 29121 22089 29124
rect 22123 29121 22135 29155
rect 22077 29115 22135 29121
rect 28813 29155 28871 29161
rect 28813 29121 28825 29155
rect 28859 29152 28871 29155
rect 28902 29152 28908 29164
rect 28859 29124 28908 29152
rect 28859 29121 28871 29124
rect 28813 29115 28871 29121
rect 28902 29112 28908 29124
rect 28960 29112 28966 29164
rect 29457 29155 29515 29161
rect 29457 29121 29469 29155
rect 29503 29121 29515 29155
rect 29457 29115 29515 29121
rect 29641 29155 29699 29161
rect 29641 29121 29653 29155
rect 29687 29152 29699 29155
rect 29687 29124 30420 29152
rect 29687 29121 29699 29124
rect 29641 29115 29699 29121
rect 18230 29084 18236 29096
rect 18064 29056 18236 29084
rect 18230 29044 18236 29056
rect 18288 29084 18294 29096
rect 19242 29084 19248 29096
rect 18288 29056 19248 29084
rect 18288 29044 18294 29056
rect 19242 29044 19248 29056
rect 19300 29044 19306 29096
rect 21818 29084 21824 29096
rect 21779 29056 21824 29084
rect 21818 29044 21824 29056
rect 21876 29044 21882 29096
rect 29472 29084 29500 29115
rect 30101 29087 30159 29093
rect 30101 29084 30113 29087
rect 25608 29056 30113 29084
rect 15013 29019 15071 29025
rect 15013 28985 15025 29019
rect 15059 29016 15071 29019
rect 15194 29016 15200 29028
rect 15059 28988 15200 29016
rect 15059 28985 15071 28988
rect 15013 28979 15071 28985
rect 15194 28976 15200 28988
rect 15252 28976 15258 29028
rect 16666 28976 16672 29028
rect 16724 29016 16730 29028
rect 16853 29019 16911 29025
rect 16853 29016 16865 29019
rect 16724 28988 16865 29016
rect 16724 28976 16730 28988
rect 16853 28985 16865 28988
rect 16899 28985 16911 29019
rect 16853 28979 16911 28985
rect 17862 28976 17868 29028
rect 17920 29016 17926 29028
rect 18322 29016 18328 29028
rect 17920 28988 18328 29016
rect 17920 28976 17926 28988
rect 18322 28976 18328 28988
rect 18380 28976 18386 29028
rect 20073 29019 20131 29025
rect 20073 28985 20085 29019
rect 20119 29016 20131 29019
rect 20530 29016 20536 29028
rect 20119 28988 20536 29016
rect 20119 28985 20131 28988
rect 20073 28979 20131 28985
rect 20530 28976 20536 28988
rect 20588 29016 20594 29028
rect 20898 29016 20904 29028
rect 20588 28988 20904 29016
rect 20588 28976 20594 28988
rect 20898 28976 20904 28988
rect 20956 28976 20962 29028
rect 24210 29016 24216 29028
rect 24171 28988 24216 29016
rect 24210 28976 24216 28988
rect 24268 28976 24274 29028
rect 24765 29019 24823 29025
rect 24765 28985 24777 29019
rect 24811 29016 24823 29019
rect 24854 29016 24860 29028
rect 24811 28988 24860 29016
rect 24811 28985 24823 28988
rect 24765 28979 24823 28985
rect 24854 28976 24860 28988
rect 24912 28976 24918 29028
rect 25608 29025 25636 29056
rect 30101 29053 30113 29056
rect 30147 29053 30159 29087
rect 30392 29084 30420 29124
rect 30466 29112 30472 29164
rect 30524 29152 30530 29164
rect 31113 29155 31171 29161
rect 31113 29152 31125 29155
rect 30524 29124 31125 29152
rect 30524 29112 30530 29124
rect 31113 29121 31125 29124
rect 31159 29121 31171 29155
rect 31113 29115 31171 29121
rect 31205 29155 31263 29161
rect 31205 29121 31217 29155
rect 31251 29152 31263 29155
rect 31478 29152 31484 29164
rect 31251 29124 31484 29152
rect 31251 29121 31263 29124
rect 31205 29115 31263 29121
rect 31478 29112 31484 29124
rect 31536 29112 31542 29164
rect 31662 29112 31668 29164
rect 31720 29152 31726 29164
rect 32309 29155 32367 29161
rect 32309 29152 32321 29155
rect 31720 29124 32321 29152
rect 31720 29112 31726 29124
rect 32309 29121 32321 29124
rect 32355 29121 32367 29155
rect 32309 29115 32367 29121
rect 32493 29155 32551 29161
rect 32493 29121 32505 29155
rect 32539 29152 32551 29155
rect 32582 29152 32588 29164
rect 32539 29124 32588 29152
rect 32539 29121 32551 29124
rect 32493 29115 32551 29121
rect 32582 29112 32588 29124
rect 32640 29112 32646 29164
rect 33318 29112 33324 29164
rect 33376 29152 33382 29164
rect 33505 29155 33563 29161
rect 33505 29152 33517 29155
rect 33376 29124 33517 29152
rect 33376 29112 33382 29124
rect 33505 29121 33517 29124
rect 33551 29121 33563 29155
rect 33870 29152 33876 29164
rect 33831 29124 33876 29152
rect 33505 29115 33563 29121
rect 33870 29112 33876 29124
rect 33928 29112 33934 29164
rect 33962 29112 33968 29164
rect 34020 29152 34026 29164
rect 34020 29124 34065 29152
rect 34020 29112 34026 29124
rect 35526 29112 35532 29164
rect 35584 29152 35590 29164
rect 35802 29152 35808 29164
rect 35584 29124 35808 29152
rect 35584 29112 35590 29124
rect 35802 29112 35808 29124
rect 35860 29152 35866 29164
rect 36648 29161 36676 29192
rect 36449 29155 36507 29161
rect 36449 29152 36461 29155
rect 35860 29124 36461 29152
rect 35860 29112 35866 29124
rect 36449 29121 36461 29124
rect 36495 29121 36507 29155
rect 36449 29115 36507 29121
rect 36633 29155 36691 29161
rect 36633 29121 36645 29155
rect 36679 29121 36691 29155
rect 36633 29115 36691 29121
rect 30392 29056 30696 29084
rect 30101 29047 30159 29053
rect 25593 29019 25651 29025
rect 25593 28985 25605 29019
rect 25639 28985 25651 29019
rect 28718 29016 28724 29028
rect 28679 28988 28724 29016
rect 25593 28979 25651 28985
rect 28718 28976 28724 28988
rect 28776 28976 28782 29028
rect 30116 29016 30144 29047
rect 30374 29016 30380 29028
rect 30116 28988 30236 29016
rect 30335 28988 30380 29016
rect 17218 28948 17224 28960
rect 17179 28920 17224 28948
rect 17218 28908 17224 28920
rect 17276 28908 17282 28960
rect 23198 28948 23204 28960
rect 23159 28920 23204 28948
rect 23198 28908 23204 28920
rect 23256 28948 23262 28960
rect 24581 28951 24639 28957
rect 24581 28948 24593 28951
rect 23256 28920 24593 28948
rect 23256 28908 23262 28920
rect 24581 28917 24593 28920
rect 24627 28917 24639 28951
rect 25406 28948 25412 28960
rect 25367 28920 25412 28948
rect 24581 28911 24639 28917
rect 25406 28908 25412 28920
rect 25464 28908 25470 28960
rect 30208 28948 30236 28988
rect 30374 28976 30380 28988
rect 30432 28976 30438 29028
rect 30466 28948 30472 28960
rect 30208 28920 30472 28948
rect 30466 28908 30472 28920
rect 30524 28908 30530 28960
rect 30668 28948 30696 29056
rect 30742 29044 30748 29096
rect 30800 29084 30806 29096
rect 31294 29084 31300 29096
rect 30800 29056 31300 29084
rect 30800 29044 30806 29056
rect 31294 29044 31300 29056
rect 31352 29044 31358 29096
rect 31389 29087 31447 29093
rect 31389 29053 31401 29087
rect 31435 29053 31447 29087
rect 31496 29084 31524 29112
rect 33226 29084 33232 29096
rect 31496 29056 33232 29084
rect 31389 29047 31447 29053
rect 31404 29016 31432 29047
rect 33226 29044 33232 29056
rect 33284 29044 33290 29096
rect 31570 29016 31576 29028
rect 31404 28988 31576 29016
rect 31570 28976 31576 28988
rect 31628 28976 31634 29028
rect 32582 29016 32588 29028
rect 31956 28988 32588 29016
rect 31956 28948 31984 28988
rect 32582 28976 32588 28988
rect 32640 28976 32646 29028
rect 33244 29016 33272 29044
rect 33962 29016 33968 29028
rect 33244 28988 33968 29016
rect 33962 28976 33968 28988
rect 34020 28976 34026 29028
rect 34149 29019 34207 29025
rect 34149 28985 34161 29019
rect 34195 29016 34207 29019
rect 34790 29016 34796 29028
rect 34195 28988 34796 29016
rect 34195 28985 34207 28988
rect 34149 28979 34207 28985
rect 34790 28976 34796 28988
rect 34848 28976 34854 29028
rect 32122 28948 32128 28960
rect 30668 28920 31984 28948
rect 32083 28920 32128 28948
rect 32122 28908 32128 28920
rect 32180 28908 32186 28960
rect 32306 28908 32312 28960
rect 32364 28948 32370 28960
rect 33597 28951 33655 28957
rect 33597 28948 33609 28951
rect 32364 28920 33609 28948
rect 32364 28908 32370 28920
rect 33597 28917 33609 28920
rect 33643 28948 33655 28951
rect 33686 28948 33692 28960
rect 33643 28920 33692 28948
rect 33643 28917 33655 28920
rect 33597 28911 33655 28917
rect 33686 28908 33692 28920
rect 33744 28908 33750 28960
rect 35621 28951 35679 28957
rect 35621 28917 35633 28951
rect 35667 28948 35679 28951
rect 35710 28948 35716 28960
rect 35667 28920 35716 28948
rect 35667 28917 35679 28920
rect 35621 28911 35679 28917
rect 35710 28908 35716 28920
rect 35768 28908 35774 28960
rect 36538 28948 36544 28960
rect 36499 28920 36544 28948
rect 36538 28908 36544 28920
rect 36596 28908 36602 28960
rect 1104 28858 44896 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 44896 28858
rect 1104 28784 44896 28806
rect 15194 28704 15200 28756
rect 15252 28744 15258 28756
rect 16482 28744 16488 28756
rect 15252 28716 16488 28744
rect 15252 28704 15258 28716
rect 16482 28704 16488 28716
rect 16540 28744 16546 28756
rect 21266 28744 21272 28756
rect 16540 28716 17816 28744
rect 16540 28704 16546 28716
rect 15657 28679 15715 28685
rect 15657 28645 15669 28679
rect 15703 28676 15715 28679
rect 16390 28676 16396 28688
rect 15703 28648 16396 28676
rect 15703 28645 15715 28648
rect 15657 28639 15715 28645
rect 16390 28636 16396 28648
rect 16448 28676 16454 28688
rect 17310 28676 17316 28688
rect 16448 28648 17316 28676
rect 16448 28636 16454 28648
rect 16500 28617 16528 28648
rect 17310 28636 17316 28648
rect 17368 28676 17374 28688
rect 17681 28679 17739 28685
rect 17681 28676 17693 28679
rect 17368 28648 17693 28676
rect 17368 28636 17374 28648
rect 17681 28645 17693 28648
rect 17727 28645 17739 28679
rect 17681 28639 17739 28645
rect 16485 28611 16543 28617
rect 16485 28577 16497 28611
rect 16531 28577 16543 28611
rect 16485 28571 16543 28577
rect 16850 28568 16856 28620
rect 16908 28608 16914 28620
rect 17218 28608 17224 28620
rect 16908 28580 17224 28608
rect 16908 28568 16914 28580
rect 17218 28568 17224 28580
rect 17276 28608 17282 28620
rect 17589 28611 17647 28617
rect 17589 28608 17601 28611
rect 17276 28580 17601 28608
rect 17276 28568 17282 28580
rect 17589 28577 17601 28580
rect 17635 28577 17647 28611
rect 17589 28571 17647 28577
rect 14274 28540 14280 28552
rect 14235 28512 14280 28540
rect 14274 28500 14280 28512
rect 14332 28500 14338 28552
rect 16574 28500 16580 28552
rect 16632 28540 16638 28552
rect 17494 28540 17500 28552
rect 16632 28512 16677 28540
rect 17407 28512 17500 28540
rect 16632 28500 16638 28512
rect 17494 28500 17500 28512
rect 17552 28500 17558 28552
rect 17788 28549 17816 28716
rect 17880 28716 20852 28744
rect 21227 28716 21272 28744
rect 17773 28543 17831 28549
rect 17773 28509 17785 28543
rect 17819 28509 17831 28543
rect 17773 28503 17831 28509
rect 14544 28475 14602 28481
rect 14544 28441 14556 28475
rect 14590 28472 14602 28475
rect 16761 28475 16819 28481
rect 16761 28472 16773 28475
rect 14590 28444 16773 28472
rect 14590 28441 14602 28444
rect 14544 28435 14602 28441
rect 16761 28441 16773 28444
rect 16807 28441 16819 28475
rect 17512 28472 17540 28500
rect 17880 28472 17908 28716
rect 20824 28676 20852 28716
rect 21266 28704 21272 28716
rect 21324 28704 21330 28756
rect 21913 28747 21971 28753
rect 21913 28713 21925 28747
rect 21959 28744 21971 28747
rect 22186 28744 22192 28756
rect 21959 28716 22192 28744
rect 21959 28713 21971 28716
rect 21913 28707 21971 28713
rect 22186 28704 22192 28716
rect 22244 28704 22250 28756
rect 27706 28744 27712 28756
rect 27667 28716 27712 28744
rect 27706 28704 27712 28716
rect 27764 28704 27770 28756
rect 27890 28744 27896 28756
rect 27851 28716 27896 28744
rect 27890 28704 27896 28716
rect 27948 28704 27954 28756
rect 30466 28704 30472 28756
rect 30524 28744 30530 28756
rect 31294 28744 31300 28756
rect 30524 28716 31300 28744
rect 30524 28704 30530 28716
rect 31294 28704 31300 28716
rect 31352 28744 31358 28756
rect 31662 28744 31668 28756
rect 31352 28716 31668 28744
rect 31352 28704 31358 28716
rect 31662 28704 31668 28716
rect 31720 28704 31726 28756
rect 34977 28747 35035 28753
rect 34977 28744 34989 28747
rect 34900 28716 34989 28744
rect 34900 28688 34928 28716
rect 34977 28713 34989 28716
rect 35023 28744 35035 28747
rect 35526 28744 35532 28756
rect 35023 28716 35532 28744
rect 35023 28713 35035 28716
rect 34977 28707 35035 28713
rect 35526 28704 35532 28716
rect 35584 28704 35590 28756
rect 35710 28744 35716 28756
rect 35671 28716 35716 28744
rect 35710 28704 35716 28716
rect 35768 28704 35774 28756
rect 35897 28747 35955 28753
rect 35897 28713 35909 28747
rect 35943 28744 35955 28747
rect 37458 28744 37464 28756
rect 35943 28716 37464 28744
rect 35943 28713 35955 28716
rect 35897 28707 35955 28713
rect 37458 28704 37464 28716
rect 37516 28704 37522 28756
rect 25406 28676 25412 28688
rect 20824 28648 25412 28676
rect 25406 28636 25412 28648
rect 25464 28636 25470 28688
rect 25774 28676 25780 28688
rect 25735 28648 25780 28676
rect 25774 28636 25780 28648
rect 25832 28636 25838 28688
rect 34882 28636 34888 28688
rect 34940 28636 34946 28688
rect 17957 28611 18015 28617
rect 17957 28577 17969 28611
rect 18003 28608 18015 28611
rect 18509 28611 18567 28617
rect 18509 28608 18521 28611
rect 18003 28580 18521 28608
rect 18003 28577 18015 28580
rect 17957 28571 18015 28577
rect 18509 28577 18521 28580
rect 18555 28577 18567 28611
rect 18509 28571 18567 28577
rect 18693 28611 18751 28617
rect 18693 28577 18705 28611
rect 18739 28608 18751 28611
rect 19058 28608 19064 28620
rect 18739 28580 19064 28608
rect 18739 28577 18751 28580
rect 18693 28571 18751 28577
rect 19058 28568 19064 28580
rect 19116 28568 19122 28620
rect 22646 28568 22652 28620
rect 22704 28608 22710 28620
rect 22704 28580 23152 28608
rect 22704 28568 22710 28580
rect 18322 28500 18328 28552
rect 18380 28540 18386 28552
rect 18417 28543 18475 28549
rect 18417 28540 18429 28543
rect 18380 28512 18429 28540
rect 18380 28500 18386 28512
rect 18417 28509 18429 28512
rect 18463 28509 18475 28543
rect 18417 28503 18475 28509
rect 19889 28543 19947 28549
rect 19889 28509 19901 28543
rect 19935 28540 19947 28543
rect 21818 28540 21824 28552
rect 19935 28512 21824 28540
rect 19935 28509 19947 28512
rect 19889 28503 19947 28509
rect 21818 28500 21824 28512
rect 21876 28500 21882 28552
rect 22278 28540 22284 28552
rect 22239 28512 22284 28540
rect 22278 28500 22284 28512
rect 22336 28500 22342 28552
rect 22833 28543 22891 28549
rect 22833 28509 22845 28543
rect 22879 28509 22891 28543
rect 23014 28540 23020 28552
rect 22975 28512 23020 28540
rect 22833 28503 22891 28509
rect 17512 28444 17908 28472
rect 20156 28475 20214 28481
rect 16761 28435 16819 28441
rect 20156 28441 20168 28475
rect 20202 28472 20214 28475
rect 20714 28472 20720 28484
rect 20202 28444 20720 28472
rect 20202 28441 20214 28444
rect 20156 28435 20214 28441
rect 20714 28432 20720 28444
rect 20772 28432 20778 28484
rect 22848 28472 22876 28503
rect 23014 28500 23020 28512
rect 23072 28500 23078 28552
rect 23124 28549 23152 28580
rect 24210 28568 24216 28620
rect 24268 28608 24274 28620
rect 24397 28611 24455 28617
rect 24397 28608 24409 28611
rect 24268 28580 24409 28608
rect 24268 28568 24274 28580
rect 24397 28577 24409 28580
rect 24443 28577 24455 28611
rect 24397 28571 24455 28577
rect 24854 28568 24860 28620
rect 24912 28608 24918 28620
rect 26145 28611 26203 28617
rect 26145 28608 26157 28611
rect 24912 28580 26157 28608
rect 24912 28568 24918 28580
rect 26145 28577 26157 28580
rect 26191 28577 26203 28611
rect 26145 28571 26203 28577
rect 27982 28568 27988 28620
rect 28040 28608 28046 28620
rect 28534 28608 28540 28620
rect 28040 28580 28540 28608
rect 28040 28568 28046 28580
rect 28534 28568 28540 28580
rect 28592 28568 28598 28620
rect 30742 28608 30748 28620
rect 30208 28580 30748 28608
rect 23109 28543 23167 28549
rect 23109 28509 23121 28543
rect 23155 28509 23167 28543
rect 23109 28503 23167 28509
rect 23201 28543 23259 28549
rect 23201 28509 23213 28543
rect 23247 28540 23259 28543
rect 23290 28540 23296 28552
rect 23247 28512 23296 28540
rect 23247 28509 23259 28512
rect 23201 28503 23259 28509
rect 23290 28500 23296 28512
rect 23348 28540 23354 28552
rect 24673 28543 24731 28549
rect 24673 28540 24685 28543
rect 23348 28512 24685 28540
rect 23348 28500 23354 28512
rect 24673 28509 24685 28512
rect 24719 28509 24731 28543
rect 24673 28503 24731 28509
rect 26050 28500 26056 28552
rect 26108 28540 26114 28552
rect 26789 28543 26847 28549
rect 26789 28540 26801 28543
rect 26108 28512 26801 28540
rect 26108 28500 26114 28512
rect 26789 28509 26801 28512
rect 26835 28509 26847 28543
rect 27062 28540 27068 28552
rect 27023 28512 27068 28540
rect 26789 28503 26847 28509
rect 27062 28500 27068 28512
rect 27120 28500 27126 28552
rect 27338 28500 27344 28552
rect 27396 28540 27402 28552
rect 30208 28549 30236 28580
rect 30742 28568 30748 28580
rect 30800 28568 30806 28620
rect 30929 28611 30987 28617
rect 30929 28577 30941 28611
rect 30975 28608 30987 28611
rect 31202 28608 31208 28620
rect 30975 28580 31208 28608
rect 30975 28577 30987 28580
rect 30929 28571 30987 28577
rect 31202 28568 31208 28580
rect 31260 28568 31266 28620
rect 31297 28611 31355 28617
rect 31297 28577 31309 28611
rect 31343 28608 31355 28611
rect 32122 28608 32128 28620
rect 31343 28580 32128 28608
rect 31343 28577 31355 28580
rect 31297 28571 31355 28577
rect 32122 28568 32128 28580
rect 32180 28568 32186 28620
rect 33594 28608 33600 28620
rect 33555 28580 33600 28608
rect 33594 28568 33600 28580
rect 33652 28568 33658 28620
rect 34790 28568 34796 28620
rect 34848 28608 34854 28620
rect 34848 28580 35112 28608
rect 34848 28568 34854 28580
rect 28721 28543 28779 28549
rect 28721 28540 28733 28543
rect 27396 28512 28733 28540
rect 27396 28500 27402 28512
rect 28721 28509 28733 28512
rect 28767 28509 28779 28543
rect 28721 28503 28779 28509
rect 30193 28543 30251 28549
rect 30193 28509 30205 28543
rect 30239 28509 30251 28543
rect 30193 28503 30251 28509
rect 30469 28543 30527 28549
rect 30469 28509 30481 28543
rect 30515 28540 30527 28543
rect 30558 28540 30564 28552
rect 30515 28512 30564 28540
rect 30515 28509 30527 28512
rect 30469 28503 30527 28509
rect 30558 28500 30564 28512
rect 30616 28540 30622 28552
rect 31570 28540 31576 28552
rect 30616 28512 31576 28540
rect 30616 28500 30622 28512
rect 31570 28500 31576 28512
rect 31628 28540 31634 28552
rect 32033 28543 32091 28549
rect 32033 28540 32045 28543
rect 31628 28512 32045 28540
rect 31628 28500 31634 28512
rect 32033 28509 32045 28512
rect 32079 28509 32091 28543
rect 32033 28503 32091 28509
rect 32217 28543 32275 28549
rect 32217 28509 32229 28543
rect 32263 28509 32275 28543
rect 32217 28503 32275 28509
rect 26881 28475 26939 28481
rect 22066 28444 25728 28472
rect 16114 28404 16120 28416
rect 16075 28376 16120 28404
rect 16114 28364 16120 28376
rect 16172 28364 16178 28416
rect 18046 28364 18052 28416
rect 18104 28404 18110 28416
rect 18693 28407 18751 28413
rect 18693 28404 18705 28407
rect 18104 28376 18705 28404
rect 18104 28364 18110 28376
rect 18693 28373 18705 28376
rect 18739 28373 18751 28407
rect 18693 28367 18751 28373
rect 21634 28364 21640 28416
rect 21692 28404 21698 28416
rect 21729 28407 21787 28413
rect 21729 28404 21741 28407
rect 21692 28376 21741 28404
rect 21692 28364 21698 28376
rect 21729 28373 21741 28376
rect 21775 28373 21787 28407
rect 21910 28404 21916 28416
rect 21871 28376 21916 28404
rect 21729 28367 21787 28373
rect 21910 28364 21916 28376
rect 21968 28404 21974 28416
rect 22066 28404 22094 28444
rect 21968 28376 22094 28404
rect 21968 28364 21974 28376
rect 23382 28364 23388 28416
rect 23440 28404 23446 28416
rect 25700 28413 25728 28444
rect 26881 28441 26893 28475
rect 26927 28472 26939 28475
rect 27877 28475 27935 28481
rect 26927 28444 27844 28472
rect 26927 28441 26939 28444
rect 26881 28435 26939 28441
rect 23477 28407 23535 28413
rect 23477 28404 23489 28407
rect 23440 28376 23489 28404
rect 23440 28364 23446 28376
rect 23477 28373 23489 28376
rect 23523 28373 23535 28407
rect 23477 28367 23535 28373
rect 25685 28407 25743 28413
rect 25685 28373 25697 28407
rect 25731 28373 25743 28407
rect 25685 28367 25743 28373
rect 27249 28407 27307 28413
rect 27249 28373 27261 28407
rect 27295 28404 27307 28407
rect 27522 28404 27528 28416
rect 27295 28376 27528 28404
rect 27295 28373 27307 28376
rect 27249 28367 27307 28373
rect 27522 28364 27528 28376
rect 27580 28364 27586 28416
rect 27816 28404 27844 28444
rect 27877 28441 27889 28475
rect 27923 28472 27935 28475
rect 27982 28472 27988 28484
rect 27923 28444 27988 28472
rect 27923 28441 27935 28444
rect 27877 28435 27935 28441
rect 27982 28432 27988 28444
rect 28040 28432 28046 28484
rect 28077 28475 28135 28481
rect 28077 28441 28089 28475
rect 28123 28472 28135 28475
rect 28902 28472 28908 28484
rect 28123 28444 28908 28472
rect 28123 28441 28135 28444
rect 28077 28435 28135 28441
rect 28092 28404 28120 28435
rect 28902 28432 28908 28444
rect 28960 28432 28966 28484
rect 30009 28475 30067 28481
rect 30009 28441 30021 28475
rect 30055 28472 30067 28475
rect 31414 28475 31472 28481
rect 31414 28472 31426 28475
rect 30055 28444 31426 28472
rect 30055 28441 30067 28444
rect 30009 28435 30067 28441
rect 31414 28441 31426 28444
rect 31460 28441 31472 28475
rect 31414 28435 31472 28441
rect 31754 28432 31760 28484
rect 31812 28472 31818 28484
rect 31938 28472 31944 28484
rect 31812 28444 31944 28472
rect 31812 28432 31818 28444
rect 31938 28432 31944 28444
rect 31996 28472 32002 28484
rect 32232 28472 32260 28503
rect 32306 28500 32312 28552
rect 32364 28540 32370 28552
rect 33318 28540 33324 28552
rect 32364 28512 32409 28540
rect 33279 28512 33324 28540
rect 32364 28500 32370 28512
rect 33318 28500 33324 28512
rect 33376 28500 33382 28552
rect 35084 28549 35112 28580
rect 34977 28543 35035 28549
rect 34977 28509 34989 28543
rect 35023 28509 35035 28543
rect 34977 28503 35035 28509
rect 35069 28543 35127 28549
rect 35069 28509 35081 28543
rect 35115 28509 35127 28543
rect 35069 28503 35127 28509
rect 36449 28543 36507 28549
rect 36449 28509 36461 28543
rect 36495 28540 36507 28543
rect 37182 28540 37188 28552
rect 36495 28512 37188 28540
rect 36495 28509 36507 28512
rect 36449 28503 36507 28509
rect 34514 28472 34520 28484
rect 31996 28444 34520 28472
rect 31996 28432 32002 28444
rect 34514 28432 34520 28444
rect 34572 28432 34578 28484
rect 34992 28472 35020 28503
rect 37182 28500 37188 28512
rect 37240 28500 37246 28552
rect 43438 28540 43444 28552
rect 43399 28512 43444 28540
rect 43438 28500 43444 28512
rect 43496 28500 43502 28552
rect 35526 28472 35532 28484
rect 34992 28444 35103 28472
rect 35487 28444 35532 28472
rect 27816 28376 28120 28404
rect 28166 28364 28172 28416
rect 28224 28404 28230 28416
rect 28537 28407 28595 28413
rect 28537 28404 28549 28407
rect 28224 28376 28549 28404
rect 28224 28364 28230 28376
rect 28537 28373 28549 28376
rect 28583 28373 28595 28407
rect 28537 28367 28595 28373
rect 30377 28407 30435 28413
rect 30377 28373 30389 28407
rect 30423 28404 30435 28407
rect 31018 28404 31024 28416
rect 30423 28376 31024 28404
rect 30423 28373 30435 28376
rect 30377 28367 30435 28373
rect 31018 28364 31024 28376
rect 31076 28364 31082 28416
rect 31110 28364 31116 28416
rect 31168 28404 31174 28416
rect 31205 28407 31263 28413
rect 31205 28404 31217 28407
rect 31168 28376 31217 28404
rect 31168 28364 31174 28376
rect 31205 28373 31217 28376
rect 31251 28373 31263 28407
rect 31205 28367 31263 28373
rect 31573 28407 31631 28413
rect 31573 28373 31585 28407
rect 31619 28404 31631 28407
rect 32490 28404 32496 28416
rect 31619 28376 32496 28404
rect 31619 28373 31631 28376
rect 31573 28367 31631 28373
rect 32490 28364 32496 28376
rect 32548 28364 32554 28416
rect 32582 28364 32588 28416
rect 32640 28404 32646 28416
rect 34422 28404 34428 28416
rect 32640 28376 34428 28404
rect 32640 28364 32646 28376
rect 34422 28364 34428 28376
rect 34480 28404 34486 28416
rect 34701 28407 34759 28413
rect 34701 28404 34713 28407
rect 34480 28376 34713 28404
rect 34480 28364 34486 28376
rect 34701 28373 34713 28376
rect 34747 28373 34759 28407
rect 35075 28404 35103 28444
rect 35526 28432 35532 28444
rect 35584 28432 35590 28484
rect 35745 28475 35803 28481
rect 35745 28441 35757 28475
rect 35791 28472 35803 28475
rect 36078 28472 36084 28484
rect 35791 28444 36084 28472
rect 35791 28441 35803 28444
rect 35745 28435 35803 28441
rect 36078 28432 36084 28444
rect 36136 28472 36142 28484
rect 36538 28472 36544 28484
rect 36136 28444 36544 28472
rect 36136 28432 36142 28444
rect 36538 28432 36544 28444
rect 36596 28432 36602 28484
rect 36722 28481 36728 28484
rect 36716 28435 36728 28481
rect 36780 28472 36786 28484
rect 36780 28444 36816 28472
rect 36722 28432 36728 28435
rect 36780 28432 36786 28444
rect 36170 28404 36176 28416
rect 35075 28376 36176 28404
rect 34701 28367 34759 28373
rect 36170 28364 36176 28376
rect 36228 28364 36234 28416
rect 37458 28364 37464 28416
rect 37516 28404 37522 28416
rect 37829 28407 37887 28413
rect 37829 28404 37841 28407
rect 37516 28376 37841 28404
rect 37516 28364 37522 28376
rect 37829 28373 37841 28376
rect 37875 28373 37887 28407
rect 37829 28367 37887 28373
rect 43533 28407 43591 28413
rect 43533 28373 43545 28407
rect 43579 28404 43591 28407
rect 43990 28404 43996 28416
rect 43579 28376 43996 28404
rect 43579 28373 43591 28376
rect 43533 28367 43591 28373
rect 43990 28364 43996 28376
rect 44048 28364 44054 28416
rect 1104 28314 44896 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 44896 28314
rect 1104 28240 44896 28262
rect 14458 28160 14464 28212
rect 14516 28200 14522 28212
rect 14829 28203 14887 28209
rect 14829 28200 14841 28203
rect 14516 28172 14841 28200
rect 14516 28160 14522 28172
rect 14829 28169 14841 28172
rect 14875 28169 14887 28203
rect 14829 28163 14887 28169
rect 16025 28203 16083 28209
rect 16025 28169 16037 28203
rect 16071 28200 16083 28203
rect 17862 28200 17868 28212
rect 16071 28172 17868 28200
rect 16071 28169 16083 28172
rect 16025 28163 16083 28169
rect 17862 28160 17868 28172
rect 17920 28160 17926 28212
rect 21177 28203 21235 28209
rect 21177 28169 21189 28203
rect 21223 28200 21235 28203
rect 21266 28200 21272 28212
rect 21223 28172 21272 28200
rect 21223 28169 21235 28172
rect 21177 28163 21235 28169
rect 21266 28160 21272 28172
rect 21324 28160 21330 28212
rect 22186 28200 22192 28212
rect 22147 28172 22192 28200
rect 22186 28160 22192 28172
rect 22244 28160 22250 28212
rect 23198 28200 23204 28212
rect 22388 28172 23204 28200
rect 17034 28092 17040 28144
rect 17092 28132 17098 28144
rect 17497 28135 17555 28141
rect 17497 28132 17509 28135
rect 17092 28104 17509 28132
rect 17092 28092 17098 28104
rect 17497 28101 17509 28104
rect 17543 28132 17555 28135
rect 21910 28132 21916 28144
rect 17543 28104 19472 28132
rect 17543 28101 17555 28104
rect 17497 28095 17555 28101
rect 19444 28076 19472 28104
rect 20824 28104 21916 28132
rect 15013 28067 15071 28073
rect 15013 28033 15025 28067
rect 15059 28064 15071 28067
rect 16022 28064 16028 28076
rect 15059 28036 16028 28064
rect 15059 28033 15071 28036
rect 15013 28027 15071 28033
rect 16022 28024 16028 28036
rect 16080 28024 16086 28076
rect 16117 28067 16175 28073
rect 16117 28033 16129 28067
rect 16163 28064 16175 28067
rect 16850 28064 16856 28076
rect 16163 28036 16856 28064
rect 16163 28033 16175 28036
rect 16117 28027 16175 28033
rect 16850 28024 16856 28036
rect 16908 28024 16914 28076
rect 17313 28067 17371 28073
rect 17313 28033 17325 28067
rect 17359 28033 17371 28067
rect 17313 28027 17371 28033
rect 17589 28067 17647 28073
rect 17589 28033 17601 28067
rect 17635 28064 17647 28067
rect 17678 28064 17684 28076
rect 17635 28036 17684 28064
rect 17635 28033 17647 28036
rect 17589 28027 17647 28033
rect 15194 27996 15200 28008
rect 15155 27968 15200 27996
rect 15194 27956 15200 27968
rect 15252 27956 15258 28008
rect 17328 27996 17356 28027
rect 17678 28024 17684 28036
rect 17736 28024 17742 28076
rect 18046 28064 18052 28076
rect 18007 28036 18052 28064
rect 18046 28024 18052 28036
rect 18104 28024 18110 28076
rect 19426 28024 19432 28076
rect 19484 28064 19490 28076
rect 20824 28073 20852 28104
rect 21910 28092 21916 28104
rect 21968 28092 21974 28144
rect 19521 28067 19579 28073
rect 19521 28064 19533 28067
rect 19484 28036 19533 28064
rect 19484 28024 19490 28036
rect 19521 28033 19533 28036
rect 19567 28033 19579 28067
rect 19521 28027 19579 28033
rect 20809 28067 20867 28073
rect 20809 28033 20821 28067
rect 20855 28033 20867 28067
rect 20809 28027 20867 28033
rect 21269 28067 21327 28073
rect 21269 28033 21281 28067
rect 21315 28064 21327 28067
rect 22278 28064 22284 28076
rect 21315 28036 22284 28064
rect 21315 28033 21327 28036
rect 21269 28027 21327 28033
rect 22278 28024 22284 28036
rect 22336 28024 22342 28076
rect 22388 28073 22416 28172
rect 23198 28160 23204 28172
rect 23256 28160 23262 28212
rect 24210 28160 24216 28212
rect 24268 28200 24274 28212
rect 24489 28203 24547 28209
rect 24489 28200 24501 28203
rect 24268 28172 24501 28200
rect 24268 28160 24274 28172
rect 24489 28169 24501 28172
rect 24535 28169 24547 28203
rect 24489 28163 24547 28169
rect 25777 28203 25835 28209
rect 25777 28169 25789 28203
rect 25823 28169 25835 28203
rect 27338 28200 27344 28212
rect 27299 28172 27344 28200
rect 25777 28163 25835 28169
rect 22557 28135 22615 28141
rect 22557 28101 22569 28135
rect 22603 28132 22615 28135
rect 22738 28132 22744 28144
rect 22603 28104 22744 28132
rect 22603 28101 22615 28104
rect 22557 28095 22615 28101
rect 22738 28092 22744 28104
rect 22796 28092 22802 28144
rect 25682 28132 25688 28144
rect 23124 28104 25688 28132
rect 22373 28067 22431 28073
rect 22373 28033 22385 28067
rect 22419 28033 22431 28067
rect 22373 28027 22431 28033
rect 22646 28024 22652 28076
rect 22704 28064 22710 28076
rect 23124 28073 23152 28104
rect 25682 28092 25688 28104
rect 25740 28092 25746 28144
rect 23382 28073 23388 28076
rect 23109 28067 23167 28073
rect 22704 28036 22749 28064
rect 22704 28024 22710 28036
rect 23109 28033 23121 28067
rect 23155 28033 23167 28067
rect 23376 28064 23388 28073
rect 23343 28036 23388 28064
rect 23109 28027 23167 28033
rect 23376 28027 23388 28036
rect 23382 28024 23388 28027
rect 23440 28024 23446 28076
rect 25133 28067 25191 28073
rect 25133 28033 25145 28067
rect 25179 28064 25191 28067
rect 25792 28064 25820 28163
rect 27338 28160 27344 28172
rect 27396 28160 27402 28212
rect 27522 28200 27528 28212
rect 27483 28172 27528 28200
rect 27522 28160 27528 28172
rect 27580 28160 27586 28212
rect 29181 28203 29239 28209
rect 29181 28169 29193 28203
rect 29227 28169 29239 28203
rect 29181 28163 29239 28169
rect 30561 28203 30619 28209
rect 30561 28169 30573 28203
rect 30607 28200 30619 28203
rect 31202 28200 31208 28212
rect 30607 28172 31208 28200
rect 30607 28169 30619 28172
rect 30561 28163 30619 28169
rect 26053 28135 26111 28141
rect 26053 28101 26065 28135
rect 26099 28132 26111 28135
rect 29196 28132 29224 28163
rect 31202 28160 31208 28172
rect 31260 28160 31266 28212
rect 32582 28200 32588 28212
rect 32324 28172 32588 28200
rect 26099 28104 29224 28132
rect 30193 28135 30251 28141
rect 26099 28101 26111 28104
rect 26053 28095 26111 28101
rect 30193 28101 30205 28135
rect 30239 28101 30251 28135
rect 30393 28135 30451 28141
rect 30393 28132 30405 28135
rect 30193 28095 30251 28101
rect 30392 28101 30405 28132
rect 30439 28101 30451 28135
rect 30392 28095 30451 28101
rect 25179 28036 25820 28064
rect 26421 28067 26479 28073
rect 25179 28033 25191 28036
rect 25133 28027 25191 28033
rect 26421 28033 26433 28067
rect 26467 28064 26479 28067
rect 27062 28064 27068 28076
rect 26467 28036 27068 28064
rect 26467 28033 26479 28036
rect 26421 28027 26479 28033
rect 27062 28024 27068 28036
rect 27120 28064 27126 28076
rect 28353 28067 28411 28073
rect 28353 28064 28365 28067
rect 27120 28036 28365 28064
rect 27120 28024 27126 28036
rect 28353 28033 28365 28036
rect 28399 28033 28411 28067
rect 28534 28064 28540 28076
rect 28495 28036 28540 28064
rect 28353 28027 28411 28033
rect 28534 28024 28540 28036
rect 28592 28024 28598 28076
rect 29546 28064 29552 28076
rect 29507 28036 29552 28064
rect 29546 28024 29552 28036
rect 29604 28024 29610 28076
rect 18064 27996 18092 28024
rect 17328 27968 18092 27996
rect 18325 27999 18383 28005
rect 18325 27965 18337 27999
rect 18371 27965 18383 27999
rect 18325 27959 18383 27965
rect 25936 27999 25994 28005
rect 25936 27965 25948 27999
rect 25982 27996 25994 27999
rect 26050 27996 26056 28008
rect 25982 27968 26056 27996
rect 25982 27965 25994 27968
rect 25936 27959 25994 27965
rect 17954 27888 17960 27940
rect 18012 27928 18018 27940
rect 18340 27928 18368 27959
rect 26050 27956 26056 27968
rect 26108 27956 26114 28008
rect 26145 27999 26203 28005
rect 26145 27965 26157 27999
rect 26191 27965 26203 27999
rect 26145 27959 26203 27965
rect 18012 27900 18368 27928
rect 18012 27888 18018 27900
rect 24854 27888 24860 27940
rect 24912 27928 24918 27940
rect 26160 27928 26188 27959
rect 27706 27956 27712 28008
rect 27764 27996 27770 28008
rect 27893 27999 27951 28005
rect 27893 27996 27905 27999
rect 27764 27968 27905 27996
rect 27764 27956 27770 27968
rect 27893 27965 27905 27968
rect 27939 27965 27951 27999
rect 27893 27959 27951 27965
rect 27982 27956 27988 28008
rect 28040 27996 28046 28008
rect 28721 27999 28779 28005
rect 28721 27996 28733 27999
rect 28040 27968 28733 27996
rect 28040 27956 28046 27968
rect 28721 27965 28733 27968
rect 28767 27996 28779 27999
rect 29457 27999 29515 28005
rect 29457 27996 29469 27999
rect 28767 27968 29469 27996
rect 28767 27965 28779 27968
rect 28721 27959 28779 27965
rect 29457 27965 29469 27968
rect 29503 27965 29515 27999
rect 30208 27996 30236 28095
rect 30392 28064 30420 28095
rect 30558 28064 30564 28076
rect 30392 28036 30564 28064
rect 30558 28024 30564 28036
rect 30616 28024 30622 28076
rect 31294 28064 31300 28076
rect 31255 28036 31300 28064
rect 31294 28024 31300 28036
rect 31352 28024 31358 28076
rect 31573 28067 31631 28073
rect 31573 28033 31585 28067
rect 31619 28064 31631 28067
rect 32324 28064 32352 28172
rect 32582 28160 32588 28172
rect 32640 28160 32646 28212
rect 33318 28160 33324 28212
rect 33376 28200 33382 28212
rect 33781 28203 33839 28209
rect 33781 28200 33793 28203
rect 33376 28172 33793 28200
rect 33376 28160 33382 28172
rect 33781 28169 33793 28172
rect 33827 28169 33839 28203
rect 33781 28163 33839 28169
rect 36078 28160 36084 28212
rect 36136 28160 36142 28212
rect 36722 28200 36728 28212
rect 36683 28172 36728 28200
rect 36722 28160 36728 28172
rect 36780 28160 36786 28212
rect 32766 28132 32772 28144
rect 32416 28104 32772 28132
rect 32416 28073 32444 28104
rect 32766 28092 32772 28104
rect 32824 28132 32830 28144
rect 34054 28132 34060 28144
rect 32824 28104 34060 28132
rect 32824 28092 32830 28104
rect 34054 28092 34060 28104
rect 34112 28092 34118 28144
rect 36096 28132 36124 28160
rect 36096 28104 36400 28132
rect 32674 28073 32680 28076
rect 31619 28036 32352 28064
rect 32401 28067 32459 28073
rect 31619 28033 31631 28036
rect 31573 28027 31631 28033
rect 32401 28033 32413 28067
rect 32447 28033 32459 28067
rect 32401 28027 32459 28033
rect 32668 28027 32680 28073
rect 32732 28064 32738 28076
rect 34422 28064 34428 28076
rect 32732 28036 32768 28064
rect 34383 28036 34428 28064
rect 32674 28024 32680 28027
rect 32732 28024 32738 28036
rect 34422 28024 34428 28036
rect 34480 28024 34486 28076
rect 34609 28067 34667 28073
rect 34609 28033 34621 28067
rect 34655 28064 34667 28067
rect 35526 28064 35532 28076
rect 34655 28036 35532 28064
rect 34655 28033 34667 28036
rect 34609 28027 34667 28033
rect 35526 28024 35532 28036
rect 35584 28064 35590 28076
rect 36081 28067 36139 28073
rect 36081 28064 36093 28067
rect 35584 28036 36093 28064
rect 35584 28024 35590 28036
rect 36081 28033 36093 28036
rect 36127 28033 36139 28067
rect 36262 28064 36268 28076
rect 36223 28036 36268 28064
rect 36081 28027 36139 28033
rect 36262 28024 36268 28036
rect 36320 28024 36326 28076
rect 36372 28073 36400 28104
rect 36357 28067 36415 28073
rect 36357 28033 36369 28067
rect 36403 28033 36415 28067
rect 36357 28027 36415 28033
rect 36449 28067 36507 28073
rect 36449 28033 36461 28067
rect 36495 28064 36507 28067
rect 37458 28064 37464 28076
rect 36495 28036 36584 28064
rect 37419 28036 37464 28064
rect 36495 28033 36507 28036
rect 36449 28027 36507 28033
rect 30742 27996 30748 28008
rect 30208 27968 30748 27996
rect 29457 27959 29515 27965
rect 30742 27956 30748 27968
rect 30800 27956 30806 28008
rect 33594 27956 33600 28008
rect 33652 27996 33658 28008
rect 34241 27999 34299 28005
rect 34241 27996 34253 27999
rect 33652 27968 34253 27996
rect 33652 27956 33658 27968
rect 34241 27965 34253 27968
rect 34287 27965 34299 27999
rect 34241 27959 34299 27965
rect 30650 27928 30656 27940
rect 24912 27900 26188 27928
rect 27540 27900 30656 27928
rect 24912 27888 24918 27900
rect 16758 27820 16764 27872
rect 16816 27860 16822 27872
rect 17129 27863 17187 27869
rect 17129 27860 17141 27863
rect 16816 27832 17141 27860
rect 16816 27820 16822 27832
rect 17129 27829 17141 27832
rect 17175 27829 17187 27863
rect 17129 27823 17187 27829
rect 18322 27820 18328 27872
rect 18380 27860 18386 27872
rect 19429 27863 19487 27869
rect 19429 27860 19441 27863
rect 18380 27832 19441 27860
rect 18380 27820 18386 27832
rect 19429 27829 19441 27832
rect 19475 27829 19487 27863
rect 19429 27823 19487 27829
rect 20898 27820 20904 27872
rect 20956 27860 20962 27872
rect 20993 27863 21051 27869
rect 20993 27860 21005 27863
rect 20956 27832 21005 27860
rect 20956 27820 20962 27832
rect 20993 27829 21005 27832
rect 21039 27829 21051 27863
rect 25314 27860 25320 27872
rect 25275 27832 25320 27860
rect 20993 27823 21051 27829
rect 25314 27820 25320 27832
rect 25372 27820 25378 27872
rect 26602 27820 26608 27872
rect 26660 27860 26666 27872
rect 27540 27869 27568 27900
rect 30650 27888 30656 27900
rect 30708 27888 30714 27940
rect 31018 27928 31024 27940
rect 30979 27900 31024 27928
rect 31018 27888 31024 27900
rect 31076 27888 31082 27940
rect 27525 27863 27583 27869
rect 27525 27860 27537 27863
rect 26660 27832 27537 27860
rect 26660 27820 26666 27832
rect 27525 27829 27537 27832
rect 27571 27829 27583 27863
rect 27525 27823 27583 27829
rect 29549 27863 29607 27869
rect 29549 27829 29561 27863
rect 29595 27860 29607 27863
rect 29822 27860 29828 27872
rect 29595 27832 29828 27860
rect 29595 27829 29607 27832
rect 29549 27823 29607 27829
rect 29822 27820 29828 27832
rect 29880 27820 29886 27872
rect 30377 27863 30435 27869
rect 30377 27829 30389 27863
rect 30423 27860 30435 27863
rect 31036 27860 31064 27888
rect 30423 27832 31064 27860
rect 31481 27863 31539 27869
rect 30423 27829 30435 27832
rect 30377 27823 30435 27829
rect 31481 27829 31493 27863
rect 31527 27860 31539 27863
rect 31846 27860 31852 27872
rect 31527 27832 31852 27860
rect 31527 27829 31539 27832
rect 31481 27823 31539 27829
rect 31846 27820 31852 27832
rect 31904 27820 31910 27872
rect 36170 27820 36176 27872
rect 36228 27860 36234 27872
rect 36556 27860 36584 28036
rect 37458 28024 37464 28036
rect 37516 28024 37522 28076
rect 37369 27863 37427 27869
rect 37369 27860 37381 27863
rect 36228 27832 37381 27860
rect 36228 27820 36234 27832
rect 37369 27829 37381 27832
rect 37415 27829 37427 27863
rect 37369 27823 37427 27829
rect 43809 27863 43867 27869
rect 43809 27829 43821 27863
rect 43855 27860 43867 27863
rect 44174 27860 44180 27872
rect 43855 27832 44180 27860
rect 43855 27829 43867 27832
rect 43809 27823 43867 27829
rect 44174 27820 44180 27832
rect 44232 27820 44238 27872
rect 1104 27770 44896 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 44896 27770
rect 1104 27696 44896 27718
rect 16114 27616 16120 27668
rect 16172 27656 16178 27668
rect 16301 27659 16359 27665
rect 16301 27656 16313 27659
rect 16172 27628 16313 27656
rect 16172 27616 16178 27628
rect 16301 27625 16313 27628
rect 16347 27625 16359 27659
rect 16301 27619 16359 27625
rect 16574 27616 16580 27668
rect 16632 27656 16638 27668
rect 17221 27659 17279 27665
rect 17221 27656 17233 27659
rect 16632 27628 17233 27656
rect 16632 27616 16638 27628
rect 17221 27625 17233 27628
rect 17267 27625 17279 27659
rect 17221 27619 17279 27625
rect 17589 27659 17647 27665
rect 17589 27625 17601 27659
rect 17635 27656 17647 27659
rect 17954 27656 17960 27668
rect 17635 27628 17960 27656
rect 17635 27625 17647 27628
rect 17589 27619 17647 27625
rect 17954 27616 17960 27628
rect 18012 27616 18018 27668
rect 21085 27659 21143 27665
rect 21085 27625 21097 27659
rect 21131 27656 21143 27659
rect 22278 27656 22284 27668
rect 21131 27628 22284 27656
rect 21131 27625 21143 27628
rect 21085 27619 21143 27625
rect 22278 27616 22284 27628
rect 22336 27656 22342 27668
rect 22465 27659 22523 27665
rect 22465 27656 22477 27659
rect 22336 27628 22477 27656
rect 22336 27616 22342 27628
rect 22465 27625 22477 27628
rect 22511 27625 22523 27659
rect 22465 27619 22523 27625
rect 22649 27659 22707 27665
rect 22649 27625 22661 27659
rect 22695 27625 22707 27659
rect 22649 27619 22707 27625
rect 16666 27588 16672 27600
rect 16627 27560 16672 27588
rect 16666 27548 16672 27560
rect 16724 27548 16730 27600
rect 18233 27591 18291 27597
rect 18233 27557 18245 27591
rect 18279 27588 18291 27591
rect 18322 27588 18328 27600
rect 18279 27560 18328 27588
rect 18279 27557 18291 27560
rect 18233 27551 18291 27557
rect 18322 27548 18328 27560
rect 18380 27548 18386 27600
rect 20714 27588 20720 27600
rect 20675 27560 20720 27588
rect 20714 27548 20720 27560
rect 20772 27548 20778 27600
rect 21726 27548 21732 27600
rect 21784 27588 21790 27600
rect 21821 27591 21879 27597
rect 21821 27588 21833 27591
rect 21784 27560 21833 27588
rect 21784 27548 21790 27560
rect 21821 27557 21833 27560
rect 21867 27557 21879 27591
rect 22664 27588 22692 27619
rect 23014 27616 23020 27668
rect 23072 27656 23078 27668
rect 23385 27659 23443 27665
rect 23385 27656 23397 27659
rect 23072 27628 23397 27656
rect 23072 27616 23078 27628
rect 23385 27625 23397 27628
rect 23431 27625 23443 27659
rect 27890 27656 27896 27668
rect 23385 27619 23443 27625
rect 27632 27628 27896 27656
rect 22738 27588 22744 27600
rect 22651 27560 22744 27588
rect 21821 27551 21879 27557
rect 22738 27548 22744 27560
rect 22796 27588 22802 27600
rect 27065 27591 27123 27597
rect 22796 27560 23152 27588
rect 22796 27548 22802 27560
rect 17862 27480 17868 27532
rect 17920 27520 17926 27532
rect 18049 27523 18107 27529
rect 18049 27520 18061 27523
rect 17920 27492 18061 27520
rect 17920 27480 17926 27492
rect 18049 27489 18061 27492
rect 18095 27489 18107 27523
rect 18049 27483 18107 27489
rect 21177 27523 21235 27529
rect 21177 27489 21189 27523
rect 21223 27520 21235 27523
rect 21266 27520 21272 27532
rect 21223 27492 21272 27520
rect 21223 27489 21235 27492
rect 21177 27483 21235 27489
rect 21266 27480 21272 27492
rect 21324 27480 21330 27532
rect 23124 27464 23152 27560
rect 27065 27557 27077 27591
rect 27111 27588 27123 27591
rect 27632 27588 27660 27628
rect 27890 27616 27896 27628
rect 27948 27616 27954 27668
rect 30650 27616 30656 27668
rect 30708 27656 30714 27668
rect 31021 27659 31079 27665
rect 31021 27656 31033 27659
rect 30708 27628 31033 27656
rect 30708 27616 30714 27628
rect 31021 27625 31033 27628
rect 31067 27656 31079 27659
rect 31110 27656 31116 27668
rect 31067 27628 31116 27656
rect 31067 27625 31079 27628
rect 31021 27619 31079 27625
rect 31110 27616 31116 27628
rect 31168 27616 31174 27668
rect 32674 27656 32680 27668
rect 32635 27628 32680 27656
rect 32674 27616 32680 27628
rect 32732 27616 32738 27668
rect 36173 27659 36231 27665
rect 36173 27625 36185 27659
rect 36219 27656 36231 27659
rect 36262 27656 36268 27668
rect 36219 27628 36268 27656
rect 36219 27625 36231 27628
rect 36173 27619 36231 27625
rect 36262 27616 36268 27628
rect 36320 27616 36326 27668
rect 27111 27560 27660 27588
rect 27111 27557 27123 27560
rect 27065 27551 27123 27557
rect 30374 27548 30380 27600
rect 30432 27588 30438 27600
rect 31573 27591 31631 27597
rect 31573 27588 31585 27591
rect 30432 27560 31585 27588
rect 30432 27548 30438 27560
rect 31573 27557 31585 27560
rect 31619 27557 31631 27591
rect 31846 27588 31852 27600
rect 31807 27560 31852 27588
rect 31573 27551 31631 27557
rect 31846 27548 31852 27560
rect 31904 27548 31910 27600
rect 25682 27520 25688 27532
rect 25643 27492 25688 27520
rect 25682 27480 25688 27492
rect 25740 27480 25746 27532
rect 28994 27480 29000 27532
rect 29052 27520 29058 27532
rect 29549 27523 29607 27529
rect 29549 27520 29561 27523
rect 29052 27492 29561 27520
rect 29052 27480 29058 27492
rect 29549 27489 29561 27492
rect 29595 27489 29607 27523
rect 29822 27520 29828 27532
rect 29783 27492 29828 27520
rect 29549 27483 29607 27489
rect 29822 27480 29828 27492
rect 29880 27480 29886 27532
rect 42702 27520 42708 27532
rect 42663 27492 42708 27520
rect 42702 27480 42708 27492
rect 42760 27480 42766 27532
rect 43990 27520 43996 27532
rect 43951 27492 43996 27520
rect 43990 27480 43996 27492
rect 44048 27480 44054 27532
rect 44174 27520 44180 27532
rect 44135 27492 44180 27520
rect 44174 27480 44180 27492
rect 44232 27480 44238 27532
rect 16485 27455 16543 27461
rect 16485 27421 16497 27455
rect 16531 27421 16543 27455
rect 16485 27415 16543 27421
rect 16500 27384 16528 27415
rect 16666 27412 16672 27464
rect 16724 27452 16730 27464
rect 16761 27455 16819 27461
rect 16761 27452 16773 27455
rect 16724 27424 16773 27452
rect 16724 27412 16730 27424
rect 16761 27421 16773 27424
rect 16807 27421 16819 27455
rect 16761 27415 16819 27421
rect 16850 27412 16856 27464
rect 16908 27452 16914 27464
rect 17405 27455 17463 27461
rect 17405 27452 17417 27455
rect 16908 27424 17417 27452
rect 16908 27412 16914 27424
rect 17405 27421 17417 27424
rect 17451 27421 17463 27455
rect 17405 27415 17463 27421
rect 17589 27455 17647 27461
rect 17589 27421 17601 27455
rect 17635 27452 17647 27455
rect 17678 27452 17684 27464
rect 17635 27424 17684 27452
rect 17635 27421 17647 27424
rect 17589 27415 17647 27421
rect 17678 27412 17684 27424
rect 17736 27412 17742 27464
rect 17954 27412 17960 27464
rect 18012 27452 18018 27464
rect 18325 27455 18383 27461
rect 18325 27452 18337 27455
rect 18012 27424 18337 27452
rect 18012 27412 18018 27424
rect 18325 27421 18337 27424
rect 18371 27421 18383 27455
rect 20898 27452 20904 27464
rect 20859 27424 20904 27452
rect 18325 27415 18383 27421
rect 20898 27412 20904 27424
rect 20956 27412 20962 27464
rect 21634 27452 21640 27464
rect 21595 27424 21640 27452
rect 21634 27412 21640 27424
rect 21692 27412 21698 27464
rect 23106 27412 23112 27464
rect 23164 27452 23170 27464
rect 23290 27452 23296 27464
rect 23164 27424 23296 27452
rect 23164 27412 23170 27424
rect 23290 27412 23296 27424
rect 23348 27412 23354 27464
rect 23382 27412 23388 27464
rect 23440 27452 23446 27464
rect 23477 27455 23535 27461
rect 23477 27452 23489 27455
rect 23440 27424 23489 27452
rect 23440 27412 23446 27424
rect 23477 27421 23489 27424
rect 23523 27421 23535 27455
rect 23477 27415 23535 27421
rect 24578 27412 24584 27464
rect 24636 27452 24642 27464
rect 25041 27455 25099 27461
rect 25041 27452 25053 27455
rect 24636 27424 25053 27452
rect 24636 27412 24642 27424
rect 25041 27421 25053 27424
rect 25087 27421 25099 27455
rect 25700 27452 25728 27480
rect 27617 27455 27675 27461
rect 27617 27452 27629 27455
rect 25700 27424 27629 27452
rect 25041 27415 25099 27421
rect 27617 27421 27629 27424
rect 27663 27421 27675 27455
rect 27617 27415 27675 27421
rect 27884 27455 27942 27461
rect 27884 27421 27896 27455
rect 27930 27452 27942 27455
rect 28166 27452 28172 27464
rect 27930 27424 28172 27452
rect 27930 27421 27942 27424
rect 27884 27415 27942 27421
rect 28166 27412 28172 27424
rect 28224 27412 28230 27464
rect 30834 27452 30840 27464
rect 30795 27424 30840 27452
rect 30834 27412 30840 27424
rect 30892 27412 30898 27464
rect 31846 27452 31852 27464
rect 31807 27424 31852 27452
rect 31846 27412 31852 27424
rect 31904 27412 31910 27464
rect 32030 27452 32036 27464
rect 31991 27424 32036 27452
rect 32030 27412 32036 27424
rect 32088 27412 32094 27464
rect 32490 27452 32496 27464
rect 32451 27424 32496 27452
rect 32490 27412 32496 27424
rect 32548 27412 32554 27464
rect 34698 27452 34704 27464
rect 34659 27424 34704 27452
rect 34698 27412 34704 27424
rect 34756 27412 34762 27464
rect 34885 27455 34943 27461
rect 34885 27421 34897 27455
rect 34931 27421 34943 27455
rect 36078 27452 36084 27464
rect 36039 27424 36084 27452
rect 34885 27415 34943 27421
rect 20162 27384 20168 27396
rect 16500 27356 20168 27384
rect 20162 27344 20168 27356
rect 20220 27384 20226 27396
rect 20622 27384 20628 27396
rect 20220 27356 20628 27384
rect 20220 27344 20226 27356
rect 20622 27344 20628 27356
rect 20680 27344 20686 27396
rect 22833 27387 22891 27393
rect 22833 27353 22845 27387
rect 22879 27384 22891 27387
rect 23198 27384 23204 27396
rect 22879 27356 23204 27384
rect 22879 27353 22891 27356
rect 22833 27347 22891 27353
rect 23198 27344 23204 27356
rect 23256 27344 23262 27396
rect 25314 27344 25320 27396
rect 25372 27384 25378 27396
rect 25930 27387 25988 27393
rect 25930 27384 25942 27387
rect 25372 27356 25942 27384
rect 25372 27344 25378 27356
rect 25930 27353 25942 27356
rect 25976 27353 25988 27387
rect 25930 27347 25988 27353
rect 34606 27344 34612 27396
rect 34664 27384 34670 27396
rect 34900 27384 34928 27415
rect 36078 27412 36084 27424
rect 36136 27412 36142 27464
rect 36170 27412 36176 27464
rect 36228 27452 36234 27464
rect 36265 27455 36323 27461
rect 36265 27452 36277 27455
rect 36228 27424 36277 27452
rect 36228 27412 36234 27424
rect 36265 27421 36277 27424
rect 36311 27421 36323 27455
rect 36265 27415 36323 27421
rect 34664 27356 34928 27384
rect 34664 27344 34670 27356
rect 17586 27276 17592 27328
rect 17644 27316 17650 27328
rect 22646 27325 22652 27328
rect 18325 27319 18383 27325
rect 18325 27316 18337 27319
rect 17644 27288 18337 27316
rect 17644 27276 17650 27288
rect 18325 27285 18337 27288
rect 18371 27285 18383 27319
rect 22633 27319 22652 27325
rect 22633 27316 22645 27319
rect 22559 27288 22645 27316
rect 18325 27279 18383 27285
rect 22633 27285 22645 27288
rect 22704 27316 22710 27328
rect 23382 27316 23388 27328
rect 22704 27288 23388 27316
rect 22633 27279 22652 27285
rect 22646 27276 22652 27279
rect 22704 27276 22710 27288
rect 23382 27276 23388 27288
rect 23440 27276 23446 27328
rect 25130 27316 25136 27328
rect 25091 27288 25136 27316
rect 25130 27276 25136 27288
rect 25188 27276 25194 27328
rect 28902 27276 28908 27328
rect 28960 27316 28966 27328
rect 28997 27319 29055 27325
rect 28997 27316 29009 27319
rect 28960 27288 29009 27316
rect 28960 27276 28966 27288
rect 28997 27285 29009 27288
rect 29043 27285 29055 27319
rect 28997 27279 29055 27285
rect 31110 27276 31116 27328
rect 31168 27316 31174 27328
rect 33502 27316 33508 27328
rect 31168 27288 33508 27316
rect 31168 27276 31174 27288
rect 33502 27276 33508 27288
rect 33560 27276 33566 27328
rect 34422 27276 34428 27328
rect 34480 27316 34486 27328
rect 34793 27319 34851 27325
rect 34793 27316 34805 27319
rect 34480 27288 34805 27316
rect 34480 27276 34486 27288
rect 34793 27285 34805 27288
rect 34839 27285 34851 27319
rect 34793 27279 34851 27285
rect 1104 27226 44896 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 44896 27226
rect 1104 27152 44896 27174
rect 16117 27115 16175 27121
rect 16117 27081 16129 27115
rect 16163 27112 16175 27115
rect 16850 27112 16856 27124
rect 16163 27084 16856 27112
rect 16163 27081 16175 27084
rect 16117 27075 16175 27081
rect 16850 27072 16856 27084
rect 16908 27072 16914 27124
rect 28629 27115 28687 27121
rect 28629 27081 28641 27115
rect 28675 27112 28687 27115
rect 28718 27112 28724 27124
rect 28675 27084 28724 27112
rect 28675 27081 28687 27084
rect 28629 27075 28687 27081
rect 28718 27072 28724 27084
rect 28776 27072 28782 27124
rect 28994 27112 29000 27124
rect 28955 27084 29000 27112
rect 28994 27072 29000 27084
rect 29052 27072 29058 27124
rect 16666 27004 16672 27056
rect 16724 27044 16730 27056
rect 17267 27047 17325 27053
rect 17267 27044 17279 27047
rect 16724 27016 17279 27044
rect 16724 27004 16730 27016
rect 17267 27013 17279 27016
rect 17313 27013 17325 27047
rect 17402 27044 17408 27056
rect 17363 27016 17408 27044
rect 17267 27007 17325 27013
rect 17402 27004 17408 27016
rect 17460 27004 17466 27056
rect 17497 27047 17555 27053
rect 17497 27013 17509 27047
rect 17543 27044 17555 27047
rect 18325 27047 18383 27053
rect 18325 27044 18337 27047
rect 17543 27016 18337 27044
rect 17543 27013 17555 27016
rect 17497 27007 17555 27013
rect 18325 27013 18337 27016
rect 18371 27013 18383 27047
rect 18325 27007 18383 27013
rect 23109 27047 23167 27053
rect 23109 27013 23121 27047
rect 23155 27044 23167 27047
rect 24026 27044 24032 27056
rect 23155 27016 24032 27044
rect 23155 27013 23167 27016
rect 23109 27007 23167 27013
rect 24026 27004 24032 27016
rect 24084 27004 24090 27056
rect 27801 27047 27859 27053
rect 27801 27013 27813 27047
rect 27847 27044 27859 27047
rect 28534 27044 28540 27056
rect 27847 27016 28540 27044
rect 27847 27013 27859 27016
rect 27801 27007 27859 27013
rect 28534 27004 28540 27016
rect 28592 27004 28598 27056
rect 32950 27004 32956 27056
rect 33008 27044 33014 27056
rect 34146 27044 34152 27056
rect 33008 27016 34152 27044
rect 33008 27004 33014 27016
rect 34146 27004 34152 27016
rect 34204 27044 34210 27056
rect 34698 27044 34704 27056
rect 34204 27016 34704 27044
rect 34204 27004 34210 27016
rect 14274 26936 14280 26988
rect 14332 26976 14338 26988
rect 14737 26979 14795 26985
rect 14737 26976 14749 26979
rect 14332 26948 14749 26976
rect 14332 26936 14338 26948
rect 14737 26945 14749 26948
rect 14783 26945 14795 26979
rect 14737 26939 14795 26945
rect 15004 26979 15062 26985
rect 15004 26945 15016 26979
rect 15050 26976 15062 26979
rect 15470 26976 15476 26988
rect 15050 26948 15476 26976
rect 15050 26945 15062 26948
rect 15004 26939 15062 26945
rect 15470 26936 15476 26948
rect 15528 26936 15534 26988
rect 17586 26936 17592 26988
rect 17644 26976 17650 26988
rect 17644 26948 17689 26976
rect 17644 26936 17650 26948
rect 17862 26936 17868 26988
rect 17920 26976 17926 26988
rect 18417 26979 18475 26985
rect 18417 26976 18429 26979
rect 17920 26948 18429 26976
rect 17920 26936 17926 26948
rect 18417 26945 18429 26948
rect 18463 26945 18475 26979
rect 18417 26939 18475 26945
rect 22925 26979 22983 26985
rect 22925 26945 22937 26979
rect 22971 26945 22983 26979
rect 22925 26939 22983 26945
rect 23201 26979 23259 26985
rect 23201 26945 23213 26979
rect 23247 26976 23259 26979
rect 23290 26976 23296 26988
rect 23247 26948 23296 26976
rect 23247 26945 23259 26948
rect 23201 26939 23259 26945
rect 17129 26911 17187 26917
rect 17129 26877 17141 26911
rect 17175 26908 17187 26911
rect 17770 26908 17776 26920
rect 17175 26880 17776 26908
rect 17175 26877 17187 26880
rect 17129 26871 17187 26877
rect 17770 26868 17776 26880
rect 17828 26868 17834 26920
rect 22940 26908 22968 26939
rect 23290 26936 23296 26948
rect 23348 26936 23354 26988
rect 28721 26979 28779 26985
rect 28721 26945 28733 26979
rect 28767 26945 28779 26979
rect 28721 26939 28779 26945
rect 23474 26908 23480 26920
rect 22940 26880 23480 26908
rect 23474 26868 23480 26880
rect 23532 26868 23538 26920
rect 27985 26911 28043 26917
rect 27985 26877 27997 26911
rect 28031 26908 28043 26911
rect 28736 26908 28764 26939
rect 28810 26936 28816 26988
rect 28868 26976 28874 26988
rect 28868 26948 28913 26976
rect 28868 26936 28874 26948
rect 30834 26936 30840 26988
rect 30892 26976 30898 26988
rect 33594 26976 33600 26988
rect 30892 26948 33600 26976
rect 30892 26936 30898 26948
rect 33594 26936 33600 26948
rect 33652 26936 33658 26988
rect 33781 26979 33839 26985
rect 33781 26945 33793 26979
rect 33827 26976 33839 26979
rect 33962 26976 33968 26988
rect 33827 26948 33968 26976
rect 33827 26945 33839 26948
rect 33781 26939 33839 26945
rect 33962 26936 33968 26948
rect 34020 26976 34026 26988
rect 34238 26976 34244 26988
rect 34020 26948 34244 26976
rect 34020 26936 34026 26948
rect 34238 26936 34244 26948
rect 34296 26936 34302 26988
rect 34422 26976 34428 26988
rect 34383 26948 34428 26976
rect 34422 26936 34428 26948
rect 34480 26936 34486 26988
rect 34532 26985 34560 27016
rect 34698 27004 34704 27016
rect 34756 27004 34762 27056
rect 34885 27047 34943 27053
rect 34885 27013 34897 27047
rect 34931 27044 34943 27047
rect 36458 27047 36516 27053
rect 36458 27044 36470 27047
rect 34931 27016 36470 27044
rect 34931 27013 34943 27016
rect 34885 27007 34943 27013
rect 36458 27013 36470 27016
rect 36504 27013 36516 27047
rect 36458 27007 36516 27013
rect 34517 26979 34575 26985
rect 34517 26945 34529 26979
rect 34563 26945 34575 26979
rect 34517 26939 34575 26945
rect 34606 26936 34612 26988
rect 34664 26976 34670 26988
rect 34664 26948 34709 26976
rect 34664 26936 34670 26948
rect 28902 26908 28908 26920
rect 28031 26880 28580 26908
rect 28736 26880 28908 26908
rect 28031 26877 28043 26880
rect 27985 26871 28043 26877
rect 28552 26852 28580 26880
rect 28902 26868 28908 26880
rect 28960 26908 28966 26920
rect 31294 26908 31300 26920
rect 28960 26880 31300 26908
rect 28960 26868 28966 26880
rect 31294 26868 31300 26880
rect 31352 26868 31358 26920
rect 33321 26911 33379 26917
rect 33321 26877 33333 26911
rect 33367 26908 33379 26911
rect 34624 26908 34652 26936
rect 33367 26880 34652 26908
rect 36725 26911 36783 26917
rect 33367 26877 33379 26880
rect 33321 26871 33379 26877
rect 36725 26877 36737 26911
rect 36771 26908 36783 26911
rect 37182 26908 37188 26920
rect 36771 26880 37188 26908
rect 36771 26877 36783 26880
rect 36725 26871 36783 26877
rect 37182 26868 37188 26880
rect 37240 26868 37246 26920
rect 27522 26800 27528 26852
rect 27580 26840 27586 26852
rect 28445 26843 28503 26849
rect 28445 26840 28457 26843
rect 27580 26812 28457 26840
rect 27580 26800 27586 26812
rect 28445 26809 28457 26812
rect 28491 26809 28503 26843
rect 28445 26803 28503 26809
rect 28534 26800 28540 26852
rect 28592 26840 28598 26852
rect 29546 26840 29552 26852
rect 28592 26812 29552 26840
rect 28592 26800 28598 26812
rect 29546 26800 29552 26812
rect 29604 26800 29610 26852
rect 31846 26800 31852 26852
rect 31904 26840 31910 26852
rect 33413 26843 33471 26849
rect 33413 26840 33425 26843
rect 31904 26812 33425 26840
rect 31904 26800 31910 26812
rect 33413 26809 33425 26812
rect 33459 26809 33471 26843
rect 33413 26803 33471 26809
rect 16206 26732 16212 26784
rect 16264 26772 16270 26784
rect 17773 26775 17831 26781
rect 17773 26772 17785 26775
rect 16264 26744 17785 26772
rect 16264 26732 16270 26744
rect 17773 26741 17785 26744
rect 17819 26741 17831 26775
rect 23014 26772 23020 26784
rect 22975 26744 23020 26772
rect 17773 26735 17831 26741
rect 23014 26732 23020 26744
rect 23072 26732 23078 26784
rect 35342 26772 35348 26784
rect 35303 26744 35348 26772
rect 35342 26732 35348 26744
rect 35400 26732 35406 26784
rect 1104 26682 44896 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 44896 26682
rect 1104 26608 44896 26630
rect 15470 26568 15476 26580
rect 15431 26540 15476 26568
rect 15470 26528 15476 26540
rect 15528 26528 15534 26580
rect 16669 26571 16727 26577
rect 16669 26537 16681 26571
rect 16715 26568 16727 26571
rect 17402 26568 17408 26580
rect 16715 26540 17408 26568
rect 16715 26537 16727 26540
rect 16669 26531 16727 26537
rect 17402 26528 17408 26540
rect 17460 26528 17466 26580
rect 17589 26571 17647 26577
rect 17589 26537 17601 26571
rect 17635 26568 17647 26571
rect 17678 26568 17684 26580
rect 17635 26540 17684 26568
rect 17635 26537 17647 26540
rect 17589 26531 17647 26537
rect 17678 26528 17684 26540
rect 17736 26528 17742 26580
rect 28629 26571 28687 26577
rect 28629 26537 28641 26571
rect 28675 26568 28687 26571
rect 28810 26568 28816 26580
rect 28675 26540 28816 26568
rect 28675 26537 28687 26540
rect 28629 26531 28687 26537
rect 28810 26528 28816 26540
rect 28868 26528 28874 26580
rect 31846 26528 31852 26580
rect 31904 26568 31910 26580
rect 32217 26571 32275 26577
rect 32217 26568 32229 26571
rect 31904 26540 32229 26568
rect 31904 26528 31910 26540
rect 32217 26537 32229 26540
rect 32263 26537 32275 26571
rect 32217 26531 32275 26537
rect 32953 26571 33011 26577
rect 32953 26537 32965 26571
rect 32999 26568 33011 26571
rect 34606 26568 34612 26580
rect 32999 26540 34612 26568
rect 32999 26537 33011 26540
rect 32953 26531 33011 26537
rect 34606 26528 34612 26540
rect 34664 26528 34670 26580
rect 34698 26528 34704 26580
rect 34756 26568 34762 26580
rect 35069 26571 35127 26577
rect 35069 26568 35081 26571
rect 34756 26540 35081 26568
rect 34756 26528 34762 26540
rect 35069 26537 35081 26540
rect 35115 26537 35127 26571
rect 35069 26531 35127 26537
rect 16114 26500 16120 26512
rect 15396 26472 16120 26500
rect 15396 26373 15424 26472
rect 16114 26460 16120 26472
rect 16172 26500 16178 26512
rect 19978 26500 19984 26512
rect 16172 26472 19984 26500
rect 16172 26460 16178 26472
rect 19978 26460 19984 26472
rect 20036 26460 20042 26512
rect 22370 26500 22376 26512
rect 21376 26472 22376 26500
rect 17862 26392 17868 26444
rect 17920 26432 17926 26444
rect 18049 26435 18107 26441
rect 18049 26432 18061 26435
rect 17920 26404 18061 26432
rect 17920 26392 17926 26404
rect 18049 26401 18061 26404
rect 18095 26432 18107 26435
rect 19521 26435 19579 26441
rect 19521 26432 19533 26435
rect 18095 26404 19533 26432
rect 18095 26401 18107 26404
rect 18049 26395 18107 26401
rect 19521 26401 19533 26404
rect 19567 26401 19579 26435
rect 19521 26395 19579 26401
rect 15381 26367 15439 26373
rect 15381 26333 15393 26367
rect 15427 26333 15439 26367
rect 15381 26327 15439 26333
rect 15565 26367 15623 26373
rect 15565 26333 15577 26367
rect 15611 26364 15623 26367
rect 16206 26364 16212 26376
rect 15611 26336 16212 26364
rect 15611 26333 15623 26336
rect 15565 26327 15623 26333
rect 16206 26324 16212 26336
rect 16264 26324 16270 26376
rect 16758 26364 16764 26376
rect 16671 26336 16764 26364
rect 16758 26324 16764 26336
rect 16816 26364 16822 26376
rect 17405 26367 17463 26373
rect 17405 26364 17417 26367
rect 16816 26336 17417 26364
rect 16816 26324 16822 26336
rect 17405 26333 17417 26336
rect 17451 26333 17463 26367
rect 17405 26327 17463 26333
rect 17034 26256 17040 26308
rect 17092 26296 17098 26308
rect 17221 26299 17279 26305
rect 17221 26296 17233 26299
rect 17092 26268 17233 26296
rect 17092 26256 17098 26268
rect 17221 26265 17233 26268
rect 17267 26296 17279 26299
rect 17880 26296 17908 26392
rect 17954 26324 17960 26376
rect 18012 26364 18018 26376
rect 18233 26367 18291 26373
rect 18233 26364 18245 26367
rect 18012 26336 18245 26364
rect 18012 26324 18018 26336
rect 18233 26333 18245 26336
rect 18279 26333 18291 26367
rect 18233 26327 18291 26333
rect 18322 26324 18328 26376
rect 18380 26364 18386 26376
rect 19242 26364 19248 26376
rect 18380 26336 18425 26364
rect 19203 26336 19248 26364
rect 18380 26324 18386 26336
rect 19242 26324 19248 26336
rect 19300 26324 19306 26376
rect 21376 26373 21404 26472
rect 22370 26460 22376 26472
rect 22428 26500 22434 26512
rect 22428 26472 23336 26500
rect 22428 26460 22434 26472
rect 23308 26441 23336 26472
rect 23750 26460 23756 26512
rect 23808 26500 23814 26512
rect 23845 26503 23903 26509
rect 23845 26500 23857 26503
rect 23808 26472 23857 26500
rect 23808 26460 23814 26472
rect 23845 26469 23857 26472
rect 23891 26469 23903 26503
rect 26786 26500 26792 26512
rect 23845 26463 23903 26469
rect 24780 26472 26792 26500
rect 24780 26441 24808 26472
rect 26786 26460 26792 26472
rect 26844 26460 26850 26512
rect 31018 26500 31024 26512
rect 30979 26472 31024 26500
rect 31018 26460 31024 26472
rect 31076 26460 31082 26512
rect 32030 26500 32036 26512
rect 31726 26472 32036 26500
rect 23293 26435 23351 26441
rect 23293 26401 23305 26435
rect 23339 26432 23351 26435
rect 24765 26435 24823 26441
rect 24765 26432 24777 26435
rect 23339 26404 24777 26432
rect 23339 26401 23351 26404
rect 23293 26395 23351 26401
rect 24765 26401 24777 26404
rect 24811 26401 24823 26435
rect 24765 26395 24823 26401
rect 25041 26435 25099 26441
rect 25041 26401 25053 26435
rect 25087 26432 25099 26435
rect 31726 26432 31754 26472
rect 32030 26460 32036 26472
rect 32088 26500 32094 26512
rect 35342 26500 35348 26512
rect 32088 26472 35348 26500
rect 32088 26460 32094 26472
rect 35342 26460 35348 26472
rect 35400 26460 35406 26512
rect 35805 26503 35863 26509
rect 35805 26469 35817 26503
rect 35851 26469 35863 26503
rect 35805 26463 35863 26469
rect 25087 26404 25728 26432
rect 25087 26401 25099 26404
rect 25041 26395 25099 26401
rect 22094 26373 22100 26376
rect 20993 26367 21051 26373
rect 20993 26333 21005 26367
rect 21039 26364 21051 26367
rect 21361 26367 21419 26373
rect 21039 26336 21312 26364
rect 21039 26333 21051 26336
rect 20993 26327 21051 26333
rect 17267 26268 17908 26296
rect 21085 26299 21143 26305
rect 17267 26265 17279 26268
rect 17221 26259 17279 26265
rect 21085 26265 21097 26299
rect 21131 26265 21143 26299
rect 21085 26259 21143 26265
rect 21177 26299 21235 26305
rect 21177 26265 21189 26299
rect 21223 26265 21235 26299
rect 21284 26296 21312 26336
rect 21361 26333 21373 26367
rect 21407 26333 21419 26367
rect 22077 26367 22100 26373
rect 21361 26327 21419 26333
rect 21468 26361 22048 26364
rect 22077 26361 22089 26367
rect 21468 26336 22089 26361
rect 21468 26296 21496 26336
rect 22020 26333 22089 26336
rect 22077 26327 22100 26333
rect 22094 26324 22100 26327
rect 22152 26324 22158 26376
rect 22189 26367 22247 26373
rect 22189 26333 22201 26367
rect 22235 26333 22247 26367
rect 22189 26327 22247 26333
rect 21284 26268 21496 26296
rect 21821 26299 21879 26305
rect 21177 26259 21235 26265
rect 21821 26265 21833 26299
rect 21867 26296 21879 26299
rect 22204 26296 22232 26327
rect 22278 26324 22284 26376
rect 22336 26364 22342 26376
rect 22465 26367 22523 26373
rect 22336 26336 22381 26364
rect 22336 26324 22342 26336
rect 22465 26333 22477 26367
rect 22511 26364 22523 26367
rect 22922 26364 22928 26376
rect 22511 26336 22928 26364
rect 22511 26333 22523 26336
rect 22465 26327 22523 26333
rect 22922 26324 22928 26336
rect 22980 26324 22986 26376
rect 23382 26324 23388 26376
rect 23440 26364 23446 26376
rect 23477 26367 23535 26373
rect 23477 26364 23489 26367
rect 23440 26336 23489 26364
rect 23440 26324 23446 26336
rect 23477 26333 23489 26336
rect 23523 26333 23535 26367
rect 23477 26327 23535 26333
rect 24486 26324 24492 26376
rect 24544 26364 24550 26376
rect 24673 26367 24731 26373
rect 24673 26364 24685 26367
rect 24544 26336 24685 26364
rect 24544 26324 24550 26336
rect 24673 26333 24685 26336
rect 24719 26333 24731 26367
rect 25498 26364 25504 26376
rect 25459 26336 25504 26364
rect 24673 26327 24731 26333
rect 25498 26324 25504 26336
rect 25556 26324 25562 26376
rect 25700 26373 25728 26404
rect 31220 26404 31754 26432
rect 25685 26367 25743 26373
rect 25685 26333 25697 26367
rect 25731 26333 25743 26367
rect 25685 26327 25743 26333
rect 25869 26367 25927 26373
rect 25869 26333 25881 26367
rect 25915 26364 25927 26367
rect 26513 26367 26571 26373
rect 26513 26364 26525 26367
rect 25915 26336 26525 26364
rect 25915 26333 25927 26336
rect 25869 26327 25927 26333
rect 26513 26333 26525 26336
rect 26559 26333 26571 26367
rect 26513 26327 26571 26333
rect 27890 26324 27896 26376
rect 27948 26364 27954 26376
rect 31220 26373 31248 26404
rect 33318 26392 33324 26444
rect 33376 26432 33382 26444
rect 33689 26435 33747 26441
rect 33689 26432 33701 26435
rect 33376 26404 33701 26432
rect 33376 26392 33382 26404
rect 33689 26401 33701 26404
rect 33735 26432 33747 26435
rect 34701 26435 34759 26441
rect 34701 26432 34713 26435
rect 33735 26404 34713 26432
rect 33735 26401 33747 26404
rect 33689 26395 33747 26401
rect 34701 26401 34713 26404
rect 34747 26401 34759 26435
rect 34701 26395 34759 26401
rect 28537 26367 28595 26373
rect 28537 26364 28549 26367
rect 27948 26336 28549 26364
rect 27948 26324 27954 26336
rect 28537 26333 28549 26336
rect 28583 26333 28595 26367
rect 28537 26327 28595 26333
rect 31205 26367 31263 26373
rect 31205 26333 31217 26367
rect 31251 26333 31263 26367
rect 31205 26327 31263 26333
rect 31297 26367 31355 26373
rect 31297 26333 31309 26367
rect 31343 26364 31355 26367
rect 31478 26364 31484 26376
rect 31343 26336 31484 26364
rect 31343 26333 31355 26336
rect 31297 26327 31355 26333
rect 31478 26324 31484 26336
rect 31536 26324 31542 26376
rect 32122 26364 32128 26376
rect 32083 26336 32128 26364
rect 32122 26324 32128 26336
rect 32180 26324 32186 26376
rect 32309 26367 32367 26373
rect 32309 26333 32321 26367
rect 32355 26333 32367 26367
rect 33594 26364 33600 26376
rect 32309 26327 32367 26333
rect 32784 26336 33456 26364
rect 33555 26336 33600 26364
rect 23014 26296 23020 26308
rect 21867 26268 22094 26296
rect 22204 26268 23020 26296
rect 21867 26265 21879 26268
rect 21821 26259 21879 26265
rect 5166 26188 5172 26240
rect 5224 26228 5230 26240
rect 16574 26228 16580 26240
rect 5224 26200 16580 26228
rect 5224 26188 5230 26200
rect 16574 26188 16580 26200
rect 16632 26188 16638 26240
rect 18046 26228 18052 26240
rect 18007 26200 18052 26228
rect 18046 26188 18052 26200
rect 18104 26188 18110 26240
rect 20806 26228 20812 26240
rect 20767 26200 20812 26228
rect 20806 26188 20812 26200
rect 20864 26188 20870 26240
rect 20990 26188 20996 26240
rect 21048 26228 21054 26240
rect 21100 26228 21128 26259
rect 21048 26200 21128 26228
rect 21192 26228 21220 26259
rect 21266 26228 21272 26240
rect 21192 26200 21272 26228
rect 21048 26188 21054 26200
rect 21266 26188 21272 26200
rect 21324 26188 21330 26240
rect 22066 26228 22094 26268
rect 23014 26256 23020 26268
rect 23072 26256 23078 26308
rect 30282 26256 30288 26308
rect 30340 26296 30346 26308
rect 31021 26299 31079 26305
rect 31021 26296 31033 26299
rect 30340 26268 31033 26296
rect 30340 26256 30346 26268
rect 31021 26265 31033 26268
rect 31067 26265 31079 26299
rect 31021 26259 31079 26265
rect 31938 26256 31944 26308
rect 31996 26296 32002 26308
rect 32324 26296 32352 26327
rect 32784 26305 32812 26336
rect 32769 26299 32827 26305
rect 32769 26296 32781 26299
rect 31996 26268 32781 26296
rect 31996 26256 32002 26268
rect 32769 26265 32781 26268
rect 32815 26265 32827 26299
rect 33428 26296 33456 26336
rect 33594 26324 33600 26336
rect 33652 26324 33658 26376
rect 33778 26324 33784 26376
rect 33836 26364 33842 26376
rect 33873 26367 33931 26373
rect 33873 26364 33885 26367
rect 33836 26336 33885 26364
rect 33836 26324 33842 26336
rect 33873 26333 33885 26336
rect 33919 26333 33931 26367
rect 34514 26364 34520 26376
rect 33873 26327 33931 26333
rect 33964 26336 34520 26364
rect 33964 26296 33992 26336
rect 34514 26324 34520 26336
rect 34572 26364 34578 26376
rect 35820 26364 35848 26463
rect 41414 26392 41420 26444
rect 41472 26432 41478 26444
rect 42061 26435 42119 26441
rect 42061 26432 42073 26435
rect 41472 26404 42073 26432
rect 41472 26392 41478 26404
rect 42061 26401 42073 26404
rect 42107 26401 42119 26435
rect 42061 26395 42119 26401
rect 37182 26364 37188 26376
rect 34572 26336 35848 26364
rect 37143 26336 37188 26364
rect 34572 26324 34578 26336
rect 37182 26324 37188 26336
rect 37240 26324 37246 26376
rect 41598 26364 41604 26376
rect 41559 26336 41604 26364
rect 41598 26324 41604 26336
rect 41656 26324 41662 26376
rect 43898 26364 43904 26376
rect 43859 26336 43904 26364
rect 43898 26324 43904 26336
rect 43956 26324 43962 26376
rect 33428 26268 33992 26296
rect 32769 26259 32827 26265
rect 34238 26256 34244 26308
rect 34296 26296 34302 26308
rect 35069 26299 35127 26305
rect 35069 26296 35081 26299
rect 34296 26268 35081 26296
rect 34296 26256 34302 26268
rect 35069 26265 35081 26268
rect 35115 26265 35127 26299
rect 35069 26259 35127 26265
rect 35986 26256 35992 26308
rect 36044 26296 36050 26308
rect 36918 26299 36976 26305
rect 36918 26296 36930 26299
rect 36044 26268 36930 26296
rect 36044 26256 36050 26268
rect 36918 26265 36930 26268
rect 36964 26265 36976 26299
rect 41782 26296 41788 26308
rect 41743 26268 41788 26296
rect 36918 26259 36976 26265
rect 41782 26256 41788 26268
rect 41840 26256 41846 26308
rect 22186 26228 22192 26240
rect 22066 26200 22192 26228
rect 22186 26188 22192 26200
rect 22244 26188 22250 26240
rect 23385 26231 23443 26237
rect 23385 26197 23397 26231
rect 23431 26228 23443 26231
rect 23474 26228 23480 26240
rect 23431 26200 23480 26228
rect 23431 26197 23443 26200
rect 23385 26191 23443 26197
rect 23474 26188 23480 26200
rect 23532 26228 23538 26240
rect 24486 26228 24492 26240
rect 23532 26200 24492 26228
rect 23532 26188 23538 26200
rect 24486 26188 24492 26200
rect 24544 26188 24550 26240
rect 26326 26228 26332 26240
rect 26287 26200 26332 26228
rect 26326 26188 26332 26200
rect 26384 26188 26390 26240
rect 29822 26188 29828 26240
rect 29880 26228 29886 26240
rect 32950 26228 32956 26240
rect 33008 26237 33014 26240
rect 33008 26231 33037 26237
rect 29880 26200 32956 26228
rect 29880 26188 29886 26200
rect 32950 26188 32956 26200
rect 33025 26197 33037 26231
rect 33008 26191 33037 26197
rect 33137 26231 33195 26237
rect 33137 26197 33149 26231
rect 33183 26228 33195 26231
rect 33318 26228 33324 26240
rect 33183 26200 33324 26228
rect 33183 26197 33195 26200
rect 33137 26191 33195 26197
rect 33008 26188 33014 26191
rect 33318 26188 33324 26200
rect 33376 26188 33382 26240
rect 33870 26188 33876 26240
rect 33928 26228 33934 26240
rect 34057 26231 34115 26237
rect 34057 26228 34069 26231
rect 33928 26200 34069 26228
rect 33928 26188 33934 26200
rect 34057 26197 34069 26200
rect 34103 26197 34115 26231
rect 34057 26191 34115 26197
rect 35253 26231 35311 26237
rect 35253 26197 35265 26231
rect 35299 26228 35311 26231
rect 35710 26228 35716 26240
rect 35299 26200 35716 26228
rect 35299 26197 35311 26200
rect 35253 26191 35311 26197
rect 35710 26188 35716 26200
rect 35768 26188 35774 26240
rect 1104 26138 44896 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 44896 26138
rect 1104 26064 44896 26086
rect 16574 25984 16580 26036
rect 16632 26024 16638 26036
rect 16632 25996 28856 26024
rect 16632 25984 16638 25996
rect 3326 25956 3332 25968
rect 3287 25928 3332 25956
rect 3326 25916 3332 25928
rect 3384 25916 3390 25968
rect 15562 25916 15568 25968
rect 15620 25956 15626 25968
rect 24026 25956 24032 25968
rect 15620 25928 19748 25956
rect 15620 25916 15626 25928
rect 5166 25848 5172 25900
rect 5224 25888 5230 25900
rect 15838 25888 15844 25900
rect 5224 25860 5269 25888
rect 15799 25860 15844 25888
rect 5224 25848 5230 25860
rect 15838 25848 15844 25860
rect 15896 25848 15902 25900
rect 15933 25891 15991 25897
rect 15933 25857 15945 25891
rect 15979 25857 15991 25891
rect 15933 25851 15991 25857
rect 16117 25891 16175 25897
rect 16117 25857 16129 25891
rect 16163 25888 16175 25891
rect 16666 25888 16672 25900
rect 16163 25860 16672 25888
rect 16163 25857 16175 25860
rect 16117 25851 16175 25857
rect 3970 25780 3976 25832
rect 4028 25820 4034 25832
rect 4985 25823 5043 25829
rect 4985 25820 4997 25823
rect 4028 25792 4997 25820
rect 4028 25780 4034 25792
rect 4985 25789 4997 25792
rect 5031 25789 5043 25823
rect 4985 25783 5043 25789
rect 15948 25752 15976 25851
rect 16666 25848 16672 25860
rect 16724 25848 16730 25900
rect 17034 25888 17040 25900
rect 16995 25860 17040 25888
rect 17034 25848 17040 25860
rect 17092 25848 17098 25900
rect 17880 25897 17908 25928
rect 17865 25891 17923 25897
rect 17865 25857 17877 25891
rect 17911 25857 17923 25891
rect 17865 25851 17923 25857
rect 17954 25848 17960 25900
rect 18012 25848 18018 25900
rect 18138 25897 18144 25900
rect 18132 25851 18144 25897
rect 18196 25888 18202 25900
rect 19720 25897 19748 25928
rect 22066 25928 22324 25956
rect 23987 25928 24032 25956
rect 19978 25897 19984 25900
rect 19705 25891 19763 25897
rect 18196 25860 18232 25888
rect 18138 25848 18144 25851
rect 18196 25848 18202 25860
rect 19705 25857 19717 25891
rect 19751 25857 19763 25891
rect 19705 25851 19763 25857
rect 19972 25851 19984 25897
rect 20036 25888 20042 25900
rect 21913 25891 21971 25897
rect 20036 25860 20072 25888
rect 19978 25848 19984 25851
rect 20036 25848 20042 25860
rect 21913 25857 21925 25891
rect 21959 25888 21971 25891
rect 22066 25888 22094 25928
rect 22186 25897 22192 25900
rect 22180 25888 22192 25897
rect 21959 25860 22094 25888
rect 22147 25860 22192 25888
rect 21959 25857 21971 25860
rect 21913 25851 21971 25857
rect 22180 25851 22192 25860
rect 22186 25848 22192 25851
rect 22244 25848 22250 25900
rect 22296 25888 22324 25928
rect 24026 25916 24032 25928
rect 24084 25916 24090 25968
rect 24486 25956 24492 25968
rect 24447 25928 24492 25956
rect 24486 25916 24492 25928
rect 24544 25916 24550 25968
rect 25308 25959 25366 25965
rect 25308 25925 25320 25959
rect 25354 25956 25366 25959
rect 26326 25956 26332 25968
rect 25354 25928 26332 25956
rect 25354 25925 25366 25928
rect 25308 25919 25366 25925
rect 26326 25916 26332 25928
rect 26384 25916 26390 25968
rect 27062 25956 27068 25968
rect 26436 25928 27068 25956
rect 23658 25888 23664 25900
rect 22296 25860 23664 25888
rect 23658 25848 23664 25860
rect 23716 25888 23722 25900
rect 25041 25891 25099 25897
rect 25041 25888 25053 25891
rect 23716 25860 25053 25888
rect 23716 25848 23722 25860
rect 25041 25857 25053 25860
rect 25087 25857 25099 25891
rect 26436 25888 26464 25928
rect 27062 25916 27068 25928
rect 27120 25916 27126 25968
rect 27249 25959 27307 25965
rect 27249 25925 27261 25959
rect 27295 25956 27307 25959
rect 28828 25956 28856 25996
rect 30558 25984 30564 26036
rect 30616 26024 30622 26036
rect 31113 26027 31171 26033
rect 31113 26024 31125 26027
rect 30616 25996 31125 26024
rect 30616 25984 30622 25996
rect 31113 25993 31125 25996
rect 31159 25993 31171 26027
rect 31113 25987 31171 25993
rect 33505 26027 33563 26033
rect 33505 25993 33517 26027
rect 33551 26024 33563 26027
rect 33778 26024 33784 26036
rect 33551 25996 33784 26024
rect 33551 25993 33563 25996
rect 33505 25987 33563 25993
rect 33778 25984 33784 25996
rect 33836 25984 33842 26036
rect 34698 26024 34704 26036
rect 34659 25996 34704 26024
rect 34698 25984 34704 25996
rect 34756 25984 34762 26036
rect 35161 26027 35219 26033
rect 35161 25993 35173 26027
rect 35207 25993 35219 26027
rect 35986 26024 35992 26036
rect 35947 25996 35992 26024
rect 35161 25987 35219 25993
rect 32030 25956 32036 25968
rect 27295 25928 28764 25956
rect 28828 25928 32036 25956
rect 27295 25925 27307 25928
rect 27249 25919 27307 25925
rect 28736 25897 28764 25928
rect 32030 25916 32036 25928
rect 32088 25916 32094 25968
rect 32122 25916 32128 25968
rect 32180 25956 32186 25968
rect 33413 25959 33471 25965
rect 33413 25956 33425 25959
rect 32180 25928 33425 25956
rect 32180 25916 32186 25928
rect 33413 25925 33425 25928
rect 33459 25956 33471 25959
rect 33594 25956 33600 25968
rect 33459 25928 33600 25956
rect 33459 25925 33471 25928
rect 33413 25919 33471 25925
rect 33594 25916 33600 25928
rect 33652 25916 33658 25968
rect 34333 25959 34391 25965
rect 34333 25925 34345 25959
rect 34379 25956 34391 25959
rect 34606 25956 34612 25968
rect 34379 25928 34612 25956
rect 34379 25925 34391 25928
rect 34333 25919 34391 25925
rect 34606 25916 34612 25928
rect 34664 25956 34670 25968
rect 35176 25956 35204 25987
rect 35986 25984 35992 25996
rect 36044 25984 36050 26036
rect 41598 25984 41604 26036
rect 41656 26024 41662 26036
rect 42429 26027 42487 26033
rect 42429 26024 42441 26027
rect 41656 25996 42441 26024
rect 41656 25984 41662 25996
rect 42429 25993 42441 25996
rect 42475 25993 42487 26027
rect 42429 25987 42487 25993
rect 34664 25928 35204 25956
rect 34664 25916 34670 25928
rect 25041 25851 25099 25857
rect 25148 25860 26464 25888
rect 26973 25891 27031 25897
rect 16758 25820 16764 25832
rect 16719 25792 16764 25820
rect 16758 25780 16764 25792
rect 16816 25780 16822 25832
rect 16945 25823 17003 25829
rect 16945 25789 16957 25823
rect 16991 25820 17003 25823
rect 17972 25820 18000 25848
rect 23937 25823 23995 25829
rect 23937 25820 23949 25823
rect 16991 25792 18000 25820
rect 23124 25792 23949 25820
rect 16991 25789 17003 25792
rect 16945 25783 17003 25789
rect 16853 25755 16911 25761
rect 16853 25752 16865 25755
rect 15948 25724 16865 25752
rect 16853 25721 16865 25724
rect 16899 25721 16911 25755
rect 19242 25752 19248 25764
rect 19203 25724 19248 25752
rect 16853 25715 16911 25721
rect 19242 25712 19248 25724
rect 19300 25712 19306 25764
rect 15838 25684 15844 25696
rect 15799 25656 15844 25684
rect 15838 25644 15844 25656
rect 15896 25644 15902 25696
rect 20990 25644 20996 25696
rect 21048 25684 21054 25696
rect 21085 25687 21143 25693
rect 21085 25684 21097 25687
rect 21048 25656 21097 25684
rect 21048 25644 21054 25656
rect 21085 25653 21097 25656
rect 21131 25684 21143 25687
rect 23124 25684 23152 25792
rect 23937 25789 23949 25792
rect 23983 25820 23995 25823
rect 25148 25820 25176 25860
rect 26973 25857 26985 25891
rect 27019 25857 27031 25891
rect 26973 25851 27031 25857
rect 28537 25891 28595 25897
rect 28537 25857 28549 25891
rect 28583 25857 28595 25891
rect 28537 25851 28595 25857
rect 28721 25891 28779 25897
rect 28721 25857 28733 25891
rect 28767 25857 28779 25891
rect 28721 25851 28779 25857
rect 28813 25891 28871 25897
rect 28813 25857 28825 25891
rect 28859 25857 28871 25891
rect 28813 25851 28871 25857
rect 23983 25792 25176 25820
rect 23983 25789 23995 25792
rect 23937 25783 23995 25789
rect 23290 25752 23296 25764
rect 23251 25724 23296 25752
rect 23290 25712 23296 25724
rect 23348 25752 23354 25764
rect 24489 25755 24547 25761
rect 24489 25752 24501 25755
rect 23348 25724 24501 25752
rect 23348 25712 23354 25724
rect 24489 25721 24501 25724
rect 24535 25721 24547 25755
rect 24489 25715 24547 25721
rect 26421 25755 26479 25761
rect 26421 25721 26433 25755
rect 26467 25752 26479 25755
rect 26510 25752 26516 25764
rect 26467 25724 26516 25752
rect 26467 25721 26479 25724
rect 26421 25715 26479 25721
rect 26510 25712 26516 25724
rect 26568 25752 26574 25764
rect 26988 25752 27016 25851
rect 27249 25823 27307 25829
rect 27249 25789 27261 25823
rect 27295 25820 27307 25823
rect 27614 25820 27620 25832
rect 27295 25792 27620 25820
rect 27295 25789 27307 25792
rect 27249 25783 27307 25789
rect 27614 25780 27620 25792
rect 27672 25780 27678 25832
rect 26568 25724 27016 25752
rect 26568 25712 26574 25724
rect 21131 25656 23152 25684
rect 21131 25653 21143 25656
rect 21085 25647 21143 25653
rect 23566 25644 23572 25696
rect 23624 25684 23630 25696
rect 23753 25687 23811 25693
rect 23753 25684 23765 25687
rect 23624 25656 23765 25684
rect 23624 25644 23630 25656
rect 23753 25653 23765 25656
rect 23799 25653 23811 25687
rect 23753 25647 23811 25653
rect 26142 25644 26148 25696
rect 26200 25684 26206 25696
rect 27065 25687 27123 25693
rect 27065 25684 27077 25687
rect 26200 25656 27077 25684
rect 26200 25644 26206 25656
rect 27065 25653 27077 25656
rect 27111 25653 27123 25687
rect 28552 25684 28580 25851
rect 28626 25712 28632 25764
rect 28684 25752 28690 25764
rect 28828 25752 28856 25851
rect 28902 25848 28908 25900
rect 28960 25888 28966 25900
rect 30653 25891 30711 25897
rect 28960 25860 29005 25888
rect 28960 25848 28966 25860
rect 30653 25857 30665 25891
rect 30699 25888 30711 25891
rect 31018 25888 31024 25900
rect 30699 25860 31024 25888
rect 30699 25857 30711 25860
rect 30653 25851 30711 25857
rect 31018 25848 31024 25860
rect 31076 25848 31082 25900
rect 31172 25891 31230 25897
rect 31172 25857 31184 25891
rect 31218 25888 31230 25891
rect 31754 25888 31760 25900
rect 31218 25860 31760 25888
rect 31218 25857 31230 25860
rect 31172 25851 31230 25857
rect 31754 25848 31760 25860
rect 31812 25848 31818 25900
rect 32309 25891 32367 25897
rect 32309 25857 32321 25891
rect 32355 25888 32367 25891
rect 33318 25888 33324 25900
rect 32355 25860 33180 25888
rect 33279 25860 33324 25888
rect 32355 25857 32367 25860
rect 32309 25851 32367 25857
rect 30466 25780 30472 25832
rect 30524 25820 30530 25832
rect 32324 25820 32352 25851
rect 30524 25792 32352 25820
rect 32493 25823 32551 25829
rect 30524 25780 30530 25792
rect 32493 25789 32505 25823
rect 32539 25820 32551 25823
rect 33042 25820 33048 25832
rect 32539 25792 33048 25820
rect 32539 25789 32551 25792
rect 32493 25783 32551 25789
rect 33042 25780 33048 25792
rect 33100 25780 33106 25832
rect 33152 25820 33180 25860
rect 33318 25848 33324 25860
rect 33376 25848 33382 25900
rect 33781 25891 33839 25897
rect 33781 25857 33793 25891
rect 33827 25888 33839 25891
rect 33962 25888 33968 25900
rect 33827 25860 33968 25888
rect 33827 25857 33839 25860
rect 33781 25851 33839 25857
rect 33962 25848 33968 25860
rect 34020 25848 34026 25900
rect 34146 25848 34152 25900
rect 34204 25888 34210 25900
rect 34241 25891 34299 25897
rect 34241 25888 34253 25891
rect 34204 25860 34253 25888
rect 34204 25848 34210 25860
rect 34241 25857 34253 25860
rect 34287 25857 34299 25891
rect 34514 25888 34520 25900
rect 34475 25860 34520 25888
rect 34241 25851 34299 25857
rect 34514 25848 34520 25860
rect 34572 25848 34578 25900
rect 35342 25888 35348 25900
rect 35303 25860 35348 25888
rect 35342 25848 35348 25860
rect 35400 25848 35406 25900
rect 35710 25848 35716 25900
rect 35768 25888 35774 25900
rect 35805 25891 35863 25897
rect 35805 25888 35817 25891
rect 35768 25860 35817 25888
rect 35768 25848 35774 25860
rect 35805 25857 35817 25860
rect 35851 25857 35863 25891
rect 37366 25888 37372 25900
rect 35805 25851 35863 25857
rect 35912 25860 37372 25888
rect 35912 25820 35940 25860
rect 37366 25848 37372 25860
rect 37424 25888 37430 25900
rect 37533 25891 37591 25897
rect 37533 25888 37545 25891
rect 37424 25860 37545 25888
rect 37424 25848 37430 25860
rect 37533 25857 37545 25860
rect 37579 25857 37591 25891
rect 37533 25851 37591 25857
rect 38930 25848 38936 25900
rect 38988 25888 38994 25900
rect 39209 25891 39267 25897
rect 39209 25888 39221 25891
rect 38988 25860 39221 25888
rect 38988 25848 38994 25860
rect 39209 25857 39221 25860
rect 39255 25857 39267 25891
rect 39209 25851 39267 25857
rect 41690 25848 41696 25900
rect 41748 25888 41754 25900
rect 42613 25891 42671 25897
rect 42613 25888 42625 25891
rect 41748 25860 42625 25888
rect 41748 25848 41754 25860
rect 42613 25857 42625 25860
rect 42659 25857 42671 25891
rect 42613 25851 42671 25857
rect 33152 25792 35940 25820
rect 37182 25780 37188 25832
rect 37240 25820 37246 25832
rect 37277 25823 37335 25829
rect 37277 25820 37289 25823
rect 37240 25792 37289 25820
rect 37240 25780 37246 25792
rect 37277 25789 37289 25792
rect 37323 25789 37335 25823
rect 37277 25783 37335 25789
rect 28684 25724 28856 25752
rect 28684 25712 28690 25724
rect 32030 25712 32036 25764
rect 32088 25752 32094 25764
rect 32088 25724 32260 25752
rect 32088 25712 32094 25724
rect 28994 25684 29000 25696
rect 28552 25656 29000 25684
rect 27065 25647 27123 25653
rect 28994 25644 29000 25656
rect 29052 25644 29058 25696
rect 29181 25687 29239 25693
rect 29181 25653 29193 25687
rect 29227 25684 29239 25687
rect 30745 25687 30803 25693
rect 30745 25684 30757 25687
rect 29227 25656 30757 25684
rect 29227 25653 29239 25656
rect 29181 25647 29239 25653
rect 30745 25653 30757 25656
rect 30791 25653 30803 25687
rect 30745 25647 30803 25653
rect 30834 25644 30840 25696
rect 30892 25684 30898 25696
rect 31297 25687 31355 25693
rect 31297 25684 31309 25687
rect 30892 25656 31309 25684
rect 30892 25644 30898 25656
rect 31297 25653 31309 25656
rect 31343 25653 31355 25687
rect 31297 25647 31355 25653
rect 31386 25644 31392 25696
rect 31444 25684 31450 25696
rect 32125 25687 32183 25693
rect 32125 25684 32137 25687
rect 31444 25656 32137 25684
rect 31444 25644 31450 25656
rect 32125 25653 32137 25656
rect 32171 25653 32183 25687
rect 32232 25684 32260 25724
rect 39393 25687 39451 25693
rect 39393 25684 39405 25687
rect 32232 25656 39405 25684
rect 32125 25647 32183 25653
rect 39393 25653 39405 25656
rect 39439 25653 39451 25687
rect 39393 25647 39451 25653
rect 43809 25687 43867 25693
rect 43809 25653 43821 25687
rect 43855 25684 43867 25687
rect 44174 25684 44180 25696
rect 43855 25656 44180 25684
rect 43855 25653 43867 25656
rect 43809 25647 43867 25653
rect 44174 25644 44180 25656
rect 44232 25644 44238 25696
rect 1104 25594 44896 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 44896 25594
rect 1104 25520 44896 25542
rect 3881 25483 3939 25489
rect 3881 25449 3893 25483
rect 3927 25480 3939 25483
rect 3970 25480 3976 25492
rect 3927 25452 3976 25480
rect 3927 25449 3939 25452
rect 3881 25443 3939 25449
rect 3970 25440 3976 25452
rect 4028 25440 4034 25492
rect 16758 25440 16764 25492
rect 16816 25480 16822 25492
rect 16945 25483 17003 25489
rect 16945 25480 16957 25483
rect 16816 25452 16957 25480
rect 16816 25440 16822 25452
rect 16945 25449 16957 25452
rect 16991 25449 17003 25483
rect 17954 25480 17960 25492
rect 17915 25452 17960 25480
rect 16945 25443 17003 25449
rect 17954 25440 17960 25452
rect 18012 25440 18018 25492
rect 18138 25440 18144 25492
rect 18196 25480 18202 25492
rect 18233 25483 18291 25489
rect 18233 25480 18245 25483
rect 18196 25452 18245 25480
rect 18196 25440 18202 25452
rect 18233 25449 18245 25452
rect 18279 25449 18291 25483
rect 21266 25480 21272 25492
rect 21227 25452 21272 25480
rect 18233 25443 18291 25449
rect 21266 25440 21272 25452
rect 21324 25440 21330 25492
rect 22094 25480 22100 25492
rect 22055 25452 22100 25480
rect 22094 25440 22100 25452
rect 22152 25440 22158 25492
rect 24486 25440 24492 25492
rect 24544 25480 24550 25492
rect 26283 25483 26341 25489
rect 26283 25480 26295 25483
rect 24544 25452 26295 25480
rect 24544 25440 24550 25452
rect 26283 25449 26295 25452
rect 26329 25449 26341 25483
rect 27614 25480 27620 25492
rect 27575 25452 27620 25480
rect 26283 25443 26341 25449
rect 27614 25440 27620 25452
rect 27672 25440 27678 25492
rect 28626 25440 28632 25492
rect 28684 25480 28690 25492
rect 29641 25483 29699 25489
rect 29641 25480 29653 25483
rect 28684 25452 29653 25480
rect 28684 25440 28690 25452
rect 29641 25449 29653 25452
rect 29687 25449 29699 25483
rect 29641 25443 29699 25449
rect 29733 25483 29791 25489
rect 29733 25449 29745 25483
rect 29779 25480 29791 25483
rect 30374 25480 30380 25492
rect 29779 25452 30380 25480
rect 29779 25449 29791 25452
rect 29733 25443 29791 25449
rect 30374 25440 30380 25452
rect 30432 25440 30438 25492
rect 30466 25440 30472 25492
rect 30524 25480 30530 25492
rect 30561 25483 30619 25489
rect 30561 25480 30573 25483
rect 30524 25452 30573 25480
rect 30524 25440 30530 25452
rect 30561 25449 30573 25452
rect 30607 25449 30619 25483
rect 38930 25480 38936 25492
rect 38891 25452 38936 25480
rect 30561 25443 30619 25449
rect 38930 25440 38936 25452
rect 38988 25440 38994 25492
rect 23014 25412 23020 25424
rect 21100 25384 23020 25412
rect 15562 25344 15568 25356
rect 15523 25316 15568 25344
rect 15562 25304 15568 25316
rect 15620 25304 15626 25356
rect 18046 25304 18052 25356
rect 18104 25344 18110 25356
rect 18141 25347 18199 25353
rect 18141 25344 18153 25347
rect 18104 25316 18153 25344
rect 18104 25304 18110 25316
rect 18141 25313 18153 25316
rect 18187 25313 18199 25347
rect 18141 25307 18199 25313
rect 19981 25347 20039 25353
rect 19981 25313 19993 25347
rect 20027 25344 20039 25347
rect 20438 25344 20444 25356
rect 20027 25316 20444 25344
rect 20027 25313 20039 25316
rect 19981 25307 20039 25313
rect 20438 25304 20444 25316
rect 20496 25304 20502 25356
rect 21100 25353 21128 25384
rect 23014 25372 23020 25384
rect 23072 25372 23078 25424
rect 25225 25415 25283 25421
rect 25225 25381 25237 25415
rect 25271 25412 25283 25415
rect 30745 25415 30803 25421
rect 25271 25384 29776 25412
rect 25271 25381 25283 25384
rect 25225 25375 25283 25381
rect 21085 25347 21143 25353
rect 21085 25313 21097 25347
rect 21131 25313 21143 25347
rect 23566 25344 23572 25356
rect 21085 25307 21143 25313
rect 22296 25316 23572 25344
rect 3970 25276 3976 25288
rect 3931 25248 3976 25276
rect 3970 25236 3976 25248
rect 4028 25236 4034 25288
rect 15838 25285 15844 25288
rect 15832 25276 15844 25285
rect 15799 25248 15844 25276
rect 15832 25239 15844 25248
rect 15838 25236 15844 25239
rect 15896 25236 15902 25288
rect 17862 25276 17868 25288
rect 17823 25248 17868 25276
rect 17862 25236 17868 25248
rect 17920 25236 17926 25288
rect 18233 25279 18291 25285
rect 18233 25245 18245 25279
rect 18279 25276 18291 25279
rect 18598 25276 18604 25288
rect 18279 25248 18604 25276
rect 18279 25245 18291 25248
rect 18233 25239 18291 25245
rect 18598 25236 18604 25248
rect 18656 25276 18662 25288
rect 19058 25276 19064 25288
rect 18656 25248 19064 25276
rect 18656 25236 18662 25248
rect 19058 25236 19064 25248
rect 19116 25236 19122 25288
rect 20165 25279 20223 25285
rect 20165 25245 20177 25279
rect 20211 25276 20223 25279
rect 20806 25276 20812 25288
rect 20211 25248 20812 25276
rect 20211 25245 20223 25248
rect 20165 25239 20223 25245
rect 20806 25236 20812 25248
rect 20864 25236 20870 25288
rect 20990 25276 20996 25288
rect 20951 25248 20996 25276
rect 20990 25236 20996 25248
rect 21048 25236 21054 25288
rect 22296 25285 22324 25316
rect 23566 25304 23572 25316
rect 23624 25304 23630 25356
rect 24765 25347 24823 25353
rect 24765 25313 24777 25347
rect 24811 25344 24823 25347
rect 25406 25344 25412 25356
rect 24811 25316 25412 25344
rect 24811 25313 24823 25316
rect 24765 25307 24823 25313
rect 25406 25304 25412 25316
rect 25464 25344 25470 25356
rect 26510 25344 26516 25356
rect 25464 25316 26372 25344
rect 26471 25316 26516 25344
rect 25464 25304 25470 25316
rect 22097 25279 22155 25285
rect 22097 25245 22109 25279
rect 22143 25245 22155 25279
rect 22097 25239 22155 25245
rect 22281 25279 22339 25285
rect 22281 25245 22293 25279
rect 22327 25245 22339 25279
rect 22281 25239 22339 25245
rect 23293 25279 23351 25285
rect 23293 25245 23305 25279
rect 23339 25276 23351 25279
rect 23382 25276 23388 25288
rect 23339 25248 23388 25276
rect 23339 25245 23351 25248
rect 23293 25239 23351 25245
rect 22112 25208 22140 25239
rect 23382 25236 23388 25248
rect 23440 25236 23446 25288
rect 24673 25279 24731 25285
rect 24673 25245 24685 25279
rect 24719 25245 24731 25279
rect 24946 25276 24952 25288
rect 24907 25248 24952 25276
rect 24673 25239 24731 25245
rect 22370 25208 22376 25220
rect 22112 25180 22376 25208
rect 22370 25168 22376 25180
rect 22428 25168 22434 25220
rect 24688 25208 24716 25239
rect 24946 25236 24952 25248
rect 25004 25236 25010 25288
rect 25041 25279 25099 25285
rect 25041 25245 25053 25279
rect 25087 25276 25099 25279
rect 26142 25276 26148 25288
rect 25087 25248 26148 25276
rect 25087 25245 25099 25248
rect 25041 25239 25099 25245
rect 26142 25236 26148 25248
rect 26200 25236 26206 25288
rect 26344 25276 26372 25316
rect 26510 25304 26516 25316
rect 26568 25304 26574 25356
rect 26896 25316 27200 25344
rect 26896 25276 26924 25316
rect 27172 25285 27200 25316
rect 27890 25304 27896 25356
rect 27948 25344 27954 25356
rect 28721 25347 28779 25353
rect 28721 25344 28733 25347
rect 27948 25316 28733 25344
rect 27948 25304 27954 25316
rect 28721 25313 28733 25316
rect 28767 25313 28779 25347
rect 28721 25307 28779 25313
rect 28902 25304 28908 25356
rect 28960 25344 28966 25356
rect 29748 25353 29776 25384
rect 30745 25381 30757 25415
rect 30791 25412 30803 25415
rect 32769 25415 32827 25421
rect 30791 25384 31340 25412
rect 30791 25381 30803 25384
rect 30745 25375 30803 25381
rect 31312 25353 31340 25384
rect 32769 25381 32781 25415
rect 32815 25381 32827 25415
rect 32769 25375 32827 25381
rect 29733 25347 29791 25353
rect 28960 25316 29592 25344
rect 28960 25304 28966 25316
rect 26344 25248 26924 25276
rect 26973 25279 27031 25285
rect 26973 25245 26985 25279
rect 27019 25245 27031 25279
rect 26973 25239 27031 25245
rect 27157 25279 27215 25285
rect 27157 25245 27169 25279
rect 27203 25245 27215 25279
rect 27430 25276 27436 25288
rect 27391 25248 27436 25276
rect 27157 25239 27215 25245
rect 25130 25208 25136 25220
rect 24688 25180 25136 25208
rect 25130 25168 25136 25180
rect 25188 25168 25194 25220
rect 20346 25140 20352 25152
rect 20307 25112 20352 25140
rect 20346 25100 20352 25112
rect 20404 25100 20410 25152
rect 23106 25100 23112 25152
rect 23164 25140 23170 25152
rect 26988 25140 27016 25239
rect 27430 25236 27436 25248
rect 27488 25236 27494 25288
rect 27522 25236 27528 25288
rect 27580 25276 27586 25288
rect 28445 25279 28503 25285
rect 28445 25276 28457 25279
rect 27580 25248 28457 25276
rect 27580 25236 27586 25248
rect 28445 25245 28457 25248
rect 28491 25245 28503 25279
rect 28626 25276 28632 25288
rect 28587 25248 28632 25276
rect 28445 25239 28503 25245
rect 28626 25236 28632 25248
rect 28684 25236 28690 25288
rect 28813 25279 28871 25285
rect 28813 25245 28825 25279
rect 28859 25276 28871 25279
rect 28859 25248 28948 25276
rect 28859 25245 28871 25248
rect 28813 25239 28871 25245
rect 27448 25208 27476 25236
rect 28920 25208 28948 25248
rect 28994 25236 29000 25288
rect 29052 25276 29058 25288
rect 29564 25285 29592 25316
rect 29733 25313 29745 25347
rect 29779 25313 29791 25347
rect 29733 25307 29791 25313
rect 31297 25347 31355 25353
rect 31297 25313 31309 25347
rect 31343 25313 31355 25347
rect 31297 25307 31355 25313
rect 31389 25347 31447 25353
rect 31389 25313 31401 25347
rect 31435 25344 31447 25347
rect 32122 25344 32128 25356
rect 31435 25316 32128 25344
rect 31435 25313 31447 25316
rect 31389 25307 31447 25313
rect 32122 25304 32128 25316
rect 32180 25344 32186 25356
rect 32784 25344 32812 25375
rect 32180 25316 32812 25344
rect 41325 25347 41383 25353
rect 32180 25304 32186 25316
rect 41325 25313 41337 25347
rect 41371 25344 41383 25347
rect 41414 25344 41420 25356
rect 41371 25316 41420 25344
rect 41371 25313 41383 25316
rect 41325 25307 41383 25313
rect 41414 25304 41420 25316
rect 41472 25304 41478 25356
rect 41877 25347 41935 25353
rect 41877 25313 41889 25347
rect 41923 25344 41935 25347
rect 43898 25344 43904 25356
rect 41923 25316 43904 25344
rect 41923 25313 41935 25316
rect 41877 25307 41935 25313
rect 43898 25304 43904 25316
rect 43956 25304 43962 25356
rect 44082 25344 44088 25356
rect 44043 25316 44088 25344
rect 44082 25304 44088 25316
rect 44140 25304 44146 25356
rect 29549 25279 29607 25285
rect 29052 25248 29097 25276
rect 29052 25236 29058 25248
rect 29549 25245 29561 25279
rect 29595 25245 29607 25279
rect 31018 25276 31024 25288
rect 29549 25239 29607 25245
rect 29932 25248 31024 25276
rect 29932 25217 29960 25248
rect 31018 25236 31024 25248
rect 31076 25236 31082 25288
rect 31478 25276 31484 25288
rect 31439 25248 31484 25276
rect 31478 25236 31484 25248
rect 31536 25236 31542 25288
rect 31573 25279 31631 25285
rect 31573 25245 31585 25279
rect 31619 25245 31631 25279
rect 31573 25239 31631 25245
rect 29917 25211 29975 25217
rect 29917 25208 29929 25211
rect 27448 25180 29929 25208
rect 29917 25177 29929 25180
rect 29963 25177 29975 25211
rect 29917 25171 29975 25177
rect 30377 25211 30435 25217
rect 30377 25177 30389 25211
rect 30423 25208 30435 25211
rect 30742 25208 30748 25220
rect 30423 25180 30748 25208
rect 30423 25177 30435 25180
rect 30377 25171 30435 25177
rect 30742 25168 30748 25180
rect 30800 25168 30806 25220
rect 31202 25168 31208 25220
rect 31260 25208 31266 25220
rect 31588 25208 31616 25239
rect 33870 25236 33876 25288
rect 33928 25285 33934 25288
rect 33928 25276 33940 25285
rect 33928 25248 33973 25276
rect 33928 25239 33940 25248
rect 33928 25236 33934 25239
rect 34054 25236 34060 25288
rect 34112 25276 34118 25288
rect 34149 25279 34207 25285
rect 34149 25276 34161 25279
rect 34112 25248 34161 25276
rect 34112 25236 34118 25248
rect 34149 25245 34161 25248
rect 34195 25245 34207 25279
rect 34149 25239 34207 25245
rect 39117 25279 39175 25285
rect 39117 25245 39129 25279
rect 39163 25245 39175 25279
rect 39298 25276 39304 25288
rect 39259 25248 39304 25276
rect 39117 25239 39175 25245
rect 31260 25180 31616 25208
rect 39132 25208 39160 25239
rect 39298 25236 39304 25248
rect 39356 25236 39362 25288
rect 42334 25276 42340 25288
rect 42295 25248 42340 25276
rect 42334 25236 42340 25248
rect 42392 25236 42398 25288
rect 40862 25208 40868 25220
rect 39132 25180 40868 25208
rect 31260 25168 31266 25180
rect 40862 25168 40868 25180
rect 40920 25168 40926 25220
rect 41693 25211 41751 25217
rect 41693 25177 41705 25211
rect 41739 25177 41751 25211
rect 42518 25208 42524 25220
rect 42479 25180 42524 25208
rect 41693 25171 41751 25177
rect 23164 25112 27016 25140
rect 28261 25143 28319 25149
rect 23164 25100 23170 25112
rect 28261 25109 28273 25143
rect 28307 25140 28319 25143
rect 30190 25140 30196 25152
rect 28307 25112 30196 25140
rect 28307 25109 28319 25112
rect 28261 25103 28319 25109
rect 30190 25100 30196 25112
rect 30248 25100 30254 25152
rect 30558 25100 30564 25152
rect 30616 25149 30622 25152
rect 30616 25143 30635 25149
rect 30623 25109 30635 25143
rect 30616 25103 30635 25109
rect 30616 25100 30622 25103
rect 31754 25100 31760 25152
rect 31812 25140 31818 25152
rect 41708 25140 41736 25171
rect 42518 25168 42524 25180
rect 42576 25168 42582 25220
rect 43990 25140 43996 25152
rect 31812 25112 31857 25140
rect 41708 25112 43996 25140
rect 31812 25100 31818 25112
rect 43990 25100 43996 25112
rect 44048 25100 44054 25152
rect 1104 25050 44896 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 44896 25050
rect 1104 24976 44896 24998
rect 19978 24896 19984 24948
rect 20036 24936 20042 24948
rect 20165 24939 20223 24945
rect 20165 24936 20177 24939
rect 20036 24908 20177 24936
rect 20036 24896 20042 24908
rect 20165 24905 20177 24908
rect 20211 24905 20223 24939
rect 20165 24899 20223 24905
rect 30374 24896 30380 24948
rect 30432 24936 30438 24948
rect 30432 24908 32444 24936
rect 30432 24896 30438 24908
rect 28626 24828 28632 24880
rect 28684 24868 28690 24880
rect 28684 24840 31248 24868
rect 28684 24828 28690 24840
rect 20346 24800 20352 24812
rect 20307 24772 20352 24800
rect 20346 24760 20352 24772
rect 20404 24760 20410 24812
rect 22370 24760 22376 24812
rect 22428 24800 22434 24812
rect 23017 24803 23075 24809
rect 23017 24800 23029 24803
rect 22428 24772 23029 24800
rect 22428 24760 22434 24772
rect 23017 24769 23029 24772
rect 23063 24769 23075 24803
rect 23290 24800 23296 24812
rect 23251 24772 23296 24800
rect 23017 24763 23075 24769
rect 23290 24760 23296 24772
rect 23348 24800 23354 24812
rect 24673 24803 24731 24809
rect 24673 24800 24685 24803
rect 23348 24772 24685 24800
rect 23348 24760 23354 24772
rect 24673 24769 24685 24772
rect 24719 24769 24731 24803
rect 24673 24763 24731 24769
rect 24765 24803 24823 24809
rect 24765 24769 24777 24803
rect 24811 24800 24823 24803
rect 24946 24800 24952 24812
rect 24811 24772 24952 24800
rect 24811 24769 24823 24772
rect 24765 24763 24823 24769
rect 24946 24760 24952 24772
rect 25004 24760 25010 24812
rect 25317 24803 25375 24809
rect 25317 24800 25329 24803
rect 25056 24772 25329 24800
rect 22278 24692 22284 24744
rect 22336 24732 22342 24744
rect 22833 24735 22891 24741
rect 22833 24732 22845 24735
rect 22336 24704 22845 24732
rect 22336 24692 22342 24704
rect 22833 24701 22845 24704
rect 22879 24701 22891 24735
rect 22833 24695 22891 24701
rect 23109 24735 23167 24741
rect 23109 24701 23121 24735
rect 23155 24701 23167 24735
rect 23109 24695 23167 24701
rect 23201 24735 23259 24741
rect 23201 24701 23213 24735
rect 23247 24732 23259 24735
rect 24026 24732 24032 24744
rect 23247 24704 24032 24732
rect 23247 24701 23259 24704
rect 23201 24695 23259 24701
rect 23124 24664 23152 24695
rect 24026 24692 24032 24704
rect 24084 24692 24090 24744
rect 24486 24664 24492 24676
rect 23124 24636 24492 24664
rect 24486 24624 24492 24636
rect 24544 24624 24550 24676
rect 23198 24556 23204 24608
rect 23256 24596 23262 24608
rect 25056 24596 25084 24772
rect 25317 24769 25329 24772
rect 25363 24769 25375 24803
rect 25590 24800 25596 24812
rect 25551 24772 25596 24800
rect 25317 24763 25375 24769
rect 25590 24760 25596 24772
rect 25648 24760 25654 24812
rect 25685 24803 25743 24809
rect 25685 24769 25697 24803
rect 25731 24800 25743 24803
rect 26142 24800 26148 24812
rect 25731 24772 26148 24800
rect 25731 24769 25743 24772
rect 25685 24763 25743 24769
rect 26142 24760 26148 24772
rect 26200 24760 26206 24812
rect 29086 24800 29092 24812
rect 29047 24772 29092 24800
rect 29086 24760 29092 24772
rect 29144 24760 29150 24812
rect 29546 24800 29552 24812
rect 29459 24772 29552 24800
rect 29546 24760 29552 24772
rect 29604 24800 29610 24812
rect 30837 24803 30895 24809
rect 30837 24800 30849 24803
rect 29604 24772 30849 24800
rect 29604 24760 29610 24772
rect 30837 24769 30849 24772
rect 30883 24769 30895 24803
rect 31018 24800 31024 24812
rect 30979 24772 31024 24800
rect 30837 24763 30895 24769
rect 31018 24760 31024 24772
rect 31076 24760 31082 24812
rect 31220 24809 31248 24840
rect 31754 24828 31760 24880
rect 31812 24868 31818 24880
rect 32125 24871 32183 24877
rect 32125 24868 32137 24871
rect 31812 24840 32137 24868
rect 31812 24828 31818 24840
rect 32125 24837 32137 24840
rect 32171 24837 32183 24871
rect 32125 24831 32183 24837
rect 31205 24803 31263 24809
rect 31205 24769 31217 24803
rect 31251 24769 31263 24803
rect 31205 24763 31263 24769
rect 31294 24760 31300 24812
rect 31352 24800 31358 24812
rect 31389 24803 31447 24809
rect 31389 24800 31401 24803
rect 31352 24772 31401 24800
rect 31352 24760 31358 24772
rect 31389 24769 31401 24772
rect 31435 24769 31447 24803
rect 32306 24800 32312 24812
rect 32267 24772 32312 24800
rect 31389 24763 31447 24769
rect 32306 24760 32312 24772
rect 32364 24760 32370 24812
rect 32416 24809 32444 24908
rect 39298 24896 39304 24948
rect 39356 24936 39362 24948
rect 39669 24939 39727 24945
rect 39669 24936 39681 24939
rect 39356 24908 39681 24936
rect 39356 24896 39362 24908
rect 39669 24905 39681 24908
rect 39715 24905 39727 24939
rect 39669 24899 39727 24905
rect 37182 24828 37188 24880
rect 37240 24868 37246 24880
rect 37240 24840 38792 24868
rect 37240 24828 37246 24840
rect 38304 24809 38332 24840
rect 38562 24809 38568 24812
rect 32401 24803 32459 24809
rect 32401 24769 32413 24803
rect 32447 24769 32459 24803
rect 32401 24763 32459 24769
rect 32861 24803 32919 24809
rect 32861 24769 32873 24803
rect 32907 24769 32919 24803
rect 32861 24763 32919 24769
rect 38289 24803 38347 24809
rect 38289 24769 38301 24803
rect 38335 24769 38347 24803
rect 38289 24763 38347 24769
rect 38556 24763 38568 24809
rect 38620 24800 38626 24812
rect 38764 24800 38792 24840
rect 38620 24772 38656 24800
rect 38764 24772 39988 24800
rect 25406 24732 25412 24744
rect 25367 24704 25412 24732
rect 25406 24692 25412 24704
rect 25464 24692 25470 24744
rect 28994 24692 29000 24744
rect 29052 24732 29058 24744
rect 29825 24735 29883 24741
rect 29825 24732 29837 24735
rect 29052 24704 29837 24732
rect 29052 24692 29058 24704
rect 29825 24701 29837 24704
rect 29871 24701 29883 24735
rect 31110 24732 31116 24744
rect 31071 24704 31116 24732
rect 29825 24695 29883 24701
rect 25866 24664 25872 24676
rect 25827 24636 25872 24664
rect 25866 24624 25872 24636
rect 25924 24624 25930 24676
rect 27614 24624 27620 24676
rect 27672 24664 27678 24676
rect 27801 24667 27859 24673
rect 27801 24664 27813 24667
rect 27672 24636 27813 24664
rect 27672 24624 27678 24636
rect 27801 24633 27813 24636
rect 27847 24664 27859 24667
rect 29454 24664 29460 24676
rect 27847 24636 29460 24664
rect 27847 24633 27859 24636
rect 27801 24627 27859 24633
rect 29454 24624 29460 24636
rect 29512 24624 29518 24676
rect 23256 24568 25084 24596
rect 29840 24596 29868 24695
rect 31110 24692 31116 24704
rect 31168 24692 31174 24744
rect 32876 24732 32904 24763
rect 38562 24760 38568 24763
rect 38620 24760 38626 24772
rect 39960 24744 39988 24772
rect 40034 24760 40040 24812
rect 40092 24800 40098 24812
rect 40385 24803 40443 24809
rect 40385 24800 40397 24803
rect 40092 24772 40397 24800
rect 40092 24760 40098 24772
rect 40385 24769 40397 24772
rect 40431 24769 40443 24803
rect 42426 24800 42432 24812
rect 42387 24772 42432 24800
rect 40385 24763 40443 24769
rect 42426 24760 42432 24772
rect 42484 24760 42490 24812
rect 43254 24800 43260 24812
rect 43215 24772 43260 24800
rect 43254 24760 43260 24772
rect 43312 24760 43318 24812
rect 43714 24760 43720 24812
rect 43772 24800 43778 24812
rect 43901 24803 43959 24809
rect 43901 24800 43913 24803
rect 43772 24772 43913 24800
rect 43772 24760 43778 24772
rect 43901 24769 43913 24772
rect 43947 24769 43959 24803
rect 43901 24763 43959 24769
rect 43990 24760 43996 24812
rect 44048 24800 44054 24812
rect 44048 24772 44093 24800
rect 44048 24760 44054 24772
rect 31312 24704 32904 24732
rect 30558 24624 30564 24676
rect 30616 24664 30622 24676
rect 31312 24664 31340 24704
rect 39942 24692 39948 24744
rect 40000 24732 40006 24744
rect 40129 24735 40187 24741
rect 40129 24732 40141 24735
rect 40000 24704 40141 24732
rect 40000 24692 40006 24704
rect 40129 24701 40141 24704
rect 40175 24701 40187 24735
rect 40129 24695 40187 24701
rect 41782 24692 41788 24744
rect 41840 24732 41846 24744
rect 42521 24735 42579 24741
rect 42521 24732 42533 24735
rect 41840 24704 42533 24732
rect 41840 24692 41846 24704
rect 42521 24701 42533 24704
rect 42567 24701 42579 24735
rect 42521 24695 42579 24701
rect 32398 24664 32404 24676
rect 30616 24636 31340 24664
rect 31404 24636 32404 24664
rect 30616 24624 30622 24636
rect 30282 24596 30288 24608
rect 29840 24568 30288 24596
rect 23256 24556 23262 24568
rect 30282 24556 30288 24568
rect 30340 24596 30346 24608
rect 31404 24596 31432 24636
rect 32398 24624 32404 24636
rect 32456 24624 32462 24676
rect 30340 24568 31432 24596
rect 31573 24599 31631 24605
rect 30340 24556 30346 24568
rect 31573 24565 31585 24599
rect 31619 24596 31631 24599
rect 32030 24596 32036 24608
rect 31619 24568 32036 24596
rect 31619 24565 31631 24568
rect 31573 24559 31631 24565
rect 32030 24556 32036 24568
rect 32088 24556 32094 24608
rect 32125 24599 32183 24605
rect 32125 24565 32137 24599
rect 32171 24596 32183 24599
rect 32306 24596 32312 24608
rect 32171 24568 32312 24596
rect 32171 24565 32183 24568
rect 32125 24559 32183 24565
rect 32306 24556 32312 24568
rect 32364 24556 32370 24608
rect 32950 24596 32956 24608
rect 32911 24568 32956 24596
rect 32950 24556 32956 24568
rect 33008 24556 33014 24608
rect 41506 24596 41512 24608
rect 41467 24568 41512 24596
rect 41506 24556 41512 24568
rect 41564 24556 41570 24608
rect 43346 24596 43352 24608
rect 43307 24568 43352 24596
rect 43346 24556 43352 24568
rect 43404 24556 43410 24608
rect 1104 24506 44896 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 44896 24506
rect 1104 24432 44896 24454
rect 26142 24392 26148 24404
rect 26103 24364 26148 24392
rect 26142 24352 26148 24364
rect 26200 24352 26206 24404
rect 26973 24395 27031 24401
rect 26973 24361 26985 24395
rect 27019 24392 27031 24395
rect 27430 24392 27436 24404
rect 27019 24364 27436 24392
rect 27019 24361 27031 24364
rect 26973 24355 27031 24361
rect 27430 24352 27436 24364
rect 27488 24352 27494 24404
rect 27890 24392 27896 24404
rect 27851 24364 27896 24392
rect 27890 24352 27896 24364
rect 27948 24352 27954 24404
rect 28813 24395 28871 24401
rect 28813 24361 28825 24395
rect 28859 24392 28871 24395
rect 29546 24392 29552 24404
rect 28859 24364 29552 24392
rect 28859 24361 28871 24364
rect 28813 24355 28871 24361
rect 29546 24352 29552 24364
rect 29604 24352 29610 24404
rect 30193 24395 30251 24401
rect 30193 24361 30205 24395
rect 30239 24392 30251 24395
rect 30558 24392 30564 24404
rect 30239 24364 30564 24392
rect 30239 24361 30251 24364
rect 30193 24355 30251 24361
rect 30558 24352 30564 24364
rect 30616 24352 30622 24404
rect 31297 24395 31355 24401
rect 31297 24361 31309 24395
rect 31343 24392 31355 24395
rect 31386 24392 31392 24404
rect 31343 24364 31392 24392
rect 31343 24361 31355 24364
rect 31297 24355 31355 24361
rect 31386 24352 31392 24364
rect 31444 24352 31450 24404
rect 31754 24352 31760 24404
rect 31812 24392 31818 24404
rect 32033 24395 32091 24401
rect 32033 24392 32045 24395
rect 31812 24364 32045 24392
rect 31812 24352 31818 24364
rect 32033 24361 32045 24364
rect 32079 24361 32091 24395
rect 32033 24355 32091 24361
rect 32125 24395 32183 24401
rect 32125 24361 32137 24395
rect 32171 24392 32183 24395
rect 32950 24392 32956 24404
rect 32171 24364 32956 24392
rect 32171 24361 32183 24364
rect 32125 24355 32183 24361
rect 26712 24296 28580 24324
rect 15562 24256 15568 24268
rect 15523 24228 15568 24256
rect 15562 24216 15568 24228
rect 15620 24216 15626 24268
rect 17957 24259 18015 24265
rect 17957 24225 17969 24259
rect 18003 24256 18015 24259
rect 18138 24256 18144 24268
rect 18003 24228 18144 24256
rect 18003 24225 18015 24228
rect 17957 24219 18015 24225
rect 18138 24216 18144 24228
rect 18196 24216 18202 24268
rect 18233 24259 18291 24265
rect 18233 24225 18245 24259
rect 18279 24225 18291 24259
rect 20162 24256 20168 24268
rect 20123 24228 20168 24256
rect 18233 24219 18291 24225
rect 16390 24148 16396 24200
rect 16448 24188 16454 24200
rect 18248 24188 18276 24219
rect 20162 24216 20168 24228
rect 20220 24216 20226 24268
rect 20438 24256 20444 24268
rect 20399 24228 20444 24256
rect 20438 24216 20444 24228
rect 20496 24216 20502 24268
rect 25225 24259 25283 24265
rect 25225 24225 25237 24259
rect 25271 24256 25283 24259
rect 25590 24256 25596 24268
rect 25271 24228 25596 24256
rect 25271 24225 25283 24228
rect 25225 24219 25283 24225
rect 25590 24216 25596 24228
rect 25648 24216 25654 24268
rect 16448 24160 18276 24188
rect 18325 24191 18383 24197
rect 16448 24148 16454 24160
rect 18325 24157 18337 24191
rect 18371 24188 18383 24191
rect 18598 24188 18604 24200
rect 18371 24160 18604 24188
rect 18371 24157 18383 24160
rect 18325 24151 18383 24157
rect 18598 24148 18604 24160
rect 18656 24148 18662 24200
rect 20180 24188 20208 24216
rect 22370 24188 22376 24200
rect 20180 24160 22376 24188
rect 22370 24148 22376 24160
rect 22428 24148 22434 24200
rect 23750 24188 23756 24200
rect 23711 24160 23756 24188
rect 23750 24148 23756 24160
rect 23808 24148 23814 24200
rect 24949 24191 25007 24197
rect 24949 24157 24961 24191
rect 24995 24157 25007 24191
rect 24949 24151 25007 24157
rect 15832 24123 15890 24129
rect 15832 24089 15844 24123
rect 15878 24120 15890 24123
rect 17954 24120 17960 24132
rect 15878 24092 17960 24120
rect 15878 24089 15890 24092
rect 15832 24083 15890 24089
rect 17954 24080 17960 24092
rect 18012 24080 18018 24132
rect 23474 24120 23480 24132
rect 23435 24092 23480 24120
rect 23474 24080 23480 24092
rect 23532 24080 23538 24132
rect 23661 24123 23719 24129
rect 23661 24089 23673 24123
rect 23707 24120 23719 24123
rect 24026 24120 24032 24132
rect 23707 24092 24032 24120
rect 23707 24089 23719 24092
rect 23661 24083 23719 24089
rect 24026 24080 24032 24092
rect 24084 24120 24090 24132
rect 24964 24120 24992 24151
rect 25406 24148 25412 24200
rect 25464 24188 25470 24200
rect 26053 24191 26111 24197
rect 26053 24188 26065 24191
rect 25464 24160 26065 24188
rect 25464 24148 25470 24160
rect 26053 24157 26065 24160
rect 26099 24157 26111 24191
rect 26234 24188 26240 24200
rect 26195 24160 26240 24188
rect 26053 24151 26111 24157
rect 24084 24092 24992 24120
rect 26068 24120 26096 24151
rect 26234 24148 26240 24160
rect 26292 24148 26298 24200
rect 26712 24197 26740 24296
rect 28552 24256 28580 24296
rect 28718 24284 28724 24336
rect 28776 24324 28782 24336
rect 30285 24327 30343 24333
rect 30285 24324 30297 24327
rect 28776 24296 30297 24324
rect 28776 24284 28782 24296
rect 30285 24293 30297 24296
rect 30331 24324 30343 24327
rect 30374 24324 30380 24336
rect 30331 24296 30380 24324
rect 30331 24293 30343 24296
rect 30285 24287 30343 24293
rect 30374 24284 30380 24296
rect 30432 24284 30438 24336
rect 26896 24228 27752 24256
rect 28552 24228 29960 24256
rect 26697 24191 26755 24197
rect 26697 24157 26709 24191
rect 26743 24157 26755 24191
rect 26697 24151 26755 24157
rect 26896 24120 26924 24228
rect 27724 24200 27752 24228
rect 27062 24148 27068 24200
rect 27120 24188 27126 24200
rect 27433 24191 27491 24197
rect 27433 24188 27445 24191
rect 27120 24160 27445 24188
rect 27120 24148 27126 24160
rect 27433 24157 27445 24160
rect 27479 24157 27491 24191
rect 27433 24151 27491 24157
rect 27522 24148 27528 24200
rect 27580 24188 27586 24200
rect 27580 24160 27625 24188
rect 27580 24148 27586 24160
rect 27706 24148 27712 24200
rect 27764 24188 27770 24200
rect 28629 24191 28687 24197
rect 27764 24160 27857 24188
rect 27764 24148 27770 24160
rect 28629 24157 28641 24191
rect 28675 24188 28687 24191
rect 28718 24188 28724 24200
rect 28675 24160 28724 24188
rect 28675 24157 28687 24160
rect 28629 24151 28687 24157
rect 28718 24148 28724 24160
rect 28776 24148 28782 24200
rect 29932 24188 29960 24228
rect 30190 24216 30196 24268
rect 30248 24256 30254 24268
rect 32030 24256 32036 24268
rect 30248 24228 31156 24256
rect 31991 24228 32036 24256
rect 30248 24216 30254 24228
rect 30377 24191 30435 24197
rect 30377 24188 30389 24191
rect 29932 24160 30389 24188
rect 30377 24157 30389 24160
rect 30423 24188 30435 24191
rect 30650 24188 30656 24200
rect 30423 24160 30656 24188
rect 30423 24157 30435 24160
rect 30377 24151 30435 24157
rect 30650 24148 30656 24160
rect 30708 24148 30714 24200
rect 31128 24197 31156 24228
rect 32030 24216 32036 24228
rect 32088 24216 32094 24268
rect 31021 24191 31079 24197
rect 31021 24157 31033 24191
rect 31067 24157 31079 24191
rect 31021 24151 31079 24157
rect 31113 24191 31171 24197
rect 31113 24157 31125 24191
rect 31159 24157 31171 24191
rect 31113 24151 31171 24157
rect 31389 24191 31447 24197
rect 31389 24157 31401 24191
rect 31435 24188 31447 24191
rect 32140 24188 32168 24355
rect 32950 24352 32956 24364
rect 33008 24352 33014 24404
rect 41049 24395 41107 24401
rect 41049 24361 41061 24395
rect 41095 24392 41107 24395
rect 41690 24392 41696 24404
rect 41095 24364 41696 24392
rect 41095 24361 41107 24364
rect 41049 24355 41107 24361
rect 41690 24352 41696 24364
rect 41748 24352 41754 24404
rect 41785 24395 41843 24401
rect 41785 24361 41797 24395
rect 41831 24392 41843 24395
rect 42518 24392 42524 24404
rect 41831 24364 42524 24392
rect 41831 24361 41843 24364
rect 41785 24355 41843 24361
rect 42518 24352 42524 24364
rect 42576 24352 42582 24404
rect 40681 24259 40739 24265
rect 40681 24225 40693 24259
rect 40727 24256 40739 24259
rect 41506 24256 41512 24268
rect 40727 24228 41512 24256
rect 40727 24225 40739 24228
rect 40681 24219 40739 24225
rect 41506 24216 41512 24228
rect 41564 24216 41570 24268
rect 42702 24256 42708 24268
rect 42663 24228 42708 24256
rect 42702 24216 42708 24228
rect 42760 24216 42766 24268
rect 43346 24216 43352 24268
rect 43404 24256 43410 24268
rect 43993 24259 44051 24265
rect 43993 24256 44005 24259
rect 43404 24228 44005 24256
rect 43404 24216 43410 24228
rect 43993 24225 44005 24228
rect 44039 24225 44051 24259
rect 44174 24256 44180 24268
rect 44135 24228 44180 24256
rect 43993 24219 44051 24225
rect 44174 24216 44180 24228
rect 44232 24216 44238 24268
rect 31435 24160 32168 24188
rect 31435 24157 31447 24160
rect 31389 24151 31447 24157
rect 26068 24092 26924 24120
rect 26973 24123 27031 24129
rect 24084 24080 24090 24092
rect 26973 24089 26985 24123
rect 27019 24120 27031 24123
rect 27338 24120 27344 24132
rect 27019 24092 27344 24120
rect 27019 24089 27031 24092
rect 26973 24083 27031 24089
rect 27338 24080 27344 24092
rect 27396 24080 27402 24132
rect 28445 24123 28503 24129
rect 28445 24089 28457 24123
rect 28491 24089 28503 24123
rect 28445 24083 28503 24089
rect 30101 24123 30159 24129
rect 30101 24089 30113 24123
rect 30147 24120 30159 24123
rect 30742 24120 30748 24132
rect 30147 24092 30748 24120
rect 30147 24089 30159 24092
rect 30101 24083 30159 24089
rect 16942 24052 16948 24064
rect 16903 24024 16948 24052
rect 16942 24012 16948 24024
rect 17000 24012 17006 24064
rect 23566 24052 23572 24064
rect 23624 24061 23630 24064
rect 23533 24024 23572 24052
rect 23566 24012 23572 24024
rect 23624 24015 23633 24061
rect 26789 24055 26847 24061
rect 26789 24021 26801 24055
rect 26835 24052 26847 24055
rect 28460 24052 28488 24083
rect 30742 24080 30748 24092
rect 30800 24080 30806 24132
rect 31036 24120 31064 24151
rect 32214 24148 32220 24200
rect 32272 24188 32278 24200
rect 35897 24191 35955 24197
rect 32272 24160 32317 24188
rect 32272 24148 32278 24160
rect 35897 24157 35909 24191
rect 35943 24188 35955 24191
rect 37182 24188 37188 24200
rect 35943 24160 37188 24188
rect 35943 24157 35955 24160
rect 35897 24151 35955 24157
rect 37182 24148 37188 24160
rect 37240 24148 37246 24200
rect 37826 24188 37832 24200
rect 37787 24160 37832 24188
rect 37826 24148 37832 24160
rect 37884 24148 37890 24200
rect 38010 24188 38016 24200
rect 37971 24160 38016 24188
rect 38010 24148 38016 24160
rect 38068 24148 38074 24200
rect 40862 24188 40868 24200
rect 40823 24160 40868 24188
rect 40862 24148 40868 24160
rect 40920 24188 40926 24200
rect 41598 24188 41604 24200
rect 40920 24160 41604 24188
rect 40920 24148 40926 24160
rect 41598 24148 41604 24160
rect 41656 24148 41662 24200
rect 41690 24148 41696 24200
rect 41748 24188 41754 24200
rect 42426 24188 42432 24200
rect 41748 24160 42432 24188
rect 41748 24148 41754 24160
rect 42426 24148 42432 24160
rect 42484 24148 42490 24200
rect 31036 24092 31524 24120
rect 30558 24052 30564 24064
rect 26835 24024 30564 24052
rect 26835 24021 26847 24024
rect 26789 24015 26847 24021
rect 23624 24012 23630 24015
rect 30558 24012 30564 24024
rect 30616 24012 30622 24064
rect 30837 24055 30895 24061
rect 30837 24021 30849 24055
rect 30883 24052 30895 24055
rect 31294 24052 31300 24064
rect 30883 24024 31300 24052
rect 30883 24021 30895 24024
rect 30837 24015 30895 24021
rect 31294 24012 31300 24024
rect 31352 24012 31358 24064
rect 31496 24052 31524 24092
rect 31570 24080 31576 24132
rect 31628 24120 31634 24132
rect 31849 24123 31907 24129
rect 31849 24120 31861 24123
rect 31628 24092 31861 24120
rect 31628 24080 31634 24092
rect 31849 24089 31861 24092
rect 31895 24089 31907 24123
rect 36142 24123 36200 24129
rect 36142 24120 36154 24123
rect 31849 24083 31907 24089
rect 35912 24092 36154 24120
rect 35912 24064 35940 24092
rect 36142 24089 36154 24092
rect 36188 24089 36200 24123
rect 36142 24083 36200 24089
rect 38197 24123 38255 24129
rect 38197 24089 38209 24123
rect 38243 24120 38255 24123
rect 38746 24120 38752 24132
rect 38243 24092 38752 24120
rect 38243 24089 38255 24092
rect 38197 24083 38255 24089
rect 38746 24080 38752 24092
rect 38804 24080 38810 24132
rect 31662 24052 31668 24064
rect 31496 24024 31668 24052
rect 31662 24012 31668 24024
rect 31720 24012 31726 24064
rect 35894 24012 35900 24064
rect 35952 24012 35958 24064
rect 1104 23962 44896 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 44896 23962
rect 1104 23888 44896 23910
rect 17954 23848 17960 23860
rect 17915 23820 17960 23848
rect 17954 23808 17960 23820
rect 18012 23808 18018 23860
rect 19426 23848 19432 23860
rect 18340 23820 19432 23848
rect 18340 23789 18368 23820
rect 19426 23808 19432 23820
rect 19484 23808 19490 23860
rect 23566 23808 23572 23860
rect 23624 23808 23630 23860
rect 25041 23851 25099 23857
rect 25041 23817 25053 23851
rect 25087 23848 25099 23851
rect 25590 23848 25596 23860
rect 25087 23820 25596 23848
rect 25087 23817 25099 23820
rect 25041 23811 25099 23817
rect 25590 23808 25596 23820
rect 25648 23808 25654 23860
rect 26234 23808 26240 23860
rect 26292 23848 26298 23860
rect 27522 23848 27528 23860
rect 26292 23820 27528 23848
rect 26292 23808 26298 23820
rect 27522 23808 27528 23820
rect 27580 23848 27586 23860
rect 30466 23848 30472 23860
rect 27580 23820 29224 23848
rect 27580 23808 27586 23820
rect 18325 23783 18383 23789
rect 18325 23749 18337 23783
rect 18371 23749 18383 23783
rect 18325 23743 18383 23749
rect 18463 23783 18521 23789
rect 18463 23749 18475 23783
rect 18509 23780 18521 23783
rect 19702 23780 19708 23792
rect 18509 23752 19708 23780
rect 18509 23749 18521 23752
rect 18463 23743 18521 23749
rect 19702 23740 19708 23752
rect 19760 23740 19766 23792
rect 20438 23780 20444 23792
rect 20180 23752 20444 23780
rect 2130 23712 2136 23724
rect 2043 23684 2136 23712
rect 2130 23672 2136 23684
rect 2188 23712 2194 23724
rect 10962 23712 10968 23724
rect 2188 23684 10968 23712
rect 2188 23672 2194 23684
rect 10962 23672 10968 23684
rect 11020 23672 11026 23724
rect 15746 23672 15752 23724
rect 15804 23712 15810 23724
rect 15933 23715 15991 23721
rect 15933 23712 15945 23715
rect 15804 23684 15945 23712
rect 15804 23672 15810 23684
rect 15933 23681 15945 23684
rect 15979 23681 15991 23715
rect 15933 23675 15991 23681
rect 15948 23644 15976 23675
rect 16022 23672 16028 23724
rect 16080 23712 16086 23724
rect 16117 23715 16175 23721
rect 16117 23712 16129 23715
rect 16080 23684 16129 23712
rect 16080 23672 16086 23684
rect 16117 23681 16129 23684
rect 16163 23681 16175 23715
rect 17218 23712 17224 23724
rect 17179 23684 17224 23712
rect 16117 23675 16175 23681
rect 17218 23672 17224 23684
rect 17276 23672 17282 23724
rect 18138 23712 18144 23724
rect 18099 23684 18144 23712
rect 18138 23672 18144 23684
rect 18196 23672 18202 23724
rect 18230 23672 18236 23724
rect 18288 23712 18294 23724
rect 19061 23715 19119 23721
rect 19061 23712 19073 23715
rect 18288 23684 18333 23712
rect 18432 23684 19073 23712
rect 18288 23672 18294 23684
rect 16390 23644 16396 23656
rect 15948 23616 16396 23644
rect 16390 23604 16396 23616
rect 16448 23644 16454 23656
rect 17037 23647 17095 23653
rect 17037 23644 17049 23647
rect 16448 23616 17049 23644
rect 16448 23604 16454 23616
rect 17037 23613 17049 23616
rect 17083 23644 17095 23647
rect 18432 23644 18460 23684
rect 19061 23681 19073 23684
rect 19107 23681 19119 23715
rect 19061 23675 19119 23681
rect 19150 23672 19156 23724
rect 19208 23712 19214 23724
rect 19337 23715 19395 23721
rect 19208 23684 19253 23712
rect 19208 23672 19214 23684
rect 19337 23681 19349 23715
rect 19383 23712 19395 23715
rect 20070 23712 20076 23724
rect 19383 23684 20076 23712
rect 19383 23681 19395 23684
rect 19337 23675 19395 23681
rect 20070 23672 20076 23684
rect 20128 23672 20134 23724
rect 20180 23721 20208 23752
rect 20438 23740 20444 23752
rect 20496 23740 20502 23792
rect 22370 23780 22376 23792
rect 22331 23752 22376 23780
rect 22370 23740 22376 23752
rect 22428 23740 22434 23792
rect 23584 23780 23612 23808
rect 23906 23783 23964 23789
rect 23906 23780 23918 23783
rect 23584 23752 23918 23780
rect 23906 23749 23918 23752
rect 23952 23749 23964 23783
rect 23906 23743 23964 23749
rect 27617 23783 27675 23789
rect 27617 23749 27629 23783
rect 27663 23780 27675 23783
rect 27706 23780 27712 23792
rect 27663 23752 27712 23780
rect 27663 23749 27675 23752
rect 27617 23743 27675 23749
rect 27706 23740 27712 23752
rect 27764 23740 27770 23792
rect 28537 23783 28595 23789
rect 28537 23780 28549 23783
rect 27816 23752 28549 23780
rect 27816 23724 27844 23752
rect 28537 23749 28549 23752
rect 28583 23749 28595 23783
rect 28537 23743 28595 23749
rect 28718 23740 28724 23792
rect 28776 23740 28782 23792
rect 20165 23715 20223 23721
rect 20165 23681 20177 23715
rect 20211 23681 20223 23715
rect 20165 23675 20223 23681
rect 20349 23715 20407 23721
rect 20349 23681 20361 23715
rect 20395 23712 20407 23715
rect 20809 23715 20867 23721
rect 20809 23712 20821 23715
rect 20395 23684 20821 23712
rect 20395 23681 20407 23684
rect 20349 23675 20407 23681
rect 20809 23681 20821 23684
rect 20855 23681 20867 23715
rect 23658 23712 23664 23724
rect 23619 23684 23664 23712
rect 20809 23675 20867 23681
rect 23658 23672 23664 23684
rect 23716 23672 23722 23724
rect 27798 23712 27804 23724
rect 27759 23684 27804 23712
rect 27798 23672 27804 23684
rect 27856 23672 27862 23724
rect 27982 23672 27988 23724
rect 28040 23712 28046 23724
rect 28736 23712 28764 23740
rect 29196 23721 29224 23820
rect 30208 23820 30472 23848
rect 28040 23684 28764 23712
rect 29181 23715 29239 23721
rect 28040 23672 28046 23684
rect 29181 23681 29193 23715
rect 29227 23681 29239 23715
rect 29181 23675 29239 23681
rect 18598 23644 18604 23656
rect 17083 23616 18460 23644
rect 18511 23616 18604 23644
rect 17083 23613 17095 23616
rect 17037 23607 17095 23613
rect 2041 23579 2099 23585
rect 2041 23545 2053 23579
rect 2087 23576 2099 23579
rect 3050 23576 3056 23588
rect 2087 23548 3056 23576
rect 2087 23545 2099 23548
rect 2041 23539 2099 23545
rect 3050 23536 3056 23548
rect 3108 23536 3114 23588
rect 18432 23576 18460 23616
rect 18598 23604 18604 23616
rect 18656 23644 18662 23656
rect 19168 23644 19196 23672
rect 18656 23616 19196 23644
rect 19981 23647 20039 23653
rect 18656 23604 18662 23616
rect 19981 23613 19993 23647
rect 20027 23613 20039 23647
rect 19981 23607 20039 23613
rect 28721 23647 28779 23653
rect 28721 23613 28733 23647
rect 28767 23644 28779 23647
rect 30208 23644 30236 23820
rect 30466 23808 30472 23820
rect 30524 23808 30530 23860
rect 30926 23808 30932 23860
rect 30984 23848 30990 23860
rect 31570 23848 31576 23860
rect 30984 23820 31248 23848
rect 31531 23820 31576 23848
rect 30984 23808 30990 23820
rect 30374 23712 30380 23724
rect 30335 23684 30380 23712
rect 30374 23672 30380 23684
rect 30432 23672 30438 23724
rect 30558 23712 30564 23724
rect 30519 23684 30564 23712
rect 30558 23672 30564 23684
rect 30616 23672 30622 23724
rect 31110 23712 31116 23724
rect 31036 23684 31116 23712
rect 28767 23616 30236 23644
rect 30469 23647 30527 23653
rect 28767 23613 28779 23616
rect 28721 23607 28779 23613
rect 30469 23613 30481 23647
rect 30515 23644 30527 23647
rect 31036 23644 31064 23684
rect 31110 23672 31116 23684
rect 31168 23672 31174 23724
rect 31220 23721 31248 23820
rect 31570 23808 31576 23820
rect 31628 23808 31634 23860
rect 37645 23851 37703 23857
rect 37645 23817 37657 23851
rect 37691 23848 37703 23851
rect 37826 23848 37832 23860
rect 37691 23820 37832 23848
rect 37691 23817 37703 23820
rect 37645 23811 37703 23817
rect 37826 23808 37832 23820
rect 37884 23808 37890 23860
rect 38473 23851 38531 23857
rect 38473 23817 38485 23851
rect 38519 23848 38531 23851
rect 38562 23848 38568 23860
rect 38519 23820 38568 23848
rect 38519 23817 38531 23820
rect 38473 23811 38531 23817
rect 38562 23808 38568 23820
rect 38620 23808 38626 23860
rect 41049 23851 41107 23857
rect 41049 23817 41061 23851
rect 41095 23848 41107 23851
rect 42334 23848 42340 23860
rect 41095 23820 42340 23848
rect 41095 23817 41107 23820
rect 41049 23811 41107 23817
rect 42334 23808 42340 23820
rect 42392 23808 42398 23860
rect 42794 23808 42800 23860
rect 42852 23848 42858 23860
rect 43346 23848 43352 23860
rect 42852 23820 43352 23848
rect 42852 23808 42858 23820
rect 43346 23808 43352 23820
rect 43404 23808 43410 23860
rect 31662 23740 31668 23792
rect 31720 23780 31726 23792
rect 32217 23783 32275 23789
rect 32217 23780 32229 23783
rect 31720 23752 32229 23780
rect 31720 23740 31726 23752
rect 32217 23749 32229 23752
rect 32263 23749 32275 23783
rect 32217 23743 32275 23749
rect 31205 23715 31263 23721
rect 31205 23681 31217 23715
rect 31251 23681 31263 23715
rect 31205 23675 31263 23681
rect 31389 23715 31447 23721
rect 31389 23681 31401 23715
rect 31435 23712 31447 23715
rect 31938 23712 31944 23724
rect 31435 23684 31944 23712
rect 31435 23681 31447 23684
rect 31389 23675 31447 23681
rect 31938 23672 31944 23684
rect 31996 23672 32002 23724
rect 32125 23715 32183 23721
rect 32125 23681 32137 23715
rect 32171 23681 32183 23715
rect 32125 23675 32183 23681
rect 32309 23715 32367 23721
rect 32309 23681 32321 23715
rect 32355 23712 32367 23715
rect 32398 23712 32404 23724
rect 32355 23684 32404 23712
rect 32355 23681 32367 23684
rect 32309 23675 32367 23681
rect 30515 23616 31064 23644
rect 31220 23616 31524 23644
rect 30515 23613 30527 23616
rect 30469 23607 30527 23613
rect 19996 23576 20024 23607
rect 18432 23548 20024 23576
rect 22094 23536 22100 23588
rect 22152 23576 22158 23588
rect 22189 23579 22247 23585
rect 22189 23576 22201 23579
rect 22152 23548 22201 23576
rect 22152 23536 22158 23548
rect 22189 23545 22201 23548
rect 22235 23545 22247 23579
rect 22189 23539 22247 23545
rect 28534 23536 28540 23588
rect 28592 23576 28598 23588
rect 31220 23576 31248 23616
rect 28592 23548 31248 23576
rect 31297 23579 31355 23585
rect 28592 23536 28598 23548
rect 31297 23545 31309 23579
rect 31343 23576 31355 23579
rect 31386 23576 31392 23588
rect 31343 23548 31392 23576
rect 31343 23545 31355 23548
rect 31297 23539 31355 23545
rect 31386 23536 31392 23548
rect 31444 23536 31450 23588
rect 31496 23576 31524 23616
rect 31570 23604 31576 23656
rect 31628 23644 31634 23656
rect 32140 23644 32168 23675
rect 32398 23672 32404 23684
rect 32456 23672 32462 23724
rect 33597 23715 33655 23721
rect 33597 23681 33609 23715
rect 33643 23681 33655 23715
rect 34054 23712 34060 23724
rect 34015 23684 34060 23712
rect 33597 23675 33655 23681
rect 33318 23644 33324 23656
rect 31628 23616 32168 23644
rect 33279 23616 33324 23644
rect 31628 23604 31634 23616
rect 33318 23604 33324 23616
rect 33376 23604 33382 23656
rect 33612 23644 33640 23675
rect 34054 23672 34060 23684
rect 34112 23672 34118 23724
rect 34146 23672 34152 23724
rect 34204 23712 34210 23724
rect 34313 23715 34371 23721
rect 34313 23712 34325 23715
rect 34204 23684 34325 23712
rect 34204 23672 34210 23684
rect 34313 23681 34325 23684
rect 34359 23681 34371 23715
rect 35897 23715 35955 23721
rect 35897 23712 35909 23715
rect 34313 23675 34371 23681
rect 35452 23684 35909 23712
rect 33962 23644 33968 23656
rect 33612 23616 33968 23644
rect 33962 23604 33968 23616
rect 34020 23604 34026 23656
rect 33505 23579 33563 23585
rect 33505 23576 33517 23579
rect 31496 23548 33517 23576
rect 33505 23545 33517 23548
rect 33551 23576 33563 23579
rect 33870 23576 33876 23588
rect 33551 23548 33876 23576
rect 33551 23545 33563 23548
rect 33505 23539 33563 23545
rect 33870 23536 33876 23548
rect 33928 23536 33934 23588
rect 35452 23585 35480 23684
rect 35897 23681 35909 23684
rect 35943 23712 35955 23715
rect 36354 23712 36360 23724
rect 35943 23684 36360 23712
rect 35943 23681 35955 23684
rect 35897 23675 35955 23681
rect 36354 23672 36360 23684
rect 36412 23712 36418 23724
rect 37277 23715 37335 23721
rect 37277 23712 37289 23715
rect 36412 23684 37289 23712
rect 36412 23672 36418 23684
rect 37277 23681 37289 23684
rect 37323 23681 37335 23715
rect 37277 23675 37335 23681
rect 37366 23672 37372 23724
rect 37424 23712 37430 23724
rect 37461 23715 37519 23721
rect 37461 23712 37473 23715
rect 37424 23684 37473 23712
rect 37424 23672 37430 23684
rect 37461 23681 37473 23684
rect 37507 23681 37519 23715
rect 37461 23675 37519 23681
rect 38657 23715 38715 23721
rect 38657 23681 38669 23715
rect 38703 23712 38715 23715
rect 39022 23712 39028 23724
rect 38703 23684 39028 23712
rect 38703 23681 38715 23684
rect 38657 23675 38715 23681
rect 39022 23672 39028 23684
rect 39080 23672 39086 23724
rect 40865 23715 40923 23721
rect 40865 23681 40877 23715
rect 40911 23712 40923 23715
rect 41509 23715 41567 23721
rect 41509 23712 41521 23715
rect 40911 23684 41521 23712
rect 40911 23681 40923 23684
rect 40865 23675 40923 23681
rect 41509 23681 41521 23684
rect 41555 23681 41567 23715
rect 41509 23675 41567 23681
rect 41598 23672 41604 23724
rect 41656 23712 41662 23724
rect 41693 23715 41751 23721
rect 41693 23712 41705 23715
rect 41656 23684 41705 23712
rect 41656 23672 41662 23684
rect 41693 23681 41705 23684
rect 41739 23681 41751 23715
rect 41693 23675 41751 23681
rect 41782 23672 41788 23724
rect 41840 23712 41846 23724
rect 42613 23715 42671 23721
rect 41840 23684 41885 23712
rect 41840 23672 41846 23684
rect 42613 23681 42625 23715
rect 42659 23712 42671 23715
rect 42794 23712 42800 23724
rect 42659 23684 42800 23712
rect 42659 23681 42671 23684
rect 42613 23675 42671 23681
rect 42794 23672 42800 23684
rect 42852 23672 42858 23724
rect 43254 23712 43260 23724
rect 43215 23684 43260 23712
rect 43254 23672 43260 23684
rect 43312 23672 43318 23724
rect 35526 23604 35532 23656
rect 35584 23644 35590 23656
rect 36173 23647 36231 23653
rect 36173 23644 36185 23647
rect 35584 23616 36185 23644
rect 35584 23604 35590 23616
rect 36173 23613 36185 23616
rect 36219 23613 36231 23647
rect 38746 23644 38752 23656
rect 38707 23616 38752 23644
rect 36173 23607 36231 23613
rect 38746 23604 38752 23616
rect 38804 23604 38810 23656
rect 38838 23604 38844 23656
rect 38896 23644 38902 23656
rect 38896 23616 38941 23644
rect 38896 23604 38902 23616
rect 35437 23579 35495 23585
rect 35437 23545 35449 23579
rect 35483 23545 35495 23579
rect 35437 23539 35495 23545
rect 2774 23508 2780 23520
rect 2735 23480 2780 23508
rect 2774 23468 2780 23480
rect 2832 23468 2838 23520
rect 15930 23468 15936 23520
rect 15988 23508 15994 23520
rect 16025 23511 16083 23517
rect 16025 23508 16037 23511
rect 15988 23480 16037 23508
rect 15988 23468 15994 23480
rect 16025 23477 16037 23480
rect 16071 23477 16083 23511
rect 16025 23471 16083 23477
rect 19337 23511 19395 23517
rect 19337 23477 19349 23511
rect 19383 23508 19395 23511
rect 19978 23508 19984 23520
rect 19383 23480 19984 23508
rect 19383 23477 19395 23480
rect 19337 23471 19395 23477
rect 19978 23468 19984 23480
rect 20036 23468 20042 23520
rect 20993 23511 21051 23517
rect 20993 23477 21005 23511
rect 21039 23508 21051 23511
rect 21266 23508 21272 23520
rect 21039 23480 21272 23508
rect 21039 23477 21051 23480
rect 20993 23471 21051 23477
rect 21266 23468 21272 23480
rect 21324 23468 21330 23520
rect 27430 23468 27436 23520
rect 27488 23508 27494 23520
rect 29181 23511 29239 23517
rect 29181 23508 29193 23511
rect 27488 23480 29193 23508
rect 27488 23468 27494 23480
rect 29181 23477 29193 23480
rect 29227 23508 29239 23511
rect 29270 23508 29276 23520
rect 29227 23480 29276 23508
rect 29227 23477 29239 23480
rect 29181 23471 29239 23477
rect 29270 23468 29276 23480
rect 29328 23468 29334 23520
rect 30742 23468 30748 23520
rect 30800 23508 30806 23520
rect 31570 23508 31576 23520
rect 30800 23480 31576 23508
rect 30800 23468 30806 23480
rect 31570 23468 31576 23480
rect 31628 23468 31634 23520
rect 33410 23508 33416 23520
rect 33371 23480 33416 23508
rect 33410 23468 33416 23480
rect 33468 23468 33474 23520
rect 42334 23468 42340 23520
rect 42392 23508 42398 23520
rect 42429 23511 42487 23517
rect 42429 23508 42441 23511
rect 42392 23480 42441 23508
rect 42392 23468 42398 23480
rect 42429 23477 42441 23480
rect 42475 23477 42487 23511
rect 42429 23471 42487 23477
rect 42518 23468 42524 23520
rect 42576 23508 42582 23520
rect 43165 23511 43223 23517
rect 43165 23508 43177 23511
rect 42576 23480 43177 23508
rect 42576 23468 42582 23480
rect 43165 23477 43177 23480
rect 43211 23477 43223 23511
rect 43165 23471 43223 23477
rect 43901 23511 43959 23517
rect 43901 23477 43913 23511
rect 43947 23508 43959 23511
rect 44174 23508 44180 23520
rect 43947 23480 44180 23508
rect 43947 23477 43959 23480
rect 43901 23471 43959 23477
rect 44174 23468 44180 23480
rect 44232 23468 44238 23520
rect 1104 23418 44896 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 44896 23418
rect 1104 23344 44896 23366
rect 16761 23307 16819 23313
rect 16761 23273 16773 23307
rect 16807 23304 16819 23307
rect 17218 23304 17224 23316
rect 16807 23276 17224 23304
rect 16807 23273 16819 23276
rect 16761 23267 16819 23273
rect 17218 23264 17224 23276
rect 17276 23264 17282 23316
rect 23474 23264 23480 23316
rect 23532 23304 23538 23316
rect 23569 23307 23627 23313
rect 23569 23304 23581 23307
rect 23532 23276 23581 23304
rect 23532 23264 23538 23276
rect 23569 23273 23581 23276
rect 23615 23273 23627 23307
rect 23569 23267 23627 23273
rect 23661 23307 23719 23313
rect 23661 23273 23673 23307
rect 23707 23304 23719 23307
rect 23750 23304 23756 23316
rect 23707 23276 23756 23304
rect 23707 23273 23719 23276
rect 23661 23267 23719 23273
rect 23750 23264 23756 23276
rect 23808 23264 23814 23316
rect 25038 23264 25044 23316
rect 25096 23304 25102 23316
rect 25961 23307 26019 23313
rect 25961 23304 25973 23307
rect 25096 23276 25973 23304
rect 25096 23264 25102 23276
rect 25961 23273 25973 23276
rect 26007 23273 26019 23307
rect 25961 23267 26019 23273
rect 26329 23307 26387 23313
rect 26329 23273 26341 23307
rect 26375 23304 26387 23307
rect 26694 23304 26700 23316
rect 26375 23276 26700 23304
rect 26375 23273 26387 23276
rect 26329 23267 26387 23273
rect 26694 23264 26700 23276
rect 26752 23264 26758 23316
rect 26973 23307 27031 23313
rect 26973 23273 26985 23307
rect 27019 23304 27031 23307
rect 27798 23304 27804 23316
rect 27019 23276 27804 23304
rect 27019 23273 27031 23276
rect 26973 23267 27031 23273
rect 27798 23264 27804 23276
rect 27856 23264 27862 23316
rect 33597 23307 33655 23313
rect 33597 23273 33609 23307
rect 33643 23304 33655 23307
rect 34146 23304 34152 23316
rect 33643 23276 34152 23304
rect 33643 23273 33655 23276
rect 33597 23267 33655 23273
rect 34146 23264 34152 23276
rect 34204 23264 34210 23316
rect 36541 23307 36599 23313
rect 36541 23273 36553 23307
rect 36587 23304 36599 23307
rect 38010 23304 38016 23316
rect 36587 23276 38016 23304
rect 36587 23273 36599 23276
rect 36541 23267 36599 23273
rect 38010 23264 38016 23276
rect 38068 23264 38074 23316
rect 41325 23307 41383 23313
rect 41325 23273 41337 23307
rect 41371 23304 41383 23307
rect 41782 23304 41788 23316
rect 41371 23276 41788 23304
rect 41371 23273 41383 23276
rect 41325 23267 41383 23273
rect 41782 23264 41788 23276
rect 41840 23264 41846 23316
rect 19426 23196 19432 23248
rect 19484 23196 19490 23248
rect 30650 23196 30656 23248
rect 30708 23236 30714 23248
rect 31113 23239 31171 23245
rect 31113 23236 31125 23239
rect 30708 23208 31125 23236
rect 30708 23196 30714 23208
rect 31113 23205 31125 23208
rect 31159 23236 31171 23239
rect 35894 23236 35900 23248
rect 31159 23208 35900 23236
rect 31159 23205 31171 23208
rect 31113 23199 31171 23205
rect 35894 23196 35900 23208
rect 35952 23196 35958 23248
rect 1394 23168 1400 23180
rect 1355 23140 1400 23168
rect 1394 23128 1400 23140
rect 1452 23128 1458 23180
rect 2774 23128 2780 23180
rect 2832 23168 2838 23180
rect 3237 23171 3295 23177
rect 3237 23168 3249 23171
rect 2832 23140 3249 23168
rect 2832 23128 2838 23140
rect 3237 23137 3249 23140
rect 3283 23137 3295 23171
rect 3237 23131 3295 23137
rect 16942 23128 16948 23180
rect 17000 23168 17006 23180
rect 17405 23171 17463 23177
rect 17405 23168 17417 23171
rect 17000 23140 17417 23168
rect 17000 23128 17006 23140
rect 17405 23137 17417 23140
rect 17451 23137 17463 23171
rect 17405 23131 17463 23137
rect 17681 23171 17739 23177
rect 17681 23137 17693 23171
rect 17727 23168 17739 23171
rect 18046 23168 18052 23180
rect 17727 23140 18052 23168
rect 17727 23137 17739 23140
rect 17681 23131 17739 23137
rect 18046 23128 18052 23140
rect 18104 23168 18110 23180
rect 18598 23168 18604 23180
rect 18104 23140 18604 23168
rect 18104 23128 18110 23140
rect 18598 23128 18604 23140
rect 18656 23128 18662 23180
rect 19444 23168 19472 23196
rect 20438 23168 20444 23180
rect 19444 23140 20444 23168
rect 15381 23103 15439 23109
rect 15381 23069 15393 23103
rect 15427 23100 15439 23103
rect 15470 23100 15476 23112
rect 15427 23072 15476 23100
rect 15427 23069 15439 23072
rect 15381 23063 15439 23069
rect 15470 23060 15476 23072
rect 15528 23060 15534 23112
rect 19334 23060 19340 23112
rect 19392 23100 19398 23112
rect 19628 23109 19656 23140
rect 20438 23128 20444 23140
rect 20496 23128 20502 23180
rect 23477 23171 23535 23177
rect 23477 23137 23489 23171
rect 23523 23168 23535 23171
rect 23842 23168 23848 23180
rect 23523 23140 23848 23168
rect 23523 23137 23535 23140
rect 23477 23131 23535 23137
rect 23842 23128 23848 23140
rect 23900 23168 23906 23180
rect 24578 23168 24584 23180
rect 23900 23140 24584 23168
rect 23900 23128 23906 23140
rect 24578 23128 24584 23140
rect 24636 23128 24642 23180
rect 26237 23171 26295 23177
rect 26237 23137 26249 23171
rect 26283 23168 26295 23171
rect 26418 23168 26424 23180
rect 26283 23140 26424 23168
rect 26283 23137 26295 23140
rect 26237 23131 26295 23137
rect 26418 23128 26424 23140
rect 26476 23128 26482 23180
rect 27338 23168 27344 23180
rect 26896 23140 27344 23168
rect 19429 23103 19487 23109
rect 19429 23100 19441 23103
rect 19392 23072 19441 23100
rect 19392 23060 19398 23072
rect 19429 23069 19441 23072
rect 19475 23069 19487 23103
rect 19429 23063 19487 23069
rect 19613 23103 19671 23109
rect 19613 23069 19625 23103
rect 19659 23069 19671 23103
rect 19613 23063 19671 23069
rect 19702 23060 19708 23112
rect 19760 23109 19766 23112
rect 19760 23103 19789 23109
rect 19777 23069 19789 23103
rect 19760 23063 19789 23069
rect 19889 23103 19947 23109
rect 19889 23069 19901 23103
rect 19935 23100 19947 23103
rect 20070 23100 20076 23112
rect 19935 23072 20076 23100
rect 19935 23069 19947 23072
rect 19889 23063 19947 23069
rect 19760 23060 19766 23063
rect 20070 23060 20076 23072
rect 20128 23060 20134 23112
rect 21266 23109 21272 23112
rect 20993 23103 21051 23109
rect 20993 23069 21005 23103
rect 21039 23069 21051 23103
rect 20993 23063 21051 23069
rect 21260 23063 21272 23109
rect 21324 23100 21330 23112
rect 23753 23103 23811 23109
rect 21324 23072 21360 23100
rect 3050 23032 3056 23044
rect 3011 23004 3056 23032
rect 3050 22992 3056 23004
rect 3108 22992 3114 23044
rect 15654 23041 15660 23044
rect 15648 22995 15660 23041
rect 15712 23032 15718 23044
rect 15712 23004 15748 23032
rect 15654 22992 15660 22995
rect 15712 22992 15718 23004
rect 18230 22992 18236 23044
rect 18288 23032 18294 23044
rect 19521 23035 19579 23041
rect 19521 23032 19533 23035
rect 18288 23004 19533 23032
rect 18288 22992 18294 23004
rect 19521 23001 19533 23004
rect 19567 23001 19579 23035
rect 19720 23032 19748 23060
rect 20346 23032 20352 23044
rect 19720 23004 20352 23032
rect 19521 22995 19579 23001
rect 20346 22992 20352 23004
rect 20404 22992 20410 23044
rect 19242 22964 19248 22976
rect 19203 22936 19248 22964
rect 19242 22924 19248 22936
rect 19300 22924 19306 22976
rect 21008 22964 21036 23063
rect 21266 23060 21272 23063
rect 21324 23060 21330 23072
rect 23753 23069 23765 23103
rect 23799 23100 23811 23103
rect 24026 23100 24032 23112
rect 23799 23072 24032 23100
rect 23799 23069 23811 23072
rect 23753 23063 23811 23069
rect 24026 23060 24032 23072
rect 24084 23060 24090 23112
rect 24394 23100 24400 23112
rect 24307 23072 24400 23100
rect 24394 23060 24400 23072
rect 24452 23100 24458 23112
rect 24854 23100 24860 23112
rect 24452 23072 24860 23100
rect 24452 23060 24458 23072
rect 24854 23060 24860 23072
rect 24912 23060 24918 23112
rect 26896 23109 26924 23140
rect 27338 23128 27344 23140
rect 27396 23168 27402 23180
rect 28353 23171 28411 23177
rect 28353 23168 28365 23171
rect 27396 23140 28365 23168
rect 27396 23128 27402 23140
rect 28353 23137 28365 23140
rect 28399 23137 28411 23171
rect 30374 23168 30380 23180
rect 28353 23131 28411 23137
rect 30208 23140 30380 23168
rect 26329 23103 26387 23109
rect 26329 23069 26341 23103
rect 26375 23069 26387 23103
rect 26329 23063 26387 23069
rect 26881 23103 26939 23109
rect 26881 23069 26893 23103
rect 26927 23069 26939 23103
rect 28074 23100 28080 23112
rect 28035 23072 28080 23100
rect 26881 23063 26939 23069
rect 23566 23032 23572 23044
rect 22066 23004 23572 23032
rect 21450 22964 21456 22976
rect 21008 22936 21456 22964
rect 21450 22924 21456 22936
rect 21508 22964 21514 22976
rect 22066 22964 22094 23004
rect 23566 22992 23572 23004
rect 23624 22992 23630 23044
rect 26234 22992 26240 23044
rect 26292 23032 26298 23044
rect 26344 23032 26372 23063
rect 28074 23060 28080 23072
rect 28132 23060 28138 23112
rect 30208 23109 30236 23140
rect 30374 23128 30380 23140
rect 30432 23168 30438 23180
rect 30926 23168 30932 23180
rect 30432 23140 30932 23168
rect 30432 23128 30438 23140
rect 30926 23128 30932 23140
rect 30984 23128 30990 23180
rect 37093 23171 37151 23177
rect 37093 23137 37105 23171
rect 37139 23168 37151 23171
rect 37826 23168 37832 23180
rect 37139 23140 37832 23168
rect 37139 23137 37151 23140
rect 37093 23131 37151 23137
rect 37826 23128 37832 23140
rect 37884 23128 37890 23180
rect 39942 23168 39948 23180
rect 39903 23140 39948 23168
rect 39942 23128 39948 23140
rect 40000 23128 40006 23180
rect 42702 23168 42708 23180
rect 42663 23140 42708 23168
rect 42702 23128 42708 23140
rect 42760 23128 42766 23180
rect 44174 23168 44180 23180
rect 44135 23140 44180 23168
rect 44174 23128 44180 23140
rect 44232 23128 44238 23180
rect 30193 23103 30251 23109
rect 30193 23069 30205 23103
rect 30239 23069 30251 23103
rect 30837 23103 30895 23109
rect 30837 23100 30849 23103
rect 30193 23063 30251 23069
rect 30300 23072 30849 23100
rect 30006 23032 30012 23044
rect 26292 23004 26372 23032
rect 29967 23004 30012 23032
rect 26292 22992 26298 23004
rect 30006 22992 30012 23004
rect 30064 23032 30070 23044
rect 30300 23032 30328 23072
rect 30837 23069 30849 23072
rect 30883 23069 30895 23103
rect 31018 23100 31024 23112
rect 30979 23072 31024 23100
rect 30837 23063 30895 23069
rect 31018 23060 31024 23072
rect 31076 23060 31082 23112
rect 33410 23060 33416 23112
rect 33468 23100 33474 23112
rect 33597 23103 33655 23109
rect 33597 23100 33609 23103
rect 33468 23072 33609 23100
rect 33468 23060 33474 23072
rect 33597 23069 33609 23072
rect 33643 23069 33655 23103
rect 33870 23100 33876 23112
rect 33831 23072 33876 23100
rect 33597 23063 33655 23069
rect 33870 23060 33876 23072
rect 33928 23100 33934 23112
rect 34422 23100 34428 23112
rect 33928 23072 34428 23100
rect 33928 23060 33934 23072
rect 34422 23060 34428 23072
rect 34480 23060 34486 23112
rect 36354 23100 36360 23112
rect 36315 23072 36360 23100
rect 36354 23060 36360 23072
rect 36412 23060 36418 23112
rect 36541 23103 36599 23109
rect 36541 23069 36553 23103
rect 36587 23069 36599 23103
rect 36541 23063 36599 23069
rect 37185 23103 37243 23109
rect 37185 23069 37197 23103
rect 37231 23100 37243 23103
rect 37642 23100 37648 23112
rect 37231 23072 37648 23100
rect 37231 23069 37243 23072
rect 37185 23063 37243 23069
rect 30064 23004 30328 23032
rect 30377 23035 30435 23041
rect 30064 22992 30070 23004
rect 30377 23001 30389 23035
rect 30423 23032 30435 23035
rect 31386 23032 31392 23044
rect 30423 23004 31392 23032
rect 30423 23001 30435 23004
rect 30377 22995 30435 23001
rect 21508 22936 22094 22964
rect 22373 22967 22431 22973
rect 21508 22924 21514 22936
rect 22373 22933 22385 22967
rect 22419 22964 22431 22967
rect 23290 22964 23296 22976
rect 22419 22936 23296 22964
rect 22419 22933 22431 22936
rect 22373 22927 22431 22933
rect 23290 22924 23296 22936
rect 23348 22924 23354 22976
rect 24578 22964 24584 22976
rect 24539 22936 24584 22964
rect 24578 22924 24584 22936
rect 24636 22924 24642 22976
rect 30190 22924 30196 22976
rect 30248 22964 30254 22976
rect 30392 22964 30420 22995
rect 31386 22992 31392 23004
rect 31444 22992 31450 23044
rect 36556 23032 36584 23063
rect 37642 23060 37648 23072
rect 37700 23060 37706 23112
rect 38657 23103 38715 23109
rect 38657 23069 38669 23103
rect 38703 23100 38715 23103
rect 38746 23100 38752 23112
rect 38703 23072 38752 23100
rect 38703 23069 38715 23072
rect 38657 23063 38715 23069
rect 38746 23060 38752 23072
rect 38804 23060 38810 23112
rect 38838 23060 38844 23112
rect 38896 23100 38902 23112
rect 38896 23072 38989 23100
rect 38896 23060 38902 23072
rect 39022 23060 39028 23112
rect 39080 23100 39086 23112
rect 39117 23103 39175 23109
rect 39117 23100 39129 23103
rect 39080 23072 39129 23100
rect 39080 23060 39086 23072
rect 39117 23069 39129 23072
rect 39163 23069 39175 23103
rect 39117 23063 39175 23069
rect 37366 23032 37372 23044
rect 36556 23004 37372 23032
rect 37366 22992 37372 23004
rect 37424 22992 37430 23044
rect 38856 23032 38884 23060
rect 38212 23004 38884 23032
rect 39301 23035 39359 23041
rect 38212 22976 38240 23004
rect 39301 23001 39313 23035
rect 39347 23032 39359 23035
rect 40190 23035 40248 23041
rect 40190 23032 40202 23035
rect 39347 23004 40202 23032
rect 39347 23001 39359 23004
rect 39301 22995 39359 23001
rect 40190 23001 40202 23004
rect 40236 23001 40248 23035
rect 40190 22995 40248 23001
rect 43438 22992 43444 23044
rect 43496 23032 43502 23044
rect 43993 23035 44051 23041
rect 43993 23032 44005 23035
rect 43496 23004 44005 23032
rect 43496 22992 43502 23004
rect 43993 23001 44005 23004
rect 44039 23001 44051 23035
rect 43993 22995 44051 23001
rect 30248 22936 30420 22964
rect 33781 22967 33839 22973
rect 30248 22924 30254 22936
rect 33781 22933 33793 22967
rect 33827 22964 33839 22967
rect 33962 22964 33968 22976
rect 33827 22936 33968 22964
rect 33827 22933 33839 22936
rect 33781 22927 33839 22933
rect 33962 22924 33968 22936
rect 34020 22924 34026 22976
rect 37553 22967 37611 22973
rect 37553 22933 37565 22967
rect 37599 22964 37611 22967
rect 38194 22964 38200 22976
rect 37599 22936 38200 22964
rect 37599 22933 37611 22936
rect 37553 22927 37611 22933
rect 38194 22924 38200 22936
rect 38252 22924 38258 22976
rect 1104 22874 44896 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 44896 22874
rect 1104 22800 44896 22822
rect 15470 22720 15476 22772
rect 15528 22760 15534 22772
rect 15528 22732 18736 22760
rect 15528 22720 15534 22732
rect 16929 22695 16987 22701
rect 16929 22661 16941 22695
rect 16975 22692 16987 22695
rect 17129 22695 17187 22701
rect 16975 22664 17080 22692
rect 16975 22661 16987 22664
rect 16929 22655 16987 22661
rect 6362 22624 6368 22636
rect 6323 22596 6368 22624
rect 6362 22584 6368 22596
rect 6420 22584 6426 22636
rect 15746 22624 15752 22636
rect 15707 22596 15752 22624
rect 15746 22584 15752 22596
rect 15804 22584 15810 22636
rect 15841 22627 15899 22633
rect 15841 22593 15853 22627
rect 15887 22593 15899 22627
rect 15841 22587 15899 22593
rect 1946 22556 1952 22568
rect 1907 22528 1952 22556
rect 1946 22516 1952 22528
rect 2004 22516 2010 22568
rect 2133 22559 2191 22565
rect 2133 22525 2145 22559
rect 2179 22556 2191 22559
rect 2866 22556 2872 22568
rect 2179 22528 2872 22556
rect 2179 22525 2191 22528
rect 2133 22519 2191 22525
rect 2866 22516 2872 22528
rect 2924 22516 2930 22568
rect 2958 22516 2964 22568
rect 3016 22556 3022 22568
rect 3016 22528 3061 22556
rect 3016 22516 3022 22528
rect 6178 22516 6184 22568
rect 6236 22556 6242 22568
rect 6549 22559 6607 22565
rect 6549 22556 6561 22559
rect 6236 22528 6561 22556
rect 6236 22516 6242 22528
rect 6549 22525 6561 22528
rect 6595 22525 6607 22559
rect 6549 22519 6607 22525
rect 15473 22559 15531 22565
rect 15473 22525 15485 22559
rect 15519 22556 15531 22559
rect 15654 22556 15660 22568
rect 15519 22528 15660 22556
rect 15519 22525 15531 22528
rect 15473 22519 15531 22525
rect 15654 22516 15660 22528
rect 15712 22516 15718 22568
rect 15856 22556 15884 22587
rect 15930 22584 15936 22636
rect 15988 22624 15994 22636
rect 15988 22596 16033 22624
rect 15988 22584 15994 22596
rect 16114 22584 16120 22636
rect 16172 22624 16178 22636
rect 17052 22624 17080 22664
rect 17129 22661 17141 22695
rect 17175 22692 17187 22695
rect 18708 22692 18736 22732
rect 19150 22720 19156 22772
rect 19208 22760 19214 22772
rect 19208 22732 20760 22760
rect 19208 22720 19214 22732
rect 19426 22692 19432 22704
rect 17175 22664 18644 22692
rect 17175 22661 17187 22664
rect 17129 22655 17187 22661
rect 17218 22624 17224 22636
rect 16172 22596 16217 22624
rect 17052 22596 17224 22624
rect 16172 22584 16178 22596
rect 17218 22584 17224 22596
rect 17276 22624 17282 22636
rect 17589 22627 17647 22633
rect 17589 22624 17601 22627
rect 17276 22596 17601 22624
rect 17276 22584 17282 22596
rect 17589 22593 17601 22596
rect 17635 22593 17647 22627
rect 17770 22624 17776 22636
rect 17731 22596 17776 22624
rect 17589 22587 17647 22593
rect 17770 22584 17776 22596
rect 17828 22584 17834 22636
rect 16298 22556 16304 22568
rect 15856 22528 16304 22556
rect 16298 22516 16304 22528
rect 16356 22516 16362 22568
rect 18046 22488 18052 22500
rect 17788 22460 18052 22488
rect 16666 22380 16672 22432
rect 16724 22420 16730 22432
rect 16761 22423 16819 22429
rect 16761 22420 16773 22423
rect 16724 22392 16773 22420
rect 16724 22380 16730 22392
rect 16761 22389 16773 22392
rect 16807 22389 16819 22423
rect 16942 22420 16948 22432
rect 16903 22392 16948 22420
rect 16761 22383 16819 22389
rect 16942 22380 16948 22392
rect 17000 22380 17006 22432
rect 17788 22429 17816 22460
rect 18046 22448 18052 22460
rect 18104 22448 18110 22500
rect 18616 22488 18644 22664
rect 18708 22664 19432 22692
rect 18708 22633 18736 22664
rect 19426 22652 19432 22664
rect 19484 22652 19490 22704
rect 18693 22627 18751 22633
rect 18693 22593 18705 22627
rect 18739 22593 18751 22627
rect 18693 22587 18751 22593
rect 18960 22627 19018 22633
rect 18960 22593 18972 22627
rect 19006 22624 19018 22627
rect 19242 22624 19248 22636
rect 19006 22596 19248 22624
rect 19006 22593 19018 22596
rect 18960 22587 19018 22593
rect 19242 22584 19248 22596
rect 19300 22584 19306 22636
rect 20732 22633 20760 22732
rect 24578 22720 24584 22772
rect 24636 22760 24642 22772
rect 33318 22760 33324 22772
rect 24636 22732 33324 22760
rect 24636 22720 24642 22732
rect 33318 22720 33324 22732
rect 33376 22720 33382 22772
rect 39393 22763 39451 22769
rect 33428 22732 36584 22760
rect 22649 22695 22707 22701
rect 22649 22661 22661 22695
rect 22695 22692 22707 22695
rect 23566 22692 23572 22704
rect 22695 22664 23572 22692
rect 22695 22661 22707 22664
rect 22649 22655 22707 22661
rect 23566 22652 23572 22664
rect 23624 22652 23630 22704
rect 25222 22652 25228 22704
rect 25280 22692 25286 22704
rect 25501 22695 25559 22701
rect 25501 22692 25513 22695
rect 25280 22664 25513 22692
rect 25280 22652 25286 22664
rect 25501 22661 25513 22664
rect 25547 22661 25559 22695
rect 26694 22692 26700 22704
rect 25501 22655 25559 22661
rect 25884 22664 26700 22692
rect 20717 22627 20775 22633
rect 20717 22593 20729 22627
rect 20763 22593 20775 22627
rect 20717 22587 20775 22593
rect 20806 22584 20812 22636
rect 20864 22624 20870 22636
rect 20901 22627 20959 22633
rect 20901 22624 20913 22627
rect 20864 22596 20913 22624
rect 20864 22584 20870 22596
rect 20901 22593 20913 22596
rect 20947 22593 20959 22627
rect 22462 22624 22468 22636
rect 22423 22596 22468 22624
rect 20901 22587 20959 22593
rect 22462 22584 22468 22596
rect 22520 22584 22526 22636
rect 23477 22627 23535 22633
rect 23477 22593 23489 22627
rect 23523 22624 23535 22627
rect 24394 22624 24400 22636
rect 23523 22596 24400 22624
rect 23523 22593 23535 22596
rect 23477 22587 23535 22593
rect 23584 22568 23612 22596
rect 24394 22584 24400 22596
rect 24452 22584 24458 22636
rect 25884 22633 25912 22664
rect 26694 22652 26700 22664
rect 26752 22652 26758 22704
rect 27062 22652 27068 22704
rect 27120 22692 27126 22704
rect 27522 22692 27528 22704
rect 27120 22664 27528 22692
rect 27120 22652 27126 22664
rect 27522 22652 27528 22664
rect 27580 22692 27586 22704
rect 28813 22695 28871 22701
rect 28813 22692 28825 22695
rect 27580 22664 28825 22692
rect 27580 22652 27586 22664
rect 28813 22661 28825 22664
rect 28859 22661 28871 22695
rect 29917 22695 29975 22701
rect 29917 22692 29929 22695
rect 28813 22655 28871 22661
rect 29196 22664 29929 22692
rect 25869 22627 25927 22633
rect 25869 22593 25881 22627
rect 25915 22593 25927 22627
rect 25869 22587 25927 22593
rect 26145 22627 26203 22633
rect 26145 22593 26157 22627
rect 26191 22624 26203 22627
rect 26418 22624 26424 22636
rect 26191 22596 26424 22624
rect 26191 22593 26203 22596
rect 26145 22587 26203 22593
rect 26418 22584 26424 22596
rect 26476 22624 26482 22636
rect 27246 22624 27252 22636
rect 26476 22596 27252 22624
rect 26476 22584 26482 22596
rect 27246 22584 27252 22596
rect 27304 22584 27310 22636
rect 27801 22627 27859 22633
rect 27801 22593 27813 22627
rect 27847 22624 27859 22627
rect 27982 22624 27988 22636
rect 27847 22596 27988 22624
rect 27847 22593 27859 22596
rect 27801 22587 27859 22593
rect 27982 22584 27988 22596
rect 28040 22584 28046 22636
rect 28626 22584 28632 22636
rect 28684 22624 28690 22636
rect 29196 22633 29224 22664
rect 29917 22661 29929 22664
rect 29963 22661 29975 22695
rect 29917 22655 29975 22661
rect 31386 22652 31392 22704
rect 31444 22692 31450 22704
rect 33428 22692 33456 22732
rect 31444 22664 33456 22692
rect 33505 22695 33563 22701
rect 31444 22652 31450 22664
rect 33505 22661 33517 22695
rect 33551 22692 33563 22695
rect 34149 22695 34207 22701
rect 34149 22692 34161 22695
rect 33551 22664 34161 22692
rect 33551 22661 33563 22664
rect 33505 22655 33563 22661
rect 34149 22661 34161 22664
rect 34195 22661 34207 22695
rect 34149 22655 34207 22661
rect 34348 22664 35756 22692
rect 34348 22636 34376 22664
rect 28905 22627 28963 22633
rect 28905 22624 28917 22627
rect 28684 22596 28917 22624
rect 28684 22584 28690 22596
rect 28905 22593 28917 22596
rect 28951 22593 28963 22627
rect 28905 22587 28963 22593
rect 29181 22627 29239 22633
rect 29181 22593 29193 22627
rect 29227 22593 29239 22627
rect 29822 22624 29828 22636
rect 29783 22596 29828 22624
rect 29181 22587 29239 22593
rect 29822 22584 29828 22596
rect 29880 22584 29886 22636
rect 30561 22627 30619 22633
rect 30561 22593 30573 22627
rect 30607 22593 30619 22627
rect 30561 22587 30619 22593
rect 23566 22516 23572 22568
rect 23624 22516 23630 22568
rect 25685 22559 25743 22565
rect 25685 22525 25697 22559
rect 25731 22556 25743 22559
rect 26234 22556 26240 22568
rect 25731 22528 26240 22556
rect 25731 22525 25743 22528
rect 25685 22519 25743 22525
rect 26234 22516 26240 22528
rect 26292 22516 26298 22568
rect 27522 22556 27528 22568
rect 27483 22528 27528 22556
rect 27522 22516 27528 22528
rect 27580 22516 27586 22568
rect 29365 22559 29423 22565
rect 29365 22525 29377 22559
rect 29411 22556 29423 22559
rect 30006 22556 30012 22568
rect 29411 22528 30012 22556
rect 29411 22525 29423 22528
rect 29365 22519 29423 22525
rect 30006 22516 30012 22528
rect 30064 22556 30070 22568
rect 30576 22556 30604 22587
rect 30742 22584 30748 22636
rect 30800 22624 30806 22636
rect 30837 22627 30895 22633
rect 30837 22624 30849 22627
rect 30800 22596 30849 22624
rect 30800 22584 30806 22596
rect 30837 22593 30849 22596
rect 30883 22624 30895 22627
rect 30926 22624 30932 22636
rect 30883 22596 30932 22624
rect 30883 22593 30895 22596
rect 30837 22587 30895 22593
rect 30926 22584 30932 22596
rect 30984 22584 30990 22636
rect 31938 22624 31944 22636
rect 31726 22596 31944 22624
rect 30064 22528 30604 22556
rect 30064 22516 30070 22528
rect 18616 22460 18736 22488
rect 17773 22423 17831 22429
rect 17773 22389 17785 22423
rect 17819 22389 17831 22423
rect 17773 22383 17831 22389
rect 17957 22423 18015 22429
rect 17957 22389 17969 22423
rect 18003 22420 18015 22423
rect 18598 22420 18604 22432
rect 18003 22392 18604 22420
rect 18003 22389 18015 22392
rect 17957 22383 18015 22389
rect 18598 22380 18604 22392
rect 18656 22380 18662 22432
rect 18708 22420 18736 22460
rect 20438 22448 20444 22500
rect 20496 22488 20502 22500
rect 23293 22491 23351 22497
rect 23293 22488 23305 22491
rect 20496 22460 23305 22488
rect 20496 22448 20502 22460
rect 23293 22457 23305 22460
rect 23339 22457 23351 22491
rect 23293 22451 23351 22457
rect 31113 22491 31171 22497
rect 31113 22457 31125 22491
rect 31159 22488 31171 22491
rect 31726 22488 31754 22596
rect 31938 22584 31944 22596
rect 31996 22624 32002 22636
rect 32401 22627 32459 22633
rect 32401 22624 32413 22627
rect 31996 22596 32413 22624
rect 31996 22584 32002 22596
rect 32401 22593 32413 22596
rect 32447 22593 32459 22627
rect 32401 22587 32459 22593
rect 32585 22627 32643 22633
rect 32585 22593 32597 22627
rect 32631 22593 32643 22627
rect 34330 22624 34336 22636
rect 34243 22596 34336 22624
rect 32585 22587 32643 22593
rect 32600 22556 32628 22587
rect 34330 22584 34336 22596
rect 34388 22584 34394 22636
rect 34517 22627 34575 22633
rect 34517 22593 34529 22627
rect 34563 22593 34575 22627
rect 34517 22587 34575 22593
rect 32600 22528 33916 22556
rect 33134 22488 33140 22500
rect 31159 22460 31754 22488
rect 33047 22460 33140 22488
rect 31159 22457 31171 22460
rect 31113 22451 31171 22457
rect 33134 22448 33140 22460
rect 33192 22488 33198 22500
rect 33778 22488 33784 22500
rect 33192 22460 33784 22488
rect 33192 22448 33198 22460
rect 33778 22448 33784 22460
rect 33836 22448 33842 22500
rect 33888 22488 33916 22528
rect 33962 22516 33968 22568
rect 34020 22556 34026 22568
rect 34532 22556 34560 22587
rect 34606 22584 34612 22636
rect 34664 22624 34670 22636
rect 35728 22633 35756 22664
rect 35894 22652 35900 22704
rect 35952 22652 35958 22704
rect 35713 22627 35771 22633
rect 34664 22596 34709 22624
rect 34664 22584 34670 22596
rect 35713 22593 35725 22627
rect 35759 22593 35771 22627
rect 35912 22624 35940 22652
rect 36556 22633 36584 22732
rect 39393 22729 39405 22763
rect 39439 22760 39451 22763
rect 40034 22760 40040 22772
rect 39439 22732 40040 22760
rect 39439 22729 39451 22732
rect 39393 22723 39451 22729
rect 40034 22720 40040 22732
rect 40092 22720 40098 22772
rect 42794 22760 42800 22772
rect 42755 22732 42800 22760
rect 42794 22720 42800 22732
rect 42852 22720 42858 22772
rect 43438 22760 43444 22772
rect 43399 22732 43444 22760
rect 43438 22720 43444 22732
rect 43496 22720 43502 22772
rect 38838 22652 38844 22704
rect 38896 22692 38902 22704
rect 39022 22692 39028 22704
rect 38896 22664 39028 22692
rect 38896 22652 38902 22664
rect 39022 22652 39028 22664
rect 39080 22652 39086 22704
rect 35713 22587 35771 22593
rect 35820 22596 35940 22624
rect 36541 22627 36599 22633
rect 35526 22556 35532 22568
rect 34020 22528 35532 22556
rect 34020 22516 34026 22528
rect 35526 22516 35532 22528
rect 35584 22516 35590 22568
rect 35820 22565 35848 22596
rect 36541 22593 36553 22627
rect 36587 22593 36599 22627
rect 36541 22587 36599 22593
rect 36725 22627 36783 22633
rect 36725 22593 36737 22627
rect 36771 22624 36783 22627
rect 37642 22624 37648 22636
rect 36771 22596 37648 22624
rect 36771 22593 36783 22596
rect 36725 22587 36783 22593
rect 35805 22559 35863 22565
rect 35805 22525 35817 22559
rect 35851 22525 35863 22559
rect 35805 22519 35863 22525
rect 35894 22516 35900 22568
rect 35952 22556 35958 22568
rect 36633 22559 36691 22565
rect 36633 22556 36645 22559
rect 35952 22528 36645 22556
rect 35952 22516 35958 22528
rect 36633 22525 36645 22528
rect 36679 22525 36691 22559
rect 36633 22519 36691 22525
rect 34790 22488 34796 22500
rect 33888 22460 34796 22488
rect 34790 22448 34796 22460
rect 34848 22448 34854 22500
rect 36081 22491 36139 22497
rect 36081 22457 36093 22491
rect 36127 22488 36139 22491
rect 36740 22488 36768 22587
rect 37642 22584 37648 22596
rect 37700 22584 37706 22636
rect 38194 22624 38200 22636
rect 38155 22596 38200 22624
rect 38194 22584 38200 22596
rect 38252 22624 38258 22636
rect 38933 22627 38991 22633
rect 38933 22624 38945 22627
rect 38252 22596 38945 22624
rect 38252 22584 38258 22596
rect 38933 22593 38945 22596
rect 38979 22593 38991 22627
rect 38933 22587 38991 22593
rect 39114 22584 39120 22636
rect 39172 22624 39178 22636
rect 39209 22627 39267 22633
rect 39209 22624 39221 22627
rect 39172 22596 39221 22624
rect 39172 22584 39178 22596
rect 39209 22593 39221 22596
rect 39255 22593 39267 22627
rect 39209 22587 39267 22593
rect 41598 22584 41604 22636
rect 41656 22624 41662 22636
rect 42613 22627 42671 22633
rect 42613 22624 42625 22627
rect 41656 22596 42625 22624
rect 41656 22584 41662 22596
rect 42613 22593 42625 22596
rect 42659 22593 42671 22627
rect 42613 22587 42671 22593
rect 43070 22584 43076 22636
rect 43128 22624 43134 22636
rect 43349 22627 43407 22633
rect 43349 22624 43361 22627
rect 43128 22596 43361 22624
rect 43128 22584 43134 22596
rect 43349 22593 43361 22596
rect 43395 22593 43407 22627
rect 43349 22587 43407 22593
rect 38289 22559 38347 22565
rect 38289 22525 38301 22559
rect 38335 22525 38347 22559
rect 38289 22519 38347 22525
rect 38381 22559 38439 22565
rect 38381 22525 38393 22559
rect 38427 22556 38439 22559
rect 38838 22556 38844 22568
rect 38427 22528 38844 22556
rect 38427 22525 38439 22528
rect 38381 22519 38439 22525
rect 36127 22460 36768 22488
rect 38304 22488 38332 22519
rect 38838 22516 38844 22528
rect 38896 22516 38902 22568
rect 42426 22556 42432 22568
rect 42387 22528 42432 22556
rect 42426 22516 42432 22528
rect 42484 22516 42490 22568
rect 38746 22488 38752 22500
rect 38304 22460 38752 22488
rect 36127 22457 36139 22460
rect 36081 22451 36139 22457
rect 38746 22448 38752 22460
rect 38804 22448 38810 22500
rect 20070 22420 20076 22432
rect 18708 22392 20076 22420
rect 20070 22380 20076 22392
rect 20128 22420 20134 22432
rect 20622 22420 20628 22432
rect 20128 22392 20628 22420
rect 20128 22380 20134 22392
rect 20622 22380 20628 22392
rect 20680 22380 20686 22432
rect 20898 22380 20904 22432
rect 20956 22420 20962 22432
rect 21085 22423 21143 22429
rect 21085 22420 21097 22423
rect 20956 22392 21097 22420
rect 20956 22380 20962 22392
rect 21085 22389 21097 22392
rect 21131 22389 21143 22423
rect 21085 22383 21143 22389
rect 30466 22380 30472 22432
rect 30524 22420 30530 22432
rect 30653 22423 30711 22429
rect 30653 22420 30665 22423
rect 30524 22392 30665 22420
rect 30524 22380 30530 22392
rect 30653 22389 30665 22392
rect 30699 22389 30711 22423
rect 30653 22383 30711 22389
rect 32401 22423 32459 22429
rect 32401 22389 32413 22423
rect 32447 22420 32459 22423
rect 32766 22420 32772 22432
rect 32447 22392 32772 22420
rect 32447 22389 32459 22392
rect 32401 22383 32459 22389
rect 32766 22380 32772 22392
rect 32824 22380 32830 22432
rect 33502 22420 33508 22432
rect 33463 22392 33508 22420
rect 33502 22380 33508 22392
rect 33560 22380 33566 22432
rect 33689 22423 33747 22429
rect 33689 22389 33701 22423
rect 33735 22420 33747 22423
rect 34698 22420 34704 22432
rect 33735 22392 34704 22420
rect 33735 22389 33747 22392
rect 33689 22383 33747 22389
rect 34698 22380 34704 22392
rect 34756 22380 34762 22432
rect 38013 22423 38071 22429
rect 38013 22389 38025 22423
rect 38059 22420 38071 22423
rect 38102 22420 38108 22432
rect 38059 22392 38108 22420
rect 38059 22389 38071 22392
rect 38013 22383 38071 22389
rect 38102 22380 38108 22392
rect 38160 22380 38166 22432
rect 1104 22330 44896 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 44896 22330
rect 1104 22256 44896 22278
rect 1946 22176 1952 22228
rect 2004 22216 2010 22228
rect 2041 22219 2099 22225
rect 2041 22216 2053 22219
rect 2004 22188 2053 22216
rect 2004 22176 2010 22188
rect 2041 22185 2053 22188
rect 2087 22185 2099 22219
rect 2041 22179 2099 22185
rect 6178 22176 6184 22228
rect 6236 22216 6242 22228
rect 6236 22188 33916 22216
rect 6236 22176 6242 22188
rect 25866 22148 25872 22160
rect 25779 22120 25872 22148
rect 25866 22108 25872 22120
rect 25924 22148 25930 22160
rect 26881 22151 26939 22157
rect 26881 22148 26893 22151
rect 25924 22120 26893 22148
rect 25924 22108 25930 22120
rect 26881 22117 26893 22120
rect 26927 22117 26939 22151
rect 26881 22111 26939 22117
rect 28074 22108 28080 22160
rect 28132 22148 28138 22160
rect 30285 22151 30343 22157
rect 28132 22120 28994 22148
rect 28132 22108 28138 22120
rect 2866 22080 2872 22092
rect 2827 22052 2872 22080
rect 2866 22040 2872 22052
rect 2924 22040 2930 22092
rect 3142 22040 3148 22092
rect 3200 22080 3206 22092
rect 6086 22080 6092 22092
rect 3200 22052 6092 22080
rect 3200 22040 3206 22052
rect 6086 22040 6092 22052
rect 6144 22080 6150 22092
rect 6457 22083 6515 22089
rect 6457 22080 6469 22083
rect 6144 22052 6469 22080
rect 6144 22040 6150 22052
rect 6457 22049 6469 22052
rect 6503 22049 6515 22083
rect 6457 22043 6515 22049
rect 16298 22040 16304 22092
rect 16356 22080 16362 22092
rect 18138 22080 18144 22092
rect 16356 22052 18144 22080
rect 16356 22040 16362 22052
rect 18138 22040 18144 22052
rect 18196 22040 18202 22092
rect 19334 22080 19340 22092
rect 19295 22052 19340 22080
rect 19334 22040 19340 22052
rect 19392 22040 19398 22092
rect 25958 22080 25964 22092
rect 25919 22052 25964 22080
rect 25958 22040 25964 22052
rect 26016 22040 26022 22092
rect 26789 22083 26847 22089
rect 26789 22049 26801 22083
rect 26835 22080 26847 22083
rect 27430 22080 27436 22092
rect 26835 22052 27436 22080
rect 26835 22049 26847 22052
rect 26789 22043 26847 22049
rect 27430 22040 27436 22052
rect 27488 22080 27494 22092
rect 27617 22083 27675 22089
rect 27617 22080 27629 22083
rect 27488 22052 27629 22080
rect 27488 22040 27494 22052
rect 27617 22049 27629 22052
rect 27663 22049 27675 22083
rect 28966 22080 28994 22120
rect 30285 22117 30297 22151
rect 30331 22148 30343 22151
rect 30374 22148 30380 22160
rect 30331 22120 30380 22148
rect 30331 22117 30343 22120
rect 30285 22111 30343 22117
rect 30009 22083 30067 22089
rect 30009 22080 30021 22083
rect 28966 22052 30021 22080
rect 27617 22043 27675 22049
rect 30009 22049 30021 22052
rect 30055 22080 30067 22083
rect 30190 22080 30196 22092
rect 30055 22052 30196 22080
rect 30055 22049 30067 22052
rect 30009 22043 30067 22049
rect 30190 22040 30196 22052
rect 30248 22040 30254 22092
rect 2961 22015 3019 22021
rect 2961 21981 2973 22015
rect 3007 22012 3019 22015
rect 3970 22012 3976 22024
rect 3007 21984 3976 22012
rect 3007 21981 3019 21984
rect 2961 21975 3019 21981
rect 3970 21972 3976 21984
rect 4028 22012 4034 22024
rect 6178 22012 6184 22024
rect 4028 21984 6184 22012
rect 4028 21972 4034 21984
rect 6178 21972 6184 21984
rect 6236 21972 6242 22024
rect 6273 22015 6331 22021
rect 6273 21981 6285 22015
rect 6319 22012 6331 22015
rect 6362 22012 6368 22024
rect 6319 21984 6368 22012
rect 6319 21981 6331 21984
rect 6273 21975 6331 21981
rect 6362 21972 6368 21984
rect 6420 21972 6426 22024
rect 15286 21972 15292 22024
rect 15344 22012 15350 22024
rect 16025 22015 16083 22021
rect 16025 22012 16037 22015
rect 15344 21984 16037 22012
rect 15344 21972 15350 21984
rect 16025 21981 16037 21984
rect 16071 21981 16083 22015
rect 16025 21975 16083 21981
rect 15746 21944 15752 21956
rect 15707 21916 15752 21944
rect 15746 21904 15752 21916
rect 15804 21904 15810 21956
rect 16040 21944 16068 21975
rect 16666 21972 16672 22024
rect 16724 22012 16730 22024
rect 17497 22015 17555 22021
rect 17497 22012 17509 22015
rect 16724 21984 17509 22012
rect 16724 21972 16730 21984
rect 17497 21981 17509 21984
rect 17543 21981 17555 22015
rect 17497 21975 17555 21981
rect 17773 22015 17831 22021
rect 17773 21981 17785 22015
rect 17819 21981 17831 22015
rect 17773 21975 17831 21981
rect 19245 22015 19303 22021
rect 19245 21981 19257 22015
rect 19291 21981 19303 22015
rect 19245 21975 19303 21981
rect 19429 22015 19487 22021
rect 19429 21981 19441 22015
rect 19475 22012 19487 22015
rect 19978 22012 19984 22024
rect 19475 21984 19984 22012
rect 19475 21981 19487 21984
rect 19429 21975 19487 21981
rect 17788 21944 17816 21975
rect 18322 21944 18328 21956
rect 16040 21916 18328 21944
rect 18322 21904 18328 21916
rect 18380 21944 18386 21956
rect 18966 21944 18972 21956
rect 18380 21916 18972 21944
rect 18380 21904 18386 21916
rect 18966 21904 18972 21916
rect 19024 21944 19030 21956
rect 19260 21944 19288 21975
rect 19978 21972 19984 21984
rect 20036 21972 20042 22024
rect 20073 22015 20131 22021
rect 20073 21981 20085 22015
rect 20119 21981 20131 22015
rect 20254 22012 20260 22024
rect 20215 21984 20260 22012
rect 20073 21975 20131 21981
rect 19024 21916 19288 21944
rect 19024 21904 19030 21916
rect 19334 21904 19340 21956
rect 19392 21944 19398 21956
rect 20088 21944 20116 21975
rect 20254 21972 20260 21984
rect 20312 21972 20318 22024
rect 20898 22012 20904 22024
rect 20859 21984 20904 22012
rect 20898 21972 20904 21984
rect 20956 21972 20962 22024
rect 21450 21972 21456 22024
rect 21508 22012 21514 22024
rect 21545 22015 21603 22021
rect 21545 22012 21557 22015
rect 21508 21984 21557 22012
rect 21508 21972 21514 21984
rect 21545 21981 21557 21984
rect 21591 21981 21603 22015
rect 21545 21975 21603 21981
rect 25777 22015 25835 22021
rect 25777 21981 25789 22015
rect 25823 22012 25835 22015
rect 26326 22012 26332 22024
rect 25823 21984 26332 22012
rect 25823 21981 25835 21984
rect 25777 21975 25835 21981
rect 26326 21972 26332 21984
rect 26384 21972 26390 22024
rect 26697 22015 26755 22021
rect 26697 22012 26709 22015
rect 26436 21984 26709 22012
rect 26436 21956 26464 21984
rect 26697 21981 26709 21984
rect 26743 21981 26755 22015
rect 26970 22012 26976 22024
rect 26931 21984 26976 22012
rect 26697 21975 26755 21981
rect 21790 21947 21848 21953
rect 21790 21944 21802 21947
rect 19392 21916 20116 21944
rect 21100 21916 21802 21944
rect 19392 21904 19398 21916
rect 14734 21836 14740 21888
rect 14792 21876 14798 21888
rect 15847 21879 15905 21885
rect 15847 21876 15859 21879
rect 14792 21848 15859 21876
rect 14792 21836 14798 21848
rect 15847 21845 15859 21848
rect 15893 21845 15905 21879
rect 15847 21839 15905 21845
rect 15933 21879 15991 21885
rect 15933 21845 15945 21879
rect 15979 21876 15991 21879
rect 16390 21876 16396 21888
rect 15979 21848 16396 21876
rect 15979 21845 15991 21848
rect 15933 21839 15991 21845
rect 16390 21836 16396 21848
rect 16448 21836 16454 21888
rect 19242 21836 19248 21888
rect 19300 21876 19306 21888
rect 21100 21885 21128 21916
rect 21790 21913 21802 21916
rect 21836 21913 21848 21947
rect 21790 21907 21848 21913
rect 26145 21947 26203 21953
rect 26145 21913 26157 21947
rect 26191 21944 26203 21947
rect 26418 21944 26424 21956
rect 26191 21916 26424 21944
rect 26191 21913 26203 21916
rect 26145 21907 26203 21913
rect 26418 21904 26424 21916
rect 26476 21904 26482 21956
rect 26712 21944 26740 21975
rect 26970 21972 26976 21984
rect 27028 22012 27034 22024
rect 27338 22012 27344 22024
rect 27028 21984 27344 22012
rect 27028 21972 27034 21984
rect 27338 21972 27344 21984
rect 27396 21972 27402 22024
rect 27893 22015 27951 22021
rect 27893 21981 27905 22015
rect 27939 21981 27951 22015
rect 27893 21975 27951 21981
rect 27522 21944 27528 21956
rect 26712 21916 27528 21944
rect 27522 21904 27528 21916
rect 27580 21904 27586 21956
rect 27908 21944 27936 21975
rect 30300 21944 30328 22111
rect 30374 22108 30380 22120
rect 30432 22108 30438 22160
rect 30469 22151 30527 22157
rect 30469 22117 30481 22151
rect 30515 22148 30527 22151
rect 31018 22148 31024 22160
rect 30515 22120 31024 22148
rect 30515 22117 30527 22120
rect 30469 22111 30527 22117
rect 31018 22108 31024 22120
rect 31076 22108 31082 22160
rect 33778 22148 33784 22160
rect 33739 22120 33784 22148
rect 33778 22108 33784 22120
rect 33836 22108 33842 22160
rect 33888 22148 33916 22188
rect 33962 22176 33968 22228
rect 34020 22216 34026 22228
rect 41690 22216 41696 22228
rect 34020 22188 34065 22216
rect 34164 22188 41696 22216
rect 34020 22176 34026 22188
rect 34164 22148 34192 22188
rect 41690 22176 41696 22188
rect 41748 22176 41754 22228
rect 41785 22219 41843 22225
rect 41785 22185 41797 22219
rect 41831 22216 41843 22219
rect 42426 22216 42432 22228
rect 41831 22188 42432 22216
rect 41831 22185 41843 22188
rect 41785 22179 41843 22185
rect 42426 22176 42432 22188
rect 42484 22176 42490 22228
rect 33888 22120 34192 22148
rect 38013 22151 38071 22157
rect 38013 22117 38025 22151
rect 38059 22148 38071 22151
rect 38746 22148 38752 22160
rect 38059 22120 38752 22148
rect 38059 22117 38071 22120
rect 38013 22111 38071 22117
rect 38746 22108 38752 22120
rect 38804 22108 38810 22160
rect 31938 22080 31944 22092
rect 31899 22052 31944 22080
rect 31938 22040 31944 22052
rect 31996 22040 32002 22092
rect 42334 22080 42340 22092
rect 32416 22052 40540 22080
rect 42295 22052 42340 22080
rect 32416 22012 32444 22052
rect 27908 21916 30328 21944
rect 30392 21984 32444 22012
rect 20165 21879 20223 21885
rect 20165 21876 20177 21879
rect 19300 21848 20177 21876
rect 19300 21836 19306 21848
rect 20165 21845 20177 21848
rect 20211 21845 20223 21879
rect 20165 21839 20223 21845
rect 21085 21879 21143 21885
rect 21085 21845 21097 21879
rect 21131 21845 21143 21879
rect 22922 21876 22928 21888
rect 22883 21848 22928 21876
rect 21085 21839 21143 21845
rect 22922 21836 22928 21848
rect 22980 21836 22986 21888
rect 26050 21876 26056 21888
rect 26011 21848 26056 21876
rect 26050 21836 26056 21848
rect 26108 21836 26114 21888
rect 27154 21876 27160 21888
rect 27115 21848 27160 21876
rect 27154 21836 27160 21848
rect 27212 21836 27218 21888
rect 27338 21836 27344 21888
rect 27396 21876 27402 21888
rect 27908 21876 27936 21916
rect 27396 21848 27936 21876
rect 27396 21836 27402 21848
rect 29086 21836 29092 21888
rect 29144 21876 29150 21888
rect 30392 21876 30420 21984
rect 32490 21972 32496 22024
rect 32548 22012 32554 22024
rect 32766 22012 32772 22024
rect 32548 21984 32593 22012
rect 32727 21984 32772 22012
rect 32548 21972 32554 21984
rect 32766 21972 32772 21984
rect 32824 21972 32830 22024
rect 34698 22012 34704 22024
rect 34659 21984 34704 22012
rect 34698 21972 34704 21984
rect 34756 21972 34762 22024
rect 35526 21972 35532 22024
rect 35584 22012 35590 22024
rect 35621 22015 35679 22021
rect 35621 22012 35633 22015
rect 35584 21984 35633 22012
rect 35584 21972 35590 21984
rect 35621 21981 35633 21984
rect 35667 21981 35679 22015
rect 35802 22012 35808 22024
rect 35763 21984 35808 22012
rect 35621 21975 35679 21981
rect 35802 21972 35808 21984
rect 35860 21972 35866 22024
rect 35986 22012 35992 22024
rect 35947 21984 35992 22012
rect 35986 21972 35992 21984
rect 36044 21972 36050 22024
rect 37642 22012 37648 22024
rect 37603 21984 37648 22012
rect 37642 21972 37648 21984
rect 37700 21972 37706 22024
rect 38838 22012 38844 22024
rect 38799 21984 38844 22012
rect 38838 21972 38844 21984
rect 38896 21972 38902 22024
rect 39114 22012 39120 22024
rect 39075 21984 39120 22012
rect 39114 21972 39120 21984
rect 39172 21972 39178 22024
rect 40402 22012 40408 22024
rect 40363 21984 40408 22012
rect 40402 21972 40408 21984
rect 40460 21972 40466 22024
rect 40512 22012 40540 22052
rect 42334 22040 42340 22052
rect 42392 22040 42398 22092
rect 42518 22080 42524 22092
rect 42479 22052 42524 22080
rect 42518 22040 42524 22052
rect 42576 22040 42582 22092
rect 42610 22040 42616 22092
rect 42668 22080 42674 22092
rect 42797 22083 42855 22089
rect 42797 22080 42809 22083
rect 42668 22052 42809 22080
rect 42668 22040 42674 22052
rect 42797 22049 42809 22052
rect 42843 22049 42855 22083
rect 42797 22043 42855 22049
rect 41414 22012 41420 22024
rect 40512 21984 41420 22012
rect 41414 21972 41420 21984
rect 41472 21972 41478 22024
rect 31386 21904 31392 21956
rect 31444 21944 31450 21956
rect 31754 21944 31760 21956
rect 31444 21916 31760 21944
rect 31444 21904 31450 21916
rect 31754 21904 31760 21916
rect 31812 21944 31818 21956
rect 31812 21916 31905 21944
rect 31812 21904 31818 21916
rect 31938 21904 31944 21956
rect 31996 21944 32002 21956
rect 32585 21947 32643 21953
rect 32585 21944 32597 21947
rect 31996 21916 32597 21944
rect 31996 21904 32002 21916
rect 32585 21913 32597 21916
rect 32631 21913 32643 21947
rect 32585 21907 32643 21913
rect 34149 21947 34207 21953
rect 34149 21913 34161 21947
rect 34195 21944 34207 21947
rect 34330 21944 34336 21956
rect 34195 21916 34336 21944
rect 34195 21913 34207 21916
rect 34149 21907 34207 21913
rect 34330 21904 34336 21916
rect 34388 21944 34394 21956
rect 35897 21947 35955 21953
rect 35897 21944 35909 21947
rect 34388 21916 35909 21944
rect 34388 21904 34394 21916
rect 35897 21913 35909 21916
rect 35943 21913 35955 21947
rect 35897 21907 35955 21913
rect 38746 21904 38752 21956
rect 38804 21944 38810 21956
rect 38933 21947 38991 21953
rect 38933 21944 38945 21947
rect 38804 21916 38945 21944
rect 38804 21904 38810 21916
rect 38933 21913 38945 21916
rect 38979 21913 38991 21947
rect 38933 21907 38991 21913
rect 40126 21904 40132 21956
rect 40184 21944 40190 21956
rect 40650 21947 40708 21953
rect 40650 21944 40662 21947
rect 40184 21916 40662 21944
rect 40184 21904 40190 21916
rect 40650 21913 40662 21916
rect 40696 21913 40708 21947
rect 40650 21907 40708 21913
rect 29144 21848 30420 21876
rect 29144 21836 29150 21848
rect 30558 21836 30564 21888
rect 30616 21876 30622 21888
rect 31297 21879 31355 21885
rect 31297 21876 31309 21879
rect 30616 21848 31309 21876
rect 30616 21836 30622 21848
rect 31297 21845 31309 21848
rect 31343 21845 31355 21879
rect 31662 21876 31668 21888
rect 31623 21848 31668 21876
rect 31297 21839 31355 21845
rect 31662 21836 31668 21848
rect 31720 21836 31726 21888
rect 32674 21885 32680 21888
rect 32670 21876 32680 21885
rect 32635 21848 32680 21876
rect 32670 21839 32680 21848
rect 32674 21836 32680 21839
rect 32732 21836 32738 21888
rect 33949 21879 34007 21885
rect 33949 21845 33961 21879
rect 33995 21876 34007 21879
rect 34422 21876 34428 21888
rect 33995 21848 34428 21876
rect 33995 21845 34007 21848
rect 33949 21839 34007 21845
rect 34422 21836 34428 21848
rect 34480 21836 34486 21888
rect 34790 21836 34796 21888
rect 34848 21876 34854 21888
rect 34885 21879 34943 21885
rect 34885 21876 34897 21879
rect 34848 21848 34897 21876
rect 34848 21836 34854 21848
rect 34885 21845 34897 21848
rect 34931 21845 34943 21879
rect 36170 21876 36176 21888
rect 36131 21848 36176 21876
rect 34885 21839 34943 21845
rect 36170 21836 36176 21848
rect 36228 21836 36234 21888
rect 38105 21879 38163 21885
rect 38105 21845 38117 21879
rect 38151 21876 38163 21879
rect 38194 21876 38200 21888
rect 38151 21848 38200 21876
rect 38151 21845 38163 21848
rect 38105 21839 38163 21845
rect 38194 21836 38200 21848
rect 38252 21836 38258 21888
rect 39301 21879 39359 21885
rect 39301 21845 39313 21879
rect 39347 21876 39359 21879
rect 39758 21876 39764 21888
rect 39347 21848 39764 21876
rect 39347 21845 39359 21848
rect 39301 21839 39359 21845
rect 39758 21836 39764 21848
rect 39816 21836 39822 21888
rect 1104 21786 44896 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 44896 21786
rect 1104 21712 44896 21734
rect 7926 21632 7932 21684
rect 7984 21672 7990 21684
rect 8021 21675 8079 21681
rect 8021 21672 8033 21675
rect 7984 21644 8033 21672
rect 7984 21632 7990 21644
rect 8021 21641 8033 21644
rect 8067 21672 8079 21675
rect 8202 21672 8208 21684
rect 8067 21644 8208 21672
rect 8067 21641 8079 21644
rect 8021 21635 8079 21641
rect 8202 21632 8208 21644
rect 8260 21632 8266 21684
rect 17770 21632 17776 21684
rect 17828 21672 17834 21684
rect 17828 21644 19380 21672
rect 17828 21632 17834 21644
rect 6362 21604 6368 21616
rect 5736 21576 6368 21604
rect 5534 21496 5540 21548
rect 5592 21536 5598 21548
rect 5736 21545 5764 21576
rect 6362 21564 6368 21576
rect 6420 21604 6426 21616
rect 6733 21607 6791 21613
rect 6733 21604 6745 21607
rect 6420 21576 6745 21604
rect 6420 21564 6426 21576
rect 6733 21573 6745 21576
rect 6779 21573 6791 21607
rect 18138 21604 18144 21616
rect 18099 21576 18144 21604
rect 6733 21567 6791 21573
rect 18138 21564 18144 21576
rect 18196 21564 18202 21616
rect 5721 21539 5779 21545
rect 5721 21536 5733 21539
rect 5592 21508 5733 21536
rect 5592 21496 5598 21508
rect 5721 21505 5733 21508
rect 5767 21505 5779 21539
rect 5721 21499 5779 21505
rect 15004 21539 15062 21545
rect 15004 21505 15016 21539
rect 15050 21536 15062 21539
rect 17865 21539 17923 21545
rect 17865 21536 17877 21539
rect 15050 21508 17877 21536
rect 15050 21505 15062 21508
rect 15004 21499 15062 21505
rect 17865 21505 17877 21508
rect 17911 21505 17923 21539
rect 17865 21499 17923 21505
rect 18049 21539 18107 21545
rect 18049 21505 18061 21539
rect 18095 21505 18107 21539
rect 18230 21536 18236 21548
rect 18191 21508 18236 21536
rect 18049 21499 18107 21505
rect 5166 21428 5172 21480
rect 5224 21468 5230 21480
rect 5445 21471 5503 21477
rect 5445 21468 5457 21471
rect 5224 21440 5457 21468
rect 5224 21428 5230 21440
rect 5445 21437 5457 21440
rect 5491 21468 5503 21471
rect 6546 21468 6552 21480
rect 5491 21440 6552 21468
rect 5491 21437 5503 21440
rect 5445 21431 5503 21437
rect 6546 21428 6552 21440
rect 6604 21428 6610 21480
rect 14737 21471 14795 21477
rect 14737 21437 14749 21471
rect 14783 21437 14795 21471
rect 14737 21431 14795 21437
rect 14752 21332 14780 21431
rect 18064 21400 18092 21499
rect 18230 21496 18236 21508
rect 18288 21496 18294 21548
rect 18524 21545 18552 21644
rect 19242 21604 19248 21616
rect 19203 21576 19248 21604
rect 19242 21564 19248 21576
rect 19300 21564 19306 21616
rect 18351 21539 18409 21545
rect 18351 21505 18363 21539
rect 18397 21536 18409 21539
rect 18509 21539 18567 21545
rect 18397 21505 18414 21536
rect 18351 21499 18414 21505
rect 18509 21505 18521 21539
rect 18555 21505 18567 21539
rect 18966 21536 18972 21548
rect 18927 21508 18972 21536
rect 18509 21499 18567 21505
rect 18386 21468 18414 21499
rect 18966 21496 18972 21508
rect 19024 21496 19030 21548
rect 19058 21496 19064 21548
rect 19116 21536 19122 21548
rect 19352 21536 19380 21644
rect 19426 21632 19432 21684
rect 19484 21672 19490 21684
rect 19797 21675 19855 21681
rect 19797 21672 19809 21675
rect 19484 21644 19809 21672
rect 19484 21632 19490 21644
rect 19797 21641 19809 21644
rect 19843 21641 19855 21675
rect 19797 21635 19855 21641
rect 25685 21675 25743 21681
rect 25685 21641 25697 21675
rect 25731 21672 25743 21675
rect 26326 21672 26332 21684
rect 25731 21644 26332 21672
rect 25731 21641 25743 21644
rect 25685 21635 25743 21641
rect 26326 21632 26332 21644
rect 26384 21672 26390 21684
rect 26970 21672 26976 21684
rect 26384 21644 26976 21672
rect 26384 21632 26390 21644
rect 26970 21632 26976 21644
rect 27028 21632 27034 21684
rect 27246 21672 27252 21684
rect 27207 21644 27252 21672
rect 27246 21632 27252 21644
rect 27304 21632 27310 21684
rect 30926 21672 30932 21684
rect 28552 21644 30932 21672
rect 19889 21607 19947 21613
rect 19889 21573 19901 21607
rect 19935 21604 19947 21607
rect 22278 21604 22284 21616
rect 19935 21576 22284 21604
rect 19935 21573 19947 21576
rect 19889 21567 19947 21573
rect 22278 21564 22284 21576
rect 22336 21604 22342 21616
rect 22462 21604 22468 21616
rect 22336 21576 22468 21604
rect 22336 21564 22342 21576
rect 22462 21564 22468 21576
rect 22520 21564 22526 21616
rect 28074 21604 28080 21616
rect 27448 21576 28080 21604
rect 20070 21536 20076 21548
rect 19116 21508 19161 21536
rect 19352 21508 20076 21536
rect 19116 21496 19122 21508
rect 20070 21496 20076 21508
rect 20128 21536 20134 21548
rect 20254 21536 20260 21548
rect 20128 21508 20260 21536
rect 20128 21496 20134 21508
rect 20254 21496 20260 21508
rect 20312 21496 20318 21548
rect 20806 21496 20812 21548
rect 20864 21536 20870 21548
rect 20901 21539 20959 21545
rect 20901 21536 20913 21539
rect 20864 21508 20913 21536
rect 20864 21496 20870 21508
rect 20901 21505 20913 21508
rect 20947 21505 20959 21539
rect 20901 21499 20959 21505
rect 21085 21539 21143 21545
rect 21085 21505 21097 21539
rect 21131 21536 21143 21539
rect 22005 21539 22063 21545
rect 22005 21536 22017 21539
rect 21131 21508 22017 21536
rect 21131 21505 21143 21508
rect 21085 21499 21143 21505
rect 22005 21505 22017 21508
rect 22051 21505 22063 21539
rect 22005 21499 22063 21505
rect 18386 21440 19380 21468
rect 19245 21403 19303 21409
rect 19245 21400 19257 21403
rect 18064 21372 19257 21400
rect 19245 21369 19257 21372
rect 19291 21369 19303 21403
rect 19352 21400 19380 21440
rect 19518 21428 19524 21480
rect 19576 21468 19582 21480
rect 20622 21468 20628 21480
rect 19576 21440 20628 21468
rect 19576 21428 19582 21440
rect 20622 21428 20628 21440
rect 20680 21468 20686 21480
rect 20717 21471 20775 21477
rect 20717 21468 20729 21471
rect 20680 21440 20729 21468
rect 20680 21428 20686 21440
rect 20717 21437 20729 21440
rect 20763 21437 20775 21471
rect 20717 21431 20775 21437
rect 20346 21400 20352 21412
rect 19352 21372 20352 21400
rect 19245 21363 19303 21369
rect 20346 21360 20352 21372
rect 20404 21360 20410 21412
rect 20916 21400 20944 21499
rect 22370 21496 22376 21548
rect 22428 21536 22434 21548
rect 24578 21545 24584 21548
rect 22721 21539 22779 21545
rect 22721 21536 22733 21539
rect 22428 21508 22733 21536
rect 22428 21496 22434 21508
rect 22721 21505 22733 21508
rect 22767 21505 22779 21539
rect 22721 21499 22779 21505
rect 24572 21499 24584 21545
rect 24636 21536 24642 21548
rect 27448 21545 27476 21576
rect 28074 21564 28080 21576
rect 28132 21564 28138 21616
rect 28552 21545 28580 21644
rect 30926 21632 30932 21644
rect 30984 21632 30990 21684
rect 32490 21672 32496 21684
rect 31036 21644 32496 21672
rect 29457 21607 29515 21613
rect 29457 21604 29469 21607
rect 28920 21576 29469 21604
rect 27433 21539 27491 21545
rect 24636 21508 24672 21536
rect 24578 21496 24584 21499
rect 24636 21496 24642 21508
rect 27433 21505 27445 21539
rect 27479 21505 27491 21539
rect 27433 21499 27491 21505
rect 27709 21539 27767 21545
rect 27709 21505 27721 21539
rect 27755 21505 27767 21539
rect 27709 21499 27767 21505
rect 28537 21539 28595 21545
rect 28537 21505 28549 21539
rect 28583 21505 28595 21539
rect 28537 21499 28595 21505
rect 21450 21428 21456 21480
rect 21508 21468 21514 21480
rect 22465 21471 22523 21477
rect 22465 21468 22477 21471
rect 21508 21440 22477 21468
rect 21508 21428 21514 21440
rect 22465 21437 22477 21440
rect 22511 21437 22523 21471
rect 22465 21431 22523 21437
rect 23658 21428 23664 21480
rect 23716 21468 23722 21480
rect 24302 21468 24308 21480
rect 23716 21440 24308 21468
rect 23716 21428 23722 21440
rect 24302 21428 24308 21440
rect 24360 21428 24366 21480
rect 25958 21428 25964 21480
rect 26016 21468 26022 21480
rect 27338 21468 27344 21480
rect 26016 21440 27344 21468
rect 26016 21428 26022 21440
rect 27338 21428 27344 21440
rect 27396 21468 27402 21480
rect 27525 21471 27583 21477
rect 27525 21468 27537 21471
rect 27396 21440 27537 21468
rect 27396 21428 27402 21440
rect 27525 21437 27537 21440
rect 27571 21437 27583 21471
rect 27525 21431 27583 21437
rect 22094 21400 22100 21412
rect 20916 21372 22100 21400
rect 22094 21360 22100 21372
rect 22152 21360 22158 21412
rect 27724 21400 27752 21499
rect 28552 21468 28580 21499
rect 27540 21372 27752 21400
rect 27816 21440 28580 21468
rect 27540 21344 27568 21372
rect 15470 21332 15476 21344
rect 14752 21304 15476 21332
rect 15470 21292 15476 21304
rect 15528 21292 15534 21344
rect 16117 21335 16175 21341
rect 16117 21301 16129 21335
rect 16163 21332 16175 21335
rect 17494 21332 17500 21344
rect 16163 21304 17500 21332
rect 16163 21301 16175 21304
rect 16117 21295 16175 21301
rect 17494 21292 17500 21304
rect 17552 21292 17558 21344
rect 18230 21292 18236 21344
rect 18288 21332 18294 21344
rect 20438 21332 20444 21344
rect 18288 21304 20444 21332
rect 18288 21292 18294 21304
rect 20438 21292 20444 21304
rect 20496 21292 20502 21344
rect 21726 21292 21732 21344
rect 21784 21332 21790 21344
rect 21821 21335 21879 21341
rect 21821 21332 21833 21335
rect 21784 21304 21833 21332
rect 21784 21292 21790 21304
rect 21821 21301 21833 21304
rect 21867 21301 21879 21335
rect 21821 21295 21879 21301
rect 23845 21335 23903 21341
rect 23845 21301 23857 21335
rect 23891 21332 23903 21335
rect 25866 21332 25872 21344
rect 23891 21304 25872 21332
rect 23891 21301 23903 21304
rect 23845 21295 23903 21301
rect 25866 21292 25872 21304
rect 25924 21292 25930 21344
rect 27522 21292 27528 21344
rect 27580 21292 27586 21344
rect 27709 21335 27767 21341
rect 27709 21301 27721 21335
rect 27755 21332 27767 21335
rect 27816 21332 27844 21440
rect 28626 21428 28632 21480
rect 28684 21468 28690 21480
rect 28920 21477 28948 21576
rect 29457 21573 29469 21576
rect 29503 21604 29515 21607
rect 29822 21604 29828 21616
rect 29503 21576 29828 21604
rect 29503 21573 29515 21576
rect 29457 21567 29515 21573
rect 29822 21564 29828 21576
rect 29880 21564 29886 21616
rect 30742 21604 30748 21616
rect 30392 21576 30748 21604
rect 29362 21496 29368 21548
rect 29420 21536 29426 21548
rect 30392 21536 30420 21576
rect 30742 21564 30748 21576
rect 30800 21564 30806 21616
rect 30834 21564 30840 21616
rect 30892 21604 30898 21616
rect 31036 21604 31064 21644
rect 32490 21632 32496 21644
rect 32548 21632 32554 21684
rect 33689 21675 33747 21681
rect 33689 21641 33701 21675
rect 33735 21672 33747 21675
rect 34330 21672 34336 21684
rect 33735 21644 34336 21672
rect 33735 21641 33747 21644
rect 33689 21635 33747 21641
rect 34330 21632 34336 21644
rect 34388 21632 34394 21684
rect 36078 21672 36084 21684
rect 34440 21644 36084 21672
rect 30892 21576 31064 21604
rect 30892 21564 30898 21576
rect 31662 21564 31668 21616
rect 31720 21604 31726 21616
rect 34440 21604 34468 21644
rect 36078 21632 36084 21644
rect 36136 21632 36142 21684
rect 38197 21675 38255 21681
rect 38197 21641 38209 21675
rect 38243 21672 38255 21675
rect 39114 21672 39120 21684
rect 38243 21644 39120 21672
rect 38243 21641 38255 21644
rect 38197 21635 38255 21641
rect 39114 21632 39120 21644
rect 39172 21632 39178 21684
rect 40126 21672 40132 21684
rect 40087 21644 40132 21672
rect 40126 21632 40132 21644
rect 40184 21632 40190 21684
rect 34790 21604 34796 21616
rect 34848 21613 34854 21616
rect 31720 21576 34468 21604
rect 34760 21576 34796 21604
rect 31720 21564 31726 21576
rect 34790 21564 34796 21576
rect 34848 21567 34860 21613
rect 38749 21607 38807 21613
rect 38749 21604 38761 21607
rect 38212 21576 38761 21604
rect 34848 21564 34854 21567
rect 38212 21548 38240 21576
rect 38749 21573 38761 21576
rect 38795 21573 38807 21607
rect 38749 21567 38807 21573
rect 30558 21536 30564 21548
rect 29420 21508 30420 21536
rect 30519 21508 30564 21536
rect 29420 21496 29426 21508
rect 30558 21496 30564 21508
rect 30616 21496 30622 21548
rect 31021 21539 31079 21545
rect 31021 21505 31033 21539
rect 31067 21536 31079 21539
rect 31938 21536 31944 21548
rect 31067 21508 31944 21536
rect 31067 21505 31079 21508
rect 31021 21499 31079 21505
rect 31938 21496 31944 21508
rect 31996 21496 32002 21548
rect 36170 21496 36176 21548
rect 36228 21536 36234 21548
rect 36357 21539 36415 21545
rect 36357 21536 36369 21539
rect 36228 21508 36369 21536
rect 36228 21496 36234 21508
rect 36357 21505 36369 21508
rect 36403 21505 36415 21539
rect 36357 21499 36415 21505
rect 38105 21539 38163 21545
rect 38105 21505 38117 21539
rect 38151 21536 38163 21539
rect 38194 21536 38200 21548
rect 38151 21508 38200 21536
rect 38151 21505 38163 21508
rect 38105 21499 38163 21505
rect 38194 21496 38200 21508
rect 38252 21496 38258 21548
rect 38289 21539 38347 21545
rect 38289 21505 38301 21539
rect 38335 21505 38347 21539
rect 38289 21499 38347 21505
rect 39945 21539 40003 21545
rect 39945 21505 39957 21539
rect 39991 21505 40003 21539
rect 39945 21499 40003 21505
rect 28905 21471 28963 21477
rect 28684 21440 28856 21468
rect 28684 21428 28690 21440
rect 28828 21400 28856 21440
rect 28905 21437 28917 21471
rect 28951 21437 28963 21471
rect 28905 21431 28963 21437
rect 30190 21428 30196 21480
rect 30248 21468 30254 21480
rect 30837 21471 30895 21477
rect 30837 21468 30849 21471
rect 30248 21440 30849 21468
rect 30248 21428 30254 21440
rect 30837 21437 30849 21440
rect 30883 21468 30895 21471
rect 32306 21468 32312 21480
rect 30883 21440 32312 21468
rect 30883 21437 30895 21440
rect 30837 21431 30895 21437
rect 32306 21428 32312 21440
rect 32364 21428 32370 21480
rect 35069 21471 35127 21477
rect 35069 21437 35081 21471
rect 35115 21468 35127 21471
rect 35342 21468 35348 21480
rect 35115 21440 35348 21468
rect 35115 21437 35127 21440
rect 35069 21431 35127 21437
rect 35342 21428 35348 21440
rect 35400 21428 35406 21480
rect 35894 21428 35900 21480
rect 35952 21468 35958 21480
rect 36265 21471 36323 21477
rect 36265 21468 36277 21471
rect 35952 21440 36277 21468
rect 35952 21428 35958 21440
rect 36265 21437 36277 21440
rect 36311 21437 36323 21471
rect 38304 21468 38332 21499
rect 38746 21468 38752 21480
rect 36265 21431 36323 21437
rect 36740 21440 38752 21468
rect 31570 21400 31576 21412
rect 28828 21372 31576 21400
rect 31570 21360 31576 21372
rect 31628 21360 31634 21412
rect 33042 21360 33048 21412
rect 33100 21400 33106 21412
rect 36740 21409 36768 21440
rect 38746 21428 38752 21440
rect 38804 21468 38810 21480
rect 39209 21471 39267 21477
rect 38804 21440 39068 21468
rect 38804 21428 38810 21440
rect 39040 21409 39068 21440
rect 39209 21437 39221 21471
rect 39255 21468 39267 21471
rect 39960 21468 39988 21499
rect 41690 21496 41696 21548
rect 41748 21536 41754 21548
rect 42429 21539 42487 21545
rect 42429 21536 42441 21539
rect 41748 21508 42441 21536
rect 41748 21496 41754 21508
rect 42429 21505 42441 21508
rect 42475 21505 42487 21539
rect 42429 21499 42487 21505
rect 39255 21440 39988 21468
rect 39255 21437 39267 21440
rect 39209 21431 39267 21437
rect 36725 21403 36783 21409
rect 33100 21372 33824 21400
rect 33100 21360 33106 21372
rect 27890 21332 27896 21344
rect 27755 21304 27896 21332
rect 27755 21301 27767 21304
rect 27709 21295 27767 21301
rect 27890 21292 27896 21304
rect 27948 21292 27954 21344
rect 29362 21292 29368 21344
rect 29420 21332 29426 21344
rect 29549 21335 29607 21341
rect 29549 21332 29561 21335
rect 29420 21304 29561 21332
rect 29420 21292 29426 21304
rect 29549 21301 29561 21304
rect 29595 21301 29607 21335
rect 29549 21295 29607 21301
rect 30374 21292 30380 21344
rect 30432 21332 30438 21344
rect 30699 21335 30757 21341
rect 30699 21332 30711 21335
rect 30432 21304 30711 21332
rect 30432 21292 30438 21304
rect 30699 21301 30711 21304
rect 30745 21332 30757 21335
rect 30834 21332 30840 21344
rect 30745 21304 30840 21332
rect 30745 21301 30757 21304
rect 30699 21295 30757 21301
rect 30834 21292 30840 21304
rect 30892 21292 30898 21344
rect 30926 21292 30932 21344
rect 30984 21332 30990 21344
rect 33796 21332 33824 21372
rect 36725 21369 36737 21403
rect 36771 21369 36783 21403
rect 36725 21363 36783 21369
rect 39025 21403 39083 21409
rect 39025 21369 39037 21403
rect 39071 21369 39083 21403
rect 39025 21363 39083 21369
rect 35434 21332 35440 21344
rect 30984 21304 31029 21332
rect 33796 21304 35440 21332
rect 30984 21292 30990 21304
rect 35434 21292 35440 21304
rect 35492 21292 35498 21344
rect 42058 21292 42064 21344
rect 42116 21332 42122 21344
rect 42521 21335 42579 21341
rect 42521 21332 42533 21335
rect 42116 21304 42533 21332
rect 42116 21292 42122 21304
rect 42521 21301 42533 21304
rect 42567 21301 42579 21335
rect 42521 21295 42579 21301
rect 42610 21292 42616 21344
rect 42668 21332 42674 21344
rect 43625 21335 43683 21341
rect 43625 21332 43637 21335
rect 42668 21304 43637 21332
rect 42668 21292 42674 21304
rect 43625 21301 43637 21304
rect 43671 21301 43683 21335
rect 43625 21295 43683 21301
rect 1104 21242 44896 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 44896 21242
rect 1104 21168 44896 21190
rect 5534 21128 5540 21140
rect 5495 21100 5540 21128
rect 5534 21088 5540 21100
rect 5592 21088 5598 21140
rect 23290 21128 23296 21140
rect 23251 21100 23296 21128
rect 23290 21088 23296 21100
rect 23348 21088 23354 21140
rect 24578 21128 24584 21140
rect 24539 21100 24584 21128
rect 24578 21088 24584 21100
rect 24636 21088 24642 21140
rect 26053 21131 26111 21137
rect 26053 21097 26065 21131
rect 26099 21097 26111 21131
rect 26234 21128 26240 21140
rect 26195 21100 26240 21128
rect 26053 21091 26111 21097
rect 22833 21063 22891 21069
rect 22833 21029 22845 21063
rect 22879 21060 22891 21063
rect 23753 21063 23811 21069
rect 22879 21032 23428 21060
rect 22879 21029 22891 21032
rect 22833 21023 22891 21029
rect 6822 20992 6828 21004
rect 6783 20964 6828 20992
rect 6822 20952 6828 20964
rect 6880 20952 6886 21004
rect 16298 20992 16304 21004
rect 15488 20964 16304 20992
rect 1670 20884 1676 20936
rect 1728 20924 1734 20936
rect 1765 20927 1823 20933
rect 1765 20924 1777 20927
rect 1728 20896 1777 20924
rect 1728 20884 1734 20896
rect 1765 20893 1777 20896
rect 1811 20893 1823 20927
rect 1765 20887 1823 20893
rect 3878 20884 3884 20936
rect 3936 20924 3942 20936
rect 5353 20927 5411 20933
rect 5353 20924 5365 20927
rect 3936 20896 5365 20924
rect 3936 20884 3942 20896
rect 5353 20893 5365 20896
rect 5399 20893 5411 20927
rect 5353 20887 5411 20893
rect 5368 20856 5396 20887
rect 5534 20884 5540 20936
rect 5592 20924 5598 20936
rect 6089 20927 6147 20933
rect 6089 20924 6101 20927
rect 5592 20896 6101 20924
rect 5592 20884 5598 20896
rect 6089 20893 6101 20896
rect 6135 20893 6147 20927
rect 11333 20927 11391 20933
rect 11333 20924 11345 20927
rect 6089 20887 6147 20893
rect 6886 20896 11345 20924
rect 6886 20856 6914 20896
rect 11333 20893 11345 20896
rect 11379 20893 11391 20927
rect 14550 20924 14556 20936
rect 14511 20896 14556 20924
rect 11333 20887 11391 20893
rect 14550 20884 14556 20896
rect 14608 20884 14614 20936
rect 14734 20924 14740 20936
rect 14695 20896 14740 20924
rect 14734 20884 14740 20896
rect 14792 20884 14798 20936
rect 15488 20933 15516 20964
rect 16298 20952 16304 20964
rect 16356 20952 16362 21004
rect 17494 20992 17500 21004
rect 17455 20964 17500 20992
rect 17494 20952 17500 20964
rect 17552 20952 17558 21004
rect 17770 20992 17776 21004
rect 17731 20964 17776 20992
rect 17770 20952 17776 20964
rect 17828 20952 17834 21004
rect 19426 20952 19432 21004
rect 19484 20992 19490 21004
rect 19613 20995 19671 21001
rect 19613 20992 19625 20995
rect 19484 20964 19625 20992
rect 19484 20952 19490 20964
rect 19613 20961 19625 20964
rect 19659 20961 19671 20995
rect 21450 20992 21456 21004
rect 21411 20964 21456 20992
rect 19613 20955 19671 20961
rect 21450 20952 21456 20964
rect 21508 20952 21514 21004
rect 23400 21001 23428 21032
rect 23753 21029 23765 21063
rect 23799 21029 23811 21063
rect 26068 21060 26096 21091
rect 26234 21088 26240 21100
rect 26292 21088 26298 21140
rect 27890 21128 27896 21140
rect 27851 21100 27896 21128
rect 27890 21088 27896 21100
rect 27948 21088 27954 21140
rect 28626 21128 28632 21140
rect 28587 21100 28632 21128
rect 28626 21088 28632 21100
rect 28684 21088 28690 21140
rect 30190 21128 30196 21140
rect 30151 21100 30196 21128
rect 30190 21088 30196 21100
rect 30248 21088 30254 21140
rect 31938 21128 31944 21140
rect 31899 21100 31944 21128
rect 31938 21088 31944 21100
rect 31996 21088 32002 21140
rect 33045 21131 33103 21137
rect 33045 21097 33057 21131
rect 33091 21128 33103 21131
rect 33134 21128 33140 21140
rect 33091 21100 33140 21128
rect 33091 21097 33103 21100
rect 33045 21091 33103 21097
rect 33134 21088 33140 21100
rect 33192 21128 33198 21140
rect 33192 21100 34100 21128
rect 33192 21088 33198 21100
rect 26142 21060 26148 21072
rect 26068 21032 26148 21060
rect 23753 21023 23811 21029
rect 23385 20995 23443 21001
rect 23385 20961 23397 20995
rect 23431 20961 23443 20995
rect 23768 20992 23796 21023
rect 26142 21020 26148 21032
rect 26200 21020 26206 21072
rect 27062 21020 27068 21072
rect 27120 21060 27126 21072
rect 27157 21063 27215 21069
rect 27157 21060 27169 21063
rect 27120 21032 27169 21060
rect 27120 21020 27126 21032
rect 27157 21029 27169 21032
rect 27203 21029 27215 21063
rect 27157 21023 27215 21029
rect 28736 21032 33916 21060
rect 25961 20995 26019 21001
rect 23768 20964 25912 20992
rect 23385 20955 23443 20961
rect 15381 20927 15439 20933
rect 15381 20893 15393 20927
rect 15427 20893 15439 20927
rect 15381 20887 15439 20893
rect 15473 20927 15531 20933
rect 15473 20893 15485 20927
rect 15519 20893 15531 20927
rect 15473 20887 15531 20893
rect 15841 20927 15899 20933
rect 15841 20893 15853 20927
rect 15887 20924 15899 20927
rect 15930 20924 15936 20936
rect 15887 20896 15936 20924
rect 15887 20893 15899 20896
rect 15841 20887 15899 20893
rect 5368 20828 6914 20856
rect 14645 20859 14703 20865
rect 14645 20825 14657 20859
rect 14691 20856 14703 20859
rect 15396 20856 15424 20887
rect 15930 20884 15936 20896
rect 15988 20884 15994 20936
rect 16666 20924 16672 20936
rect 16627 20896 16672 20924
rect 16666 20884 16672 20896
rect 16724 20884 16730 20936
rect 21726 20933 21732 20936
rect 21720 20924 21732 20933
rect 21687 20896 21732 20924
rect 21720 20887 21732 20896
rect 21726 20884 21732 20887
rect 21784 20884 21790 20936
rect 22922 20884 22928 20936
rect 22980 20924 22986 20936
rect 23569 20927 23627 20933
rect 23569 20924 23581 20927
rect 22980 20896 23581 20924
rect 22980 20884 22986 20896
rect 23569 20893 23581 20896
rect 23615 20893 23627 20927
rect 24394 20924 24400 20936
rect 24355 20896 24400 20924
rect 23569 20887 23627 20893
rect 24394 20884 24400 20896
rect 24452 20884 24458 20936
rect 25884 20933 25912 20964
rect 25961 20961 25973 20995
rect 26007 20992 26019 20995
rect 26786 20992 26792 21004
rect 26007 20964 26792 20992
rect 26007 20961 26019 20964
rect 25961 20955 26019 20961
rect 26786 20952 26792 20964
rect 26844 20952 26850 21004
rect 26970 20952 26976 21004
rect 27028 20992 27034 21004
rect 27028 20964 27292 20992
rect 27028 20952 27034 20964
rect 25869 20927 25927 20933
rect 25869 20893 25881 20927
rect 25915 20893 25927 20927
rect 25869 20887 25927 20893
rect 26050 20884 26056 20936
rect 26108 20924 26114 20936
rect 26881 20927 26939 20933
rect 26881 20924 26893 20927
rect 26108 20896 26893 20924
rect 26108 20884 26114 20896
rect 26881 20893 26893 20896
rect 26927 20893 26939 20927
rect 27154 20924 27160 20936
rect 27115 20896 27160 20924
rect 26881 20887 26939 20893
rect 27154 20884 27160 20896
rect 27212 20884 27218 20936
rect 27264 20924 27292 20964
rect 27430 20952 27436 21004
rect 27488 20992 27494 21004
rect 27488 20964 28672 20992
rect 27488 20952 27494 20964
rect 28644 20933 28672 20964
rect 28445 20927 28503 20933
rect 28445 20924 28457 20927
rect 27264 20896 28457 20924
rect 28445 20893 28457 20896
rect 28491 20893 28503 20927
rect 28445 20887 28503 20893
rect 28629 20927 28687 20933
rect 28629 20893 28641 20927
rect 28675 20893 28687 20927
rect 28629 20887 28687 20893
rect 15562 20856 15568 20868
rect 14691 20828 15424 20856
rect 15523 20828 15568 20856
rect 14691 20825 14703 20828
rect 14645 20819 14703 20825
rect 15562 20816 15568 20828
rect 15620 20816 15626 20868
rect 15654 20816 15660 20868
rect 15712 20865 15718 20868
rect 15712 20859 15741 20865
rect 15729 20825 15741 20859
rect 15712 20819 15741 20825
rect 16853 20859 16911 20865
rect 16853 20825 16865 20859
rect 16899 20856 16911 20859
rect 17402 20856 17408 20868
rect 16899 20828 17408 20856
rect 16899 20825 16911 20828
rect 16853 20819 16911 20825
rect 15712 20816 15718 20819
rect 17402 20816 17408 20828
rect 17460 20816 17466 20868
rect 19880 20859 19938 20865
rect 19880 20825 19892 20859
rect 19926 20856 19938 20859
rect 19978 20856 19984 20868
rect 19926 20828 19984 20856
rect 19926 20825 19938 20828
rect 19880 20819 19938 20825
rect 19978 20816 19984 20828
rect 20036 20816 20042 20868
rect 23290 20856 23296 20868
rect 23251 20828 23296 20856
rect 23290 20816 23296 20828
rect 23348 20816 23354 20868
rect 25958 20816 25964 20868
rect 26016 20856 26022 20868
rect 27801 20859 27859 20865
rect 27801 20856 27813 20859
rect 26016 20828 27813 20856
rect 26016 20816 26022 20828
rect 27801 20825 27813 20828
rect 27847 20825 27859 20859
rect 27801 20819 27859 20825
rect 11514 20788 11520 20800
rect 11475 20760 11520 20788
rect 11514 20748 11520 20760
rect 11572 20748 11578 20800
rect 15194 20788 15200 20800
rect 15155 20760 15200 20788
rect 15194 20748 15200 20760
rect 15252 20748 15258 20800
rect 17037 20791 17095 20797
rect 17037 20757 17049 20791
rect 17083 20788 17095 20791
rect 18138 20788 18144 20800
rect 17083 20760 18144 20788
rect 17083 20757 17095 20760
rect 17037 20751 17095 20757
rect 18138 20748 18144 20760
rect 18196 20748 18202 20800
rect 20438 20748 20444 20800
rect 20496 20788 20502 20800
rect 20993 20791 21051 20797
rect 20993 20788 21005 20791
rect 20496 20760 21005 20788
rect 20496 20748 20502 20760
rect 20993 20757 21005 20760
rect 21039 20757 21051 20791
rect 20993 20751 21051 20757
rect 23382 20748 23388 20800
rect 23440 20788 23446 20800
rect 28736 20788 28764 21032
rect 29825 20995 29883 21001
rect 29825 20961 29837 20995
rect 29871 20992 29883 20995
rect 31386 20992 31392 21004
rect 29871 20964 31064 20992
rect 31347 20964 31392 20992
rect 29871 20961 29883 20964
rect 29825 20955 29883 20961
rect 30009 20927 30067 20933
rect 30009 20893 30021 20927
rect 30055 20893 30067 20927
rect 30009 20887 30067 20893
rect 30285 20927 30343 20933
rect 30285 20893 30297 20927
rect 30331 20924 30343 20927
rect 30374 20924 30380 20936
rect 30331 20896 30380 20924
rect 30331 20893 30343 20896
rect 30285 20887 30343 20893
rect 30024 20856 30052 20887
rect 30374 20884 30380 20896
rect 30432 20884 30438 20936
rect 30926 20924 30932 20936
rect 30887 20896 30932 20924
rect 30926 20884 30932 20896
rect 30984 20884 30990 20936
rect 31036 20933 31064 20964
rect 31386 20952 31392 20964
rect 31444 20952 31450 21004
rect 33781 20995 33839 21001
rect 33781 20992 33793 20995
rect 32876 20964 33793 20992
rect 31021 20927 31079 20933
rect 31021 20893 31033 20927
rect 31067 20893 31079 20927
rect 31294 20924 31300 20936
rect 31255 20896 31300 20924
rect 31021 20887 31079 20893
rect 31294 20884 31300 20896
rect 31352 20924 31358 20936
rect 31662 20924 31668 20936
rect 31352 20896 31668 20924
rect 31352 20884 31358 20896
rect 31662 20884 31668 20896
rect 31720 20924 31726 20936
rect 32876 20933 32904 20964
rect 33781 20961 33793 20964
rect 33827 20961 33839 20995
rect 33781 20955 33839 20961
rect 32033 20927 32091 20933
rect 32033 20924 32045 20927
rect 31720 20896 32045 20924
rect 31720 20884 31726 20896
rect 32033 20893 32045 20896
rect 32079 20893 32091 20927
rect 32033 20887 32091 20893
rect 32861 20927 32919 20933
rect 32861 20893 32873 20927
rect 32907 20893 32919 20927
rect 32861 20887 32919 20893
rect 33137 20927 33195 20933
rect 33137 20893 33149 20927
rect 33183 20924 33195 20927
rect 33597 20927 33655 20933
rect 33183 20896 33548 20924
rect 33183 20893 33195 20896
rect 33137 20887 33195 20893
rect 30558 20856 30564 20868
rect 30024 20828 30564 20856
rect 30558 20816 30564 20828
rect 30616 20816 30622 20868
rect 32677 20859 32735 20865
rect 32677 20825 32689 20859
rect 32723 20856 32735 20859
rect 33410 20856 33416 20868
rect 32723 20828 33416 20856
rect 32723 20825 32735 20828
rect 32677 20819 32735 20825
rect 33410 20816 33416 20828
rect 33468 20816 33474 20868
rect 30742 20788 30748 20800
rect 23440 20760 28764 20788
rect 30703 20760 30748 20788
rect 23440 20748 23446 20760
rect 30742 20748 30748 20760
rect 30800 20748 30806 20800
rect 30834 20748 30840 20800
rect 30892 20788 30898 20800
rect 33042 20788 33048 20800
rect 30892 20760 33048 20788
rect 30892 20748 30898 20760
rect 33042 20748 33048 20760
rect 33100 20748 33106 20800
rect 33520 20788 33548 20896
rect 33597 20893 33609 20927
rect 33643 20924 33655 20927
rect 33888 20924 33916 21032
rect 34072 20933 34100 21100
rect 38838 21088 38844 21140
rect 38896 21128 38902 21140
rect 38933 21131 38991 21137
rect 38933 21128 38945 21131
rect 38896 21100 38945 21128
rect 38896 21088 38902 21100
rect 38933 21097 38945 21100
rect 38979 21097 38991 21131
rect 38933 21091 38991 21097
rect 35894 21060 35900 21072
rect 35855 21032 35900 21060
rect 35894 21020 35900 21032
rect 35952 21020 35958 21072
rect 35434 20992 35440 21004
rect 35395 20964 35440 20992
rect 35434 20952 35440 20964
rect 35492 20952 35498 21004
rect 40405 20995 40463 21001
rect 40405 20961 40417 20995
rect 40451 20992 40463 20995
rect 41046 20992 41052 21004
rect 40451 20964 41052 20992
rect 40451 20961 40463 20964
rect 40405 20955 40463 20961
rect 41046 20952 41052 20964
rect 41104 20952 41110 21004
rect 42337 20995 42395 21001
rect 42337 20961 42349 20995
rect 42383 20992 42395 20995
rect 42610 20992 42616 21004
rect 42383 20964 42616 20992
rect 42383 20961 42395 20964
rect 42337 20955 42395 20961
rect 42610 20952 42616 20964
rect 42668 20952 42674 21004
rect 44082 20992 44088 21004
rect 44043 20964 44088 20992
rect 44082 20952 44088 20964
rect 44140 20952 44146 21004
rect 33643 20896 33916 20924
rect 34057 20927 34115 20933
rect 33643 20893 33655 20896
rect 33597 20887 33655 20893
rect 34057 20893 34069 20927
rect 34103 20893 34115 20927
rect 35529 20927 35587 20933
rect 35529 20924 35541 20927
rect 34057 20887 34115 20893
rect 35268 20896 35541 20924
rect 35268 20800 35296 20896
rect 35529 20893 35541 20896
rect 35575 20893 35587 20927
rect 38746 20924 38752 20936
rect 38707 20896 38752 20924
rect 35529 20887 35587 20893
rect 38746 20884 38752 20896
rect 38804 20884 38810 20936
rect 40589 20927 40647 20933
rect 40589 20893 40601 20927
rect 40635 20893 40647 20927
rect 40589 20887 40647 20893
rect 40126 20816 40132 20868
rect 40184 20856 40190 20868
rect 40604 20856 40632 20887
rect 40184 20828 40632 20856
rect 42521 20859 42579 20865
rect 40184 20816 40190 20828
rect 42521 20825 42533 20859
rect 42567 20856 42579 20859
rect 43070 20856 43076 20868
rect 42567 20828 43076 20856
rect 42567 20825 42579 20828
rect 42521 20819 42579 20825
rect 43070 20816 43076 20828
rect 43128 20816 43134 20868
rect 33965 20791 34023 20797
rect 33965 20788 33977 20791
rect 33520 20760 33977 20788
rect 33965 20757 33977 20760
rect 34011 20788 34023 20791
rect 35250 20788 35256 20800
rect 34011 20760 35256 20788
rect 34011 20757 34023 20760
rect 33965 20751 34023 20757
rect 35250 20748 35256 20760
rect 35308 20748 35314 20800
rect 40773 20791 40831 20797
rect 40773 20757 40785 20791
rect 40819 20788 40831 20791
rect 41322 20788 41328 20800
rect 40819 20760 41328 20788
rect 40819 20757 40831 20760
rect 40773 20751 40831 20757
rect 41322 20748 41328 20760
rect 41380 20748 41386 20800
rect 1104 20698 44896 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 44896 20698
rect 1104 20624 44896 20646
rect 15933 20587 15991 20593
rect 15933 20553 15945 20587
rect 15979 20584 15991 20587
rect 16298 20584 16304 20596
rect 15979 20556 16304 20584
rect 15979 20553 15991 20556
rect 15933 20547 15991 20553
rect 16298 20544 16304 20556
rect 16356 20544 16362 20596
rect 16390 20544 16396 20596
rect 16448 20584 16454 20596
rect 18509 20587 18567 20593
rect 16448 20556 17632 20584
rect 16448 20544 16454 20556
rect 15470 20516 15476 20528
rect 14016 20488 15476 20516
rect 1670 20448 1676 20460
rect 1631 20420 1676 20448
rect 1670 20408 1676 20420
rect 1728 20408 1734 20460
rect 11514 20408 11520 20460
rect 11572 20448 11578 20460
rect 12250 20448 12256 20460
rect 11572 20420 12256 20448
rect 11572 20408 11578 20420
rect 12250 20408 12256 20420
rect 12308 20448 12314 20460
rect 14016 20457 14044 20488
rect 15470 20476 15476 20488
rect 15528 20476 15534 20528
rect 17494 20516 17500 20528
rect 17328 20488 17500 20516
rect 12345 20451 12403 20457
rect 12345 20448 12357 20451
rect 12308 20420 12357 20448
rect 12308 20408 12314 20420
rect 12345 20417 12357 20420
rect 12391 20417 12403 20451
rect 12345 20411 12403 20417
rect 14001 20451 14059 20457
rect 14001 20417 14013 20451
rect 14047 20417 14059 20451
rect 14001 20411 14059 20417
rect 14090 20408 14096 20460
rect 14148 20408 14154 20460
rect 14268 20451 14326 20457
rect 14268 20417 14280 20451
rect 14314 20448 14326 20451
rect 15194 20448 15200 20460
rect 14314 20420 15200 20448
rect 14314 20417 14326 20420
rect 14268 20411 14326 20417
rect 15194 20408 15200 20420
rect 15252 20408 15258 20460
rect 15378 20408 15384 20460
rect 15436 20448 15442 20460
rect 16025 20451 16083 20457
rect 16025 20448 16037 20451
rect 15436 20420 16037 20448
rect 15436 20408 15442 20420
rect 16025 20417 16037 20420
rect 16071 20417 16083 20451
rect 16025 20411 16083 20417
rect 1857 20383 1915 20389
rect 1857 20349 1869 20383
rect 1903 20380 1915 20383
rect 2038 20380 2044 20392
rect 1903 20352 2044 20380
rect 1903 20349 1915 20352
rect 1857 20343 1915 20349
rect 2038 20340 2044 20352
rect 2096 20340 2102 20392
rect 2774 20380 2780 20392
rect 2735 20352 2780 20380
rect 2774 20340 2780 20352
rect 2832 20340 2838 20392
rect 12526 20340 12532 20392
rect 12584 20380 12590 20392
rect 12621 20383 12679 20389
rect 12621 20380 12633 20383
rect 12584 20352 12633 20380
rect 12584 20340 12590 20352
rect 12621 20349 12633 20352
rect 12667 20380 12679 20383
rect 14108 20380 14136 20408
rect 12667 20352 14136 20380
rect 16040 20380 16068 20411
rect 17126 20408 17132 20460
rect 17184 20448 17190 20460
rect 17328 20457 17356 20488
rect 17494 20476 17500 20488
rect 17552 20476 17558 20528
rect 17604 20525 17632 20556
rect 18509 20553 18521 20587
rect 18555 20584 18567 20587
rect 18690 20584 18696 20596
rect 18555 20556 18696 20584
rect 18555 20553 18567 20556
rect 18509 20547 18567 20553
rect 18690 20544 18696 20556
rect 18748 20584 18754 20596
rect 19334 20584 19340 20596
rect 18748 20556 19340 20584
rect 18748 20544 18754 20556
rect 19334 20544 19340 20556
rect 19392 20544 19398 20596
rect 19705 20587 19763 20593
rect 19705 20553 19717 20587
rect 19751 20584 19763 20587
rect 19978 20584 19984 20596
rect 19751 20556 19984 20584
rect 19751 20553 19763 20556
rect 19705 20547 19763 20553
rect 19978 20544 19984 20556
rect 20036 20544 20042 20596
rect 37918 20584 37924 20596
rect 22066 20556 37924 20584
rect 17589 20519 17647 20525
rect 17589 20485 17601 20519
rect 17635 20516 17647 20519
rect 19058 20516 19064 20528
rect 17635 20488 19064 20516
rect 17635 20485 17647 20488
rect 17589 20479 17647 20485
rect 19058 20476 19064 20488
rect 19116 20476 19122 20528
rect 19429 20519 19487 20525
rect 19429 20485 19441 20519
rect 19475 20516 19487 20519
rect 22066 20516 22094 20556
rect 37918 20544 37924 20556
rect 37976 20584 37982 20596
rect 41046 20584 41052 20596
rect 37976 20556 40540 20584
rect 41007 20556 41052 20584
rect 37976 20544 37982 20556
rect 19475 20488 20760 20516
rect 19475 20485 19487 20488
rect 19429 20479 19487 20485
rect 17313 20451 17371 20457
rect 17313 20448 17325 20451
rect 17184 20420 17325 20448
rect 17184 20408 17190 20420
rect 17313 20417 17325 20420
rect 17359 20417 17371 20451
rect 17313 20411 17371 20417
rect 17402 20408 17408 20460
rect 17460 20448 17466 20460
rect 18322 20448 18328 20460
rect 17460 20420 18184 20448
rect 18283 20420 18328 20448
rect 17460 20408 17466 20420
rect 17862 20380 17868 20392
rect 16040 20352 17868 20380
rect 12667 20349 12679 20352
rect 12621 20343 12679 20349
rect 17862 20340 17868 20352
rect 17920 20340 17926 20392
rect 18156 20389 18184 20420
rect 18322 20408 18328 20420
rect 18380 20408 18386 20460
rect 19150 20448 19156 20460
rect 19111 20420 19156 20448
rect 19150 20408 19156 20420
rect 19208 20408 19214 20460
rect 19334 20448 19340 20460
rect 19295 20420 19340 20448
rect 19334 20408 19340 20420
rect 19392 20408 19398 20460
rect 19521 20451 19579 20457
rect 19521 20417 19533 20451
rect 19567 20448 19579 20451
rect 19978 20448 19984 20460
rect 19567 20420 19984 20448
rect 19567 20417 19579 20420
rect 19521 20411 19579 20417
rect 19978 20408 19984 20420
rect 20036 20448 20042 20460
rect 20254 20448 20260 20460
rect 20036 20420 20260 20448
rect 20036 20408 20042 20420
rect 20254 20408 20260 20420
rect 20312 20408 20318 20460
rect 20438 20448 20444 20460
rect 20399 20420 20444 20448
rect 20438 20408 20444 20420
rect 20496 20408 20502 20460
rect 18141 20383 18199 20389
rect 18141 20349 18153 20383
rect 18187 20380 18199 20383
rect 20456 20380 20484 20408
rect 20732 20389 20760 20488
rect 21928 20488 22094 20516
rect 18187 20352 20484 20380
rect 20717 20383 20775 20389
rect 18187 20349 18199 20352
rect 18141 20343 18199 20349
rect 20717 20349 20729 20383
rect 20763 20380 20775 20383
rect 20898 20380 20904 20392
rect 20763 20352 20904 20380
rect 20763 20349 20775 20352
rect 20717 20343 20775 20349
rect 20898 20340 20904 20352
rect 20956 20380 20962 20392
rect 21821 20383 21879 20389
rect 21821 20380 21833 20383
rect 20956 20352 21833 20380
rect 20956 20340 20962 20352
rect 21821 20349 21833 20352
rect 21867 20349 21879 20383
rect 21821 20343 21879 20349
rect 21928 20312 21956 20488
rect 22186 20476 22192 20528
rect 22244 20516 22250 20528
rect 26602 20516 26608 20528
rect 22244 20488 26608 20516
rect 22244 20476 22250 20488
rect 26602 20476 26608 20488
rect 26660 20476 26666 20528
rect 29362 20516 29368 20528
rect 29420 20525 29426 20528
rect 29332 20488 29368 20516
rect 29362 20476 29368 20488
rect 29420 20479 29432 20525
rect 31389 20519 31447 20525
rect 31389 20485 31401 20519
rect 31435 20516 31447 20519
rect 32217 20519 32275 20525
rect 32217 20516 32229 20519
rect 31435 20488 32229 20516
rect 31435 20485 31447 20488
rect 31389 20479 31447 20485
rect 32217 20485 32229 20488
rect 32263 20516 32275 20519
rect 32490 20516 32496 20528
rect 32263 20488 32496 20516
rect 32263 20485 32275 20488
rect 32217 20479 32275 20485
rect 29420 20476 29426 20479
rect 32490 20476 32496 20488
rect 32548 20476 32554 20528
rect 35342 20516 35348 20528
rect 33888 20488 35348 20516
rect 22002 20408 22008 20460
rect 22060 20448 22066 20460
rect 23017 20451 23075 20457
rect 23017 20448 23029 20451
rect 22060 20420 23029 20448
rect 22060 20408 22066 20420
rect 23017 20417 23029 20420
rect 23063 20417 23075 20451
rect 23017 20411 23075 20417
rect 24946 20408 24952 20460
rect 25004 20448 25010 20460
rect 25297 20451 25355 20457
rect 25297 20448 25309 20451
rect 25004 20420 25309 20448
rect 25004 20408 25010 20420
rect 25297 20417 25309 20420
rect 25343 20417 25355 20451
rect 25297 20411 25355 20417
rect 29546 20408 29552 20460
rect 29604 20448 29610 20460
rect 29641 20451 29699 20457
rect 29641 20448 29653 20451
rect 29604 20420 29653 20448
rect 29604 20408 29610 20420
rect 29641 20417 29653 20420
rect 29687 20417 29699 20451
rect 29641 20411 29699 20417
rect 30377 20451 30435 20457
rect 30377 20417 30389 20451
rect 30423 20448 30435 20451
rect 30558 20448 30564 20460
rect 30423 20420 30564 20448
rect 30423 20417 30435 20420
rect 30377 20411 30435 20417
rect 30558 20408 30564 20420
rect 30616 20408 30622 20460
rect 31202 20448 31208 20460
rect 31163 20420 31208 20448
rect 31202 20408 31208 20420
rect 31260 20408 31266 20460
rect 31294 20408 31300 20460
rect 31352 20448 31358 20460
rect 31570 20448 31576 20460
rect 31352 20420 31397 20448
rect 31531 20420 31576 20448
rect 31352 20408 31358 20420
rect 31570 20408 31576 20420
rect 31628 20408 31634 20460
rect 31662 20408 31668 20460
rect 31720 20448 31726 20460
rect 32125 20451 32183 20457
rect 32125 20448 32137 20451
rect 31720 20420 32137 20448
rect 31720 20408 31726 20420
rect 32125 20417 32137 20420
rect 32171 20417 32183 20451
rect 32306 20448 32312 20460
rect 32267 20420 32312 20448
rect 32125 20411 32183 20417
rect 32306 20408 32312 20420
rect 32364 20408 32370 20460
rect 33318 20408 33324 20460
rect 33376 20448 33382 20460
rect 33888 20457 33916 20488
rect 35342 20476 35348 20488
rect 35400 20516 35406 20528
rect 40402 20516 40408 20528
rect 35400 20488 40408 20516
rect 35400 20476 35406 20488
rect 37844 20457 37872 20488
rect 38102 20457 38108 20460
rect 33873 20451 33931 20457
rect 33873 20448 33885 20451
rect 33376 20420 33885 20448
rect 33376 20408 33382 20420
rect 33873 20417 33885 20420
rect 33919 20417 33931 20451
rect 34140 20451 34198 20457
rect 34140 20448 34152 20451
rect 33873 20411 33931 20417
rect 33980 20420 34152 20448
rect 23474 20340 23480 20392
rect 23532 20380 23538 20392
rect 24302 20380 24308 20392
rect 23532 20352 24308 20380
rect 23532 20340 23538 20352
rect 24302 20340 24308 20352
rect 24360 20380 24366 20392
rect 24762 20380 24768 20392
rect 24360 20352 24768 20380
rect 24360 20340 24366 20352
rect 24762 20340 24768 20352
rect 24820 20380 24826 20392
rect 25041 20383 25099 20389
rect 25041 20380 25053 20383
rect 24820 20352 25053 20380
rect 24820 20340 24826 20352
rect 25041 20349 25053 20352
rect 25087 20349 25099 20383
rect 25041 20343 25099 20349
rect 30469 20383 30527 20389
rect 30469 20349 30481 20383
rect 30515 20380 30527 20383
rect 31312 20380 31340 20408
rect 30515 20352 31340 20380
rect 30515 20349 30527 20352
rect 30469 20343 30527 20349
rect 33410 20340 33416 20392
rect 33468 20380 33474 20392
rect 33980 20380 34008 20420
rect 34140 20417 34152 20420
rect 34186 20417 34198 20451
rect 34140 20411 34198 20417
rect 37829 20451 37887 20457
rect 37829 20417 37841 20451
rect 37875 20417 37887 20451
rect 38096 20448 38108 20457
rect 38063 20420 38108 20448
rect 37829 20411 37887 20417
rect 38096 20411 38108 20420
rect 38102 20408 38108 20411
rect 38160 20408 38166 20460
rect 39684 20457 39712 20488
rect 40402 20476 40408 20488
rect 40460 20476 40466 20528
rect 39669 20451 39727 20457
rect 39669 20417 39681 20451
rect 39715 20417 39727 20451
rect 39669 20411 39727 20417
rect 39758 20408 39764 20460
rect 39816 20448 39822 20460
rect 39925 20451 39983 20457
rect 39925 20448 39937 20451
rect 39816 20420 39937 20448
rect 39816 20408 39822 20420
rect 39925 20417 39937 20420
rect 39971 20417 39983 20451
rect 40512 20448 40540 20556
rect 41046 20544 41052 20556
rect 41104 20544 41110 20596
rect 43070 20584 43076 20596
rect 43031 20556 43076 20584
rect 43070 20544 43076 20556
rect 43128 20544 43134 20596
rect 42981 20451 43039 20457
rect 42981 20448 42993 20451
rect 40512 20420 42993 20448
rect 39925 20411 39983 20417
rect 42981 20417 42993 20420
rect 43027 20417 43039 20451
rect 42981 20411 43039 20417
rect 33468 20352 34008 20380
rect 33468 20340 33474 20352
rect 15304 20284 21956 20312
rect 8202 20204 8208 20256
rect 8260 20244 8266 20256
rect 15304 20244 15332 20284
rect 22094 20272 22100 20324
rect 22152 20312 22158 20324
rect 22189 20315 22247 20321
rect 22189 20312 22201 20315
rect 22152 20284 22201 20312
rect 22152 20272 22158 20284
rect 22189 20281 22201 20284
rect 22235 20312 22247 20315
rect 23382 20312 23388 20324
rect 22235 20284 23388 20312
rect 22235 20281 22247 20284
rect 22189 20275 22247 20281
rect 23382 20272 23388 20284
rect 23440 20272 23446 20324
rect 26418 20312 26424 20324
rect 26379 20284 26424 20312
rect 26418 20272 26424 20284
rect 26476 20272 26482 20324
rect 35250 20312 35256 20324
rect 35211 20284 35256 20312
rect 35250 20272 35256 20284
rect 35308 20272 35314 20324
rect 8260 20216 15332 20244
rect 15381 20247 15439 20253
rect 8260 20204 8266 20216
rect 15381 20213 15393 20247
rect 15427 20244 15439 20247
rect 15838 20244 15844 20256
rect 15427 20216 15844 20244
rect 15427 20213 15439 20216
rect 15381 20207 15439 20213
rect 15838 20204 15844 20216
rect 15896 20204 15902 20256
rect 22281 20247 22339 20253
rect 22281 20213 22293 20247
rect 22327 20244 22339 20247
rect 22830 20244 22836 20256
rect 22327 20216 22836 20244
rect 22327 20213 22339 20216
rect 22281 20207 22339 20213
rect 22830 20204 22836 20216
rect 22888 20204 22894 20256
rect 23477 20247 23535 20253
rect 23477 20213 23489 20247
rect 23523 20244 23535 20247
rect 24394 20244 24400 20256
rect 23523 20216 24400 20244
rect 23523 20213 23535 20216
rect 23477 20207 23535 20213
rect 24394 20204 24400 20216
rect 24452 20204 24458 20256
rect 31021 20247 31079 20253
rect 31021 20213 31033 20247
rect 31067 20244 31079 20247
rect 31202 20244 31208 20256
rect 31067 20216 31208 20244
rect 31067 20213 31079 20216
rect 31021 20207 31079 20213
rect 31202 20204 31208 20216
rect 31260 20204 31266 20256
rect 39209 20247 39267 20253
rect 39209 20213 39221 20247
rect 39255 20244 39267 20247
rect 39298 20244 39304 20256
rect 39255 20216 39304 20244
rect 39255 20213 39267 20216
rect 39209 20207 39267 20213
rect 39298 20204 39304 20216
rect 39356 20204 39362 20256
rect 43622 20244 43628 20256
rect 43583 20216 43628 20244
rect 43622 20204 43628 20216
rect 43680 20204 43686 20256
rect 1104 20154 44896 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 44896 20154
rect 1104 20080 44896 20102
rect 2038 20040 2044 20052
rect 1999 20012 2044 20040
rect 2038 20000 2044 20012
rect 2096 20000 2102 20052
rect 14550 20000 14556 20052
rect 14608 20040 14614 20052
rect 15013 20043 15071 20049
rect 15013 20040 15025 20043
rect 14608 20012 15025 20040
rect 14608 20000 14614 20012
rect 15013 20009 15025 20012
rect 15059 20009 15071 20043
rect 15013 20003 15071 20009
rect 15197 20043 15255 20049
rect 15197 20009 15209 20043
rect 15243 20040 15255 20043
rect 16390 20040 16396 20052
rect 15243 20012 16396 20040
rect 15243 20009 15255 20012
rect 15197 20003 15255 20009
rect 16390 20000 16396 20012
rect 16448 20000 16454 20052
rect 17221 20043 17279 20049
rect 17221 20009 17233 20043
rect 17267 20040 17279 20043
rect 17402 20040 17408 20052
rect 17267 20012 17408 20040
rect 17267 20009 17279 20012
rect 17221 20003 17279 20009
rect 17402 20000 17408 20012
rect 17460 20000 17466 20052
rect 17862 20000 17868 20052
rect 17920 20040 17926 20052
rect 18325 20043 18383 20049
rect 18325 20040 18337 20043
rect 17920 20012 18337 20040
rect 17920 20000 17926 20012
rect 18325 20009 18337 20012
rect 18371 20009 18383 20043
rect 18325 20003 18383 20009
rect 18509 20043 18567 20049
rect 18509 20009 18521 20043
rect 18555 20040 18567 20043
rect 19334 20040 19340 20052
rect 18555 20012 19340 20040
rect 18555 20009 18567 20012
rect 18509 20003 18567 20009
rect 19334 20000 19340 20012
rect 19392 20000 19398 20052
rect 20070 20040 20076 20052
rect 20031 20012 20076 20040
rect 20070 20000 20076 20012
rect 20128 20000 20134 20052
rect 21818 20040 21824 20052
rect 20180 20012 21824 20040
rect 15562 19932 15568 19984
rect 15620 19972 15626 19984
rect 20180 19972 20208 20012
rect 21818 20000 21824 20012
rect 21876 20000 21882 20052
rect 22278 20040 22284 20052
rect 22239 20012 22284 20040
rect 22278 20000 22284 20012
rect 22336 20000 22342 20052
rect 22738 20000 22744 20052
rect 22796 20040 22802 20052
rect 27430 20040 27436 20052
rect 22796 20012 27016 20040
rect 27391 20012 27436 20040
rect 22796 20000 22802 20012
rect 15620 19944 20208 19972
rect 20257 19975 20315 19981
rect 15620 19932 15626 19944
rect 20257 19941 20269 19975
rect 20303 19972 20315 19975
rect 21174 19972 21180 19984
rect 20303 19944 21180 19972
rect 20303 19941 20315 19944
rect 20257 19935 20315 19941
rect 21174 19932 21180 19944
rect 21232 19932 21238 19984
rect 26988 19972 27016 20012
rect 27430 20000 27436 20012
rect 27488 20000 27494 20052
rect 31205 20043 31263 20049
rect 31205 20009 31217 20043
rect 31251 20040 31263 20043
rect 31570 20040 31576 20052
rect 31251 20012 31576 20040
rect 31251 20009 31263 20012
rect 31205 20003 31263 20009
rect 31570 20000 31576 20012
rect 31628 20000 31634 20052
rect 41414 20040 41420 20052
rect 31726 20012 41420 20040
rect 31726 19972 31754 20012
rect 41414 20000 41420 20012
rect 41472 20000 41478 20052
rect 26988 19944 31754 19972
rect 8846 19864 8852 19916
rect 8904 19904 8910 19916
rect 15838 19904 15844 19916
rect 8904 19876 12434 19904
rect 15799 19876 15844 19904
rect 8904 19864 8910 19876
rect 2130 19836 2136 19848
rect 2091 19808 2136 19836
rect 2130 19796 2136 19808
rect 2188 19836 2194 19848
rect 3970 19836 3976 19848
rect 2188 19808 3976 19836
rect 2188 19796 2194 19808
rect 3970 19796 3976 19808
rect 4028 19796 4034 19848
rect 12250 19836 12256 19848
rect 12211 19808 12256 19836
rect 12250 19796 12256 19808
rect 12308 19796 12314 19848
rect 12406 19768 12434 19876
rect 15838 19864 15844 19876
rect 15896 19904 15902 19916
rect 15896 19876 17448 19904
rect 15896 19864 15902 19876
rect 16117 19839 16175 19845
rect 16117 19805 16129 19839
rect 16163 19805 16175 19839
rect 17126 19836 17132 19848
rect 17087 19808 17132 19836
rect 16117 19799 16175 19805
rect 12802 19768 12808 19780
rect 12406 19740 12808 19768
rect 12802 19728 12808 19740
rect 12860 19768 12866 19780
rect 12897 19771 12955 19777
rect 12897 19768 12909 19771
rect 12860 19740 12909 19768
rect 12860 19728 12866 19740
rect 12897 19737 12909 19740
rect 12943 19737 12955 19771
rect 12897 19731 12955 19737
rect 15181 19771 15239 19777
rect 15181 19737 15193 19771
rect 15227 19768 15239 19771
rect 15286 19768 15292 19780
rect 15227 19740 15292 19768
rect 15227 19737 15239 19740
rect 15181 19731 15239 19737
rect 15286 19728 15292 19740
rect 15344 19728 15350 19780
rect 15381 19771 15439 19777
rect 15381 19737 15393 19771
rect 15427 19768 15439 19771
rect 15930 19768 15936 19780
rect 15427 19740 15936 19768
rect 15427 19737 15439 19740
rect 15381 19731 15439 19737
rect 15930 19728 15936 19740
rect 15988 19768 15994 19780
rect 16132 19768 16160 19799
rect 17126 19796 17132 19808
rect 17184 19796 17190 19848
rect 17420 19845 17448 19876
rect 19904 19876 20944 19904
rect 19904 19845 19932 19876
rect 20916 19848 20944 19876
rect 24762 19864 24768 19916
rect 24820 19904 24826 19916
rect 26053 19907 26111 19913
rect 26053 19904 26065 19907
rect 24820 19876 26065 19904
rect 24820 19864 24826 19876
rect 26053 19873 26065 19876
rect 26099 19873 26111 19907
rect 32490 19904 32496 19916
rect 32451 19876 32496 19904
rect 26053 19867 26111 19873
rect 32490 19864 32496 19876
rect 32548 19864 32554 19916
rect 32950 19904 32956 19916
rect 32911 19876 32956 19904
rect 32950 19864 32956 19876
rect 33008 19864 33014 19916
rect 35342 19864 35348 19916
rect 35400 19904 35406 19916
rect 35437 19907 35495 19913
rect 35437 19904 35449 19907
rect 35400 19876 35449 19904
rect 35400 19864 35406 19876
rect 35437 19873 35449 19876
rect 35483 19873 35495 19907
rect 39298 19904 39304 19916
rect 39259 19876 39304 19904
rect 35437 19867 35495 19873
rect 39298 19864 39304 19876
rect 39356 19864 39362 19916
rect 40405 19907 40463 19913
rect 40405 19904 40417 19907
rect 40052 19876 40417 19904
rect 17405 19839 17463 19845
rect 17405 19805 17417 19839
rect 17451 19805 17463 19839
rect 17405 19799 17463 19805
rect 19889 19839 19947 19845
rect 19889 19805 19901 19839
rect 19935 19805 19947 19839
rect 19889 19799 19947 19805
rect 19981 19839 20039 19845
rect 19981 19805 19993 19839
rect 20027 19805 20039 19839
rect 19981 19799 20039 19805
rect 18138 19768 18144 19780
rect 15988 19740 17724 19768
rect 18099 19740 18144 19768
rect 15988 19728 15994 19740
rect 17696 19712 17724 19740
rect 18138 19728 18144 19740
rect 18196 19728 18202 19780
rect 18322 19728 18328 19780
rect 18380 19777 18386 19780
rect 18380 19771 18404 19777
rect 18392 19737 18404 19771
rect 19996 19768 20024 19799
rect 20070 19796 20076 19848
rect 20128 19836 20134 19848
rect 20717 19839 20775 19845
rect 20717 19836 20729 19839
rect 20128 19808 20729 19836
rect 20128 19796 20134 19808
rect 20717 19805 20729 19808
rect 20763 19805 20775 19839
rect 20898 19836 20904 19848
rect 20859 19808 20904 19836
rect 20717 19799 20775 19805
rect 20898 19796 20904 19808
rect 20956 19796 20962 19848
rect 21545 19839 21603 19845
rect 21545 19805 21557 19839
rect 21591 19836 21603 19839
rect 21591 19808 22784 19836
rect 21591 19805 21603 19808
rect 21545 19799 21603 19805
rect 22189 19771 22247 19777
rect 22189 19768 22201 19771
rect 18380 19731 18404 19737
rect 18432 19740 20024 19768
rect 22066 19740 22201 19768
rect 18380 19728 18386 19731
rect 17494 19660 17500 19712
rect 17552 19700 17558 19712
rect 17589 19703 17647 19709
rect 17589 19700 17601 19703
rect 17552 19672 17601 19700
rect 17552 19660 17558 19672
rect 17589 19669 17601 19672
rect 17635 19669 17647 19703
rect 17589 19663 17647 19669
rect 17678 19660 17684 19712
rect 17736 19700 17742 19712
rect 18432 19700 18460 19740
rect 17736 19672 18460 19700
rect 17736 19660 17742 19672
rect 19058 19660 19064 19712
rect 19116 19700 19122 19712
rect 20254 19700 20260 19712
rect 19116 19672 20260 19700
rect 19116 19660 19122 19672
rect 20254 19660 20260 19672
rect 20312 19660 20318 19712
rect 20346 19660 20352 19712
rect 20404 19700 20410 19712
rect 20809 19703 20867 19709
rect 20809 19700 20821 19703
rect 20404 19672 20821 19700
rect 20404 19660 20410 19672
rect 20809 19669 20821 19672
rect 20855 19669 20867 19703
rect 20809 19663 20867 19669
rect 21453 19703 21511 19709
rect 21453 19669 21465 19703
rect 21499 19700 21511 19703
rect 21634 19700 21640 19712
rect 21499 19672 21640 19700
rect 21499 19669 21511 19672
rect 21453 19663 21511 19669
rect 21634 19660 21640 19672
rect 21692 19700 21698 19712
rect 22066 19700 22094 19740
rect 22189 19737 22201 19740
rect 22235 19737 22247 19771
rect 22756 19768 22784 19808
rect 22830 19796 22836 19848
rect 22888 19836 22894 19848
rect 22888 19808 22933 19836
rect 22888 19796 22894 19808
rect 30558 19796 30564 19848
rect 30616 19836 30622 19848
rect 31021 19839 31079 19845
rect 31021 19836 31033 19839
rect 30616 19808 31033 19836
rect 30616 19796 30622 19808
rect 31021 19805 31033 19808
rect 31067 19805 31079 19839
rect 31021 19799 31079 19805
rect 32585 19839 32643 19845
rect 32585 19805 32597 19839
rect 32631 19836 32643 19839
rect 32674 19836 32680 19848
rect 32631 19808 32680 19836
rect 32631 19805 32643 19808
rect 32585 19799 32643 19805
rect 32674 19796 32680 19808
rect 32732 19836 32738 19848
rect 35693 19839 35751 19845
rect 35693 19836 35705 19839
rect 32732 19808 35705 19836
rect 32732 19796 32738 19808
rect 35693 19805 35705 19808
rect 35739 19805 35751 19839
rect 35693 19799 35751 19805
rect 39117 19839 39175 19845
rect 39117 19805 39129 19839
rect 39163 19836 39175 19839
rect 40052 19836 40080 19876
rect 40405 19873 40417 19876
rect 40451 19904 40463 19907
rect 41598 19904 41604 19916
rect 40451 19876 41604 19904
rect 40451 19873 40463 19876
rect 40405 19867 40463 19873
rect 41598 19864 41604 19876
rect 41656 19864 41662 19916
rect 42058 19904 42064 19916
rect 42019 19876 42064 19904
rect 42058 19864 42064 19876
rect 42116 19864 42122 19916
rect 43070 19904 43076 19916
rect 43031 19876 43076 19904
rect 43070 19864 43076 19876
rect 43128 19864 43134 19916
rect 39163 19808 40080 19836
rect 39163 19805 39175 19808
rect 39117 19799 39175 19805
rect 40126 19796 40132 19848
rect 40184 19836 40190 19848
rect 40184 19808 40229 19836
rect 40184 19796 40190 19808
rect 41506 19796 41512 19848
rect 41564 19836 41570 19848
rect 41877 19839 41935 19845
rect 41877 19836 41889 19839
rect 41564 19808 41889 19836
rect 41564 19796 41570 19808
rect 41877 19805 41889 19808
rect 41923 19805 41935 19839
rect 41877 19799 41935 19805
rect 25314 19768 25320 19780
rect 22756 19740 25320 19768
rect 22189 19731 22247 19737
rect 25314 19728 25320 19740
rect 25372 19728 25378 19780
rect 26326 19777 26332 19780
rect 26320 19731 26332 19777
rect 26384 19768 26390 19780
rect 26384 19740 26420 19768
rect 26326 19728 26332 19731
rect 26384 19728 26390 19740
rect 30374 19728 30380 19780
rect 30432 19768 30438 19780
rect 30837 19771 30895 19777
rect 30837 19768 30849 19771
rect 30432 19740 30849 19768
rect 30432 19728 30438 19740
rect 30837 19737 30849 19740
rect 30883 19737 30895 19771
rect 30837 19731 30895 19737
rect 23014 19700 23020 19712
rect 21692 19672 22094 19700
rect 22975 19672 23020 19700
rect 21692 19660 21698 19672
rect 23014 19660 23020 19672
rect 23072 19660 23078 19712
rect 36817 19703 36875 19709
rect 36817 19669 36829 19703
rect 36863 19700 36875 19703
rect 36906 19700 36912 19712
rect 36863 19672 36912 19700
rect 36863 19669 36875 19672
rect 36817 19663 36875 19669
rect 36906 19660 36912 19672
rect 36964 19660 36970 19712
rect 38930 19700 38936 19712
rect 38891 19672 38936 19700
rect 38930 19660 38936 19672
rect 38988 19660 38994 19712
rect 1104 19610 44896 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 44896 19610
rect 1104 19536 44896 19558
rect 20898 19496 20904 19508
rect 15120 19468 19380 19496
rect 12710 19428 12716 19440
rect 12623 19400 12716 19428
rect 12710 19388 12716 19400
rect 12768 19428 12774 19440
rect 15120 19428 15148 19468
rect 12768 19400 15148 19428
rect 12768 19388 12774 19400
rect 15286 19388 15292 19440
rect 15344 19428 15350 19440
rect 15499 19431 15557 19437
rect 15344 19400 15389 19428
rect 15344 19388 15350 19400
rect 15499 19397 15511 19431
rect 15545 19428 15557 19431
rect 15654 19428 15660 19440
rect 15545 19400 15660 19428
rect 15545 19397 15557 19400
rect 15499 19391 15557 19397
rect 15654 19388 15660 19400
rect 15712 19428 15718 19440
rect 17218 19428 17224 19440
rect 15712 19400 17224 19428
rect 15712 19388 15718 19400
rect 17218 19388 17224 19400
rect 17276 19388 17282 19440
rect 18322 19388 18328 19440
rect 18380 19428 18386 19440
rect 18417 19431 18475 19437
rect 18417 19428 18429 19431
rect 18380 19400 18429 19428
rect 18380 19388 18386 19400
rect 18417 19397 18429 19400
rect 18463 19397 18475 19431
rect 18417 19391 18475 19397
rect 12161 19363 12219 19369
rect 12161 19329 12173 19363
rect 12207 19360 12219 19363
rect 12250 19360 12256 19372
rect 12207 19332 12256 19360
rect 12207 19329 12219 19332
rect 12161 19323 12219 19329
rect 12250 19320 12256 19332
rect 12308 19360 12314 19372
rect 12618 19360 12624 19372
rect 12308 19332 12624 19360
rect 12308 19320 12314 19332
rect 12618 19320 12624 19332
rect 12676 19360 12682 19372
rect 13265 19363 13323 19369
rect 13265 19360 13277 19363
rect 12676 19332 13277 19360
rect 12676 19320 12682 19332
rect 13265 19329 13277 19332
rect 13311 19329 13323 19363
rect 13538 19360 13544 19372
rect 13499 19332 13544 19360
rect 13265 19323 13323 19329
rect 13538 19320 13544 19332
rect 13596 19320 13602 19372
rect 15013 19363 15071 19369
rect 15013 19329 15025 19363
rect 15059 19360 15071 19363
rect 15102 19360 15108 19372
rect 15059 19332 15108 19360
rect 15059 19329 15071 19332
rect 15013 19323 15071 19329
rect 15102 19320 15108 19332
rect 15160 19320 15166 19372
rect 15197 19363 15255 19369
rect 15197 19329 15209 19363
rect 15243 19329 15255 19363
rect 15197 19323 15255 19329
rect 15381 19363 15439 19369
rect 15381 19329 15393 19363
rect 15427 19350 15439 19363
rect 18690 19360 18696 19372
rect 15427 19329 15516 19350
rect 18651 19332 18696 19360
rect 15381 19323 15516 19329
rect 15212 19224 15240 19323
rect 15396 19322 15516 19323
rect 15488 19292 15516 19322
rect 18690 19320 18696 19332
rect 18748 19320 18754 19372
rect 15562 19292 15568 19304
rect 15488 19264 15568 19292
rect 15562 19252 15568 19264
rect 15620 19252 15626 19304
rect 15657 19295 15715 19301
rect 15657 19261 15669 19295
rect 15703 19292 15715 19295
rect 16114 19292 16120 19304
rect 15703 19264 16120 19292
rect 15703 19261 15715 19264
rect 15657 19255 15715 19261
rect 16114 19252 16120 19264
rect 16172 19252 16178 19304
rect 19352 19292 19380 19468
rect 19628 19468 20904 19496
rect 19426 19320 19432 19372
rect 19484 19360 19490 19372
rect 19628 19369 19656 19468
rect 20898 19456 20904 19468
rect 20956 19456 20962 19508
rect 41506 19496 41512 19508
rect 22066 19468 41414 19496
rect 41467 19468 41512 19496
rect 22066 19428 22094 19468
rect 19812 19400 20392 19428
rect 19812 19369 19840 19400
rect 20364 19372 20392 19400
rect 20456 19400 22094 19428
rect 19521 19363 19579 19369
rect 19521 19360 19533 19363
rect 19484 19332 19533 19360
rect 19484 19320 19490 19332
rect 19521 19329 19533 19332
rect 19567 19329 19579 19363
rect 19521 19323 19579 19329
rect 19613 19363 19671 19369
rect 19613 19329 19625 19363
rect 19659 19329 19671 19363
rect 19613 19323 19671 19329
rect 19797 19363 19855 19369
rect 19797 19329 19809 19363
rect 19843 19329 19855 19363
rect 19797 19323 19855 19329
rect 19889 19363 19947 19369
rect 19889 19329 19901 19363
rect 19935 19360 19947 19363
rect 20070 19360 20076 19372
rect 19935 19332 20076 19360
rect 19935 19329 19947 19332
rect 19889 19323 19947 19329
rect 20070 19320 20076 19332
rect 20128 19320 20134 19372
rect 20346 19360 20352 19372
rect 20307 19332 20352 19360
rect 20346 19320 20352 19332
rect 20404 19320 20410 19372
rect 20456 19292 20484 19400
rect 22186 19388 22192 19440
rect 22244 19428 22250 19440
rect 22244 19400 22289 19428
rect 22244 19388 22250 19400
rect 23014 19388 23020 19440
rect 23072 19428 23078 19440
rect 23722 19431 23780 19437
rect 23722 19428 23734 19431
rect 23072 19400 23734 19428
rect 23072 19388 23078 19400
rect 23722 19397 23734 19400
rect 23768 19397 23780 19431
rect 23722 19391 23780 19397
rect 30460 19431 30518 19437
rect 30460 19397 30472 19431
rect 30506 19428 30518 19431
rect 30926 19428 30932 19440
rect 30506 19400 30932 19428
rect 30506 19397 30518 19400
rect 30460 19391 30518 19397
rect 30926 19388 30932 19400
rect 30984 19388 30990 19440
rect 32950 19388 32956 19440
rect 33008 19428 33014 19440
rect 33566 19431 33624 19437
rect 33566 19428 33578 19431
rect 33008 19400 33578 19428
rect 33008 19388 33014 19400
rect 33566 19397 33578 19400
rect 33612 19397 33624 19431
rect 41386 19428 41414 19468
rect 41506 19456 41512 19468
rect 41564 19456 41570 19508
rect 43714 19428 43720 19440
rect 41386 19400 43720 19428
rect 33566 19391 33624 19397
rect 43714 19388 43720 19400
rect 43772 19388 43778 19440
rect 20625 19363 20683 19369
rect 20625 19329 20637 19363
rect 20671 19360 20683 19363
rect 21542 19360 21548 19372
rect 20671 19332 21548 19360
rect 20671 19329 20683 19332
rect 20625 19323 20683 19329
rect 21542 19320 21548 19332
rect 21600 19320 21606 19372
rect 23474 19360 23480 19372
rect 23435 19332 23480 19360
rect 23474 19320 23480 19332
rect 23532 19320 23538 19372
rect 26694 19320 26700 19372
rect 26752 19360 26758 19372
rect 27157 19363 27215 19369
rect 27157 19360 27169 19363
rect 26752 19332 27169 19360
rect 26752 19320 26758 19332
rect 27157 19329 27169 19332
rect 27203 19329 27215 19363
rect 27157 19323 27215 19329
rect 27341 19363 27399 19369
rect 27341 19329 27353 19363
rect 27387 19360 27399 19363
rect 28350 19360 28356 19372
rect 27387 19332 28356 19360
rect 27387 19329 27399 19332
rect 27341 19323 27399 19329
rect 28350 19320 28356 19332
rect 28408 19320 28414 19372
rect 33318 19360 33324 19372
rect 33279 19332 33324 19360
rect 33318 19320 33324 19332
rect 33376 19320 33382 19372
rect 38930 19360 38936 19372
rect 38891 19332 38936 19360
rect 38930 19320 38936 19332
rect 38988 19320 38994 19372
rect 41322 19360 41328 19372
rect 41283 19332 41328 19360
rect 41322 19320 41328 19332
rect 41380 19320 41386 19372
rect 41414 19320 41420 19372
rect 41472 19360 41478 19372
rect 42889 19363 42947 19369
rect 42889 19360 42901 19363
rect 41472 19332 42901 19360
rect 41472 19320 41478 19332
rect 42889 19329 42901 19332
rect 42935 19329 42947 19363
rect 42889 19323 42947 19329
rect 42978 19320 42984 19372
rect 43036 19360 43042 19372
rect 43036 19332 43081 19360
rect 43036 19320 43042 19332
rect 19352 19264 20484 19292
rect 20809 19295 20867 19301
rect 20809 19261 20821 19295
rect 20855 19292 20867 19295
rect 23106 19292 23112 19304
rect 20855 19264 23112 19292
rect 20855 19261 20867 19264
rect 20809 19255 20867 19261
rect 23106 19252 23112 19264
rect 23164 19252 23170 19304
rect 26973 19295 27031 19301
rect 26973 19261 26985 19295
rect 27019 19292 27031 19295
rect 27062 19292 27068 19304
rect 27019 19264 27068 19292
rect 27019 19261 27031 19264
rect 26973 19255 27031 19261
rect 27062 19252 27068 19264
rect 27120 19252 27126 19304
rect 29546 19252 29552 19304
rect 29604 19292 29610 19304
rect 30193 19295 30251 19301
rect 30193 19292 30205 19295
rect 29604 19264 30205 19292
rect 29604 19252 29610 19264
rect 30193 19261 30205 19264
rect 30239 19261 30251 19295
rect 30193 19255 30251 19261
rect 15286 19224 15292 19236
rect 15212 19196 15292 19224
rect 15286 19184 15292 19196
rect 15344 19184 15350 19236
rect 20254 19184 20260 19236
rect 20312 19224 20318 19236
rect 20441 19227 20499 19233
rect 20441 19224 20453 19227
rect 20312 19196 20453 19224
rect 20312 19184 20318 19196
rect 20441 19193 20453 19196
rect 20487 19193 20499 19227
rect 20441 19187 20499 19193
rect 21082 19184 21088 19236
rect 21140 19224 21146 19236
rect 21821 19227 21879 19233
rect 21821 19224 21833 19227
rect 21140 19196 21833 19224
rect 21140 19184 21146 19196
rect 21821 19193 21833 19196
rect 21867 19193 21879 19227
rect 21821 19187 21879 19193
rect 19334 19156 19340 19168
rect 19295 19128 19340 19156
rect 19334 19116 19340 19128
rect 19392 19116 19398 19168
rect 21174 19116 21180 19168
rect 21232 19156 21238 19168
rect 22189 19159 22247 19165
rect 22189 19156 22201 19159
rect 21232 19128 22201 19156
rect 21232 19116 21238 19128
rect 22189 19125 22201 19128
rect 22235 19125 22247 19159
rect 22189 19119 22247 19125
rect 22373 19159 22431 19165
rect 22373 19125 22385 19159
rect 22419 19156 22431 19159
rect 23014 19156 23020 19168
rect 22419 19128 23020 19156
rect 22419 19125 22431 19128
rect 22373 19119 22431 19125
rect 23014 19116 23020 19128
rect 23072 19116 23078 19168
rect 24854 19156 24860 19168
rect 24815 19128 24860 19156
rect 24854 19116 24860 19128
rect 24912 19116 24918 19168
rect 31570 19156 31576 19168
rect 31531 19128 31576 19156
rect 31570 19116 31576 19128
rect 31628 19116 31634 19168
rect 34698 19156 34704 19168
rect 34659 19128 34704 19156
rect 34698 19116 34704 19128
rect 34756 19116 34762 19168
rect 38746 19156 38752 19168
rect 38707 19128 38752 19156
rect 38746 19116 38752 19128
rect 38804 19116 38810 19168
rect 43809 19159 43867 19165
rect 43809 19125 43821 19159
rect 43855 19156 43867 19159
rect 44174 19156 44180 19168
rect 43855 19128 44180 19156
rect 43855 19125 43867 19128
rect 43809 19119 43867 19125
rect 44174 19116 44180 19128
rect 44232 19116 44238 19168
rect 1104 19066 44896 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 44896 19066
rect 1104 18992 44896 19014
rect 13538 18912 13544 18964
rect 13596 18952 13602 18964
rect 13596 18924 15516 18952
rect 13596 18912 13602 18924
rect 15488 18884 15516 18924
rect 16942 18912 16948 18964
rect 17000 18952 17006 18964
rect 17129 18955 17187 18961
rect 17129 18952 17141 18955
rect 17000 18924 17141 18952
rect 17000 18912 17006 18924
rect 17129 18921 17141 18924
rect 17175 18921 17187 18955
rect 17129 18915 17187 18921
rect 18509 18955 18567 18961
rect 18509 18921 18521 18955
rect 18555 18952 18567 18955
rect 19334 18952 19340 18964
rect 18555 18924 19340 18952
rect 18555 18921 18567 18924
rect 18509 18915 18567 18921
rect 19334 18912 19340 18924
rect 19392 18912 19398 18964
rect 25823 18955 25881 18961
rect 25823 18921 25835 18955
rect 25869 18952 25881 18955
rect 26418 18952 26424 18964
rect 25869 18924 26424 18952
rect 25869 18921 25881 18924
rect 25823 18915 25881 18921
rect 26418 18912 26424 18924
rect 26476 18912 26482 18964
rect 27448 18924 37780 18952
rect 23842 18884 23848 18896
rect 15488 18856 18736 18884
rect 15470 18816 15476 18828
rect 15431 18788 15476 18816
rect 15470 18776 15476 18788
rect 15528 18776 15534 18828
rect 17313 18819 17371 18825
rect 17313 18785 17325 18819
rect 17359 18816 17371 18819
rect 17678 18816 17684 18828
rect 17359 18788 17684 18816
rect 17359 18785 17371 18788
rect 17313 18779 17371 18785
rect 17678 18776 17684 18788
rect 17736 18776 17742 18828
rect 2038 18748 2044 18760
rect 1999 18720 2044 18748
rect 2038 18708 2044 18720
rect 2096 18708 2102 18760
rect 12618 18708 12624 18760
rect 12676 18748 12682 18760
rect 12713 18751 12771 18757
rect 12713 18748 12725 18751
rect 12676 18720 12725 18748
rect 12676 18708 12682 18720
rect 12713 18717 12725 18720
rect 12759 18717 12771 18751
rect 12713 18711 12771 18717
rect 15194 18708 15200 18760
rect 15252 18757 15258 18760
rect 15252 18748 15264 18757
rect 15933 18751 15991 18757
rect 15252 18720 15297 18748
rect 15252 18711 15264 18720
rect 15933 18717 15945 18751
rect 15979 18717 15991 18751
rect 16114 18748 16120 18760
rect 16075 18720 16120 18748
rect 15933 18711 15991 18717
rect 15252 18708 15258 18711
rect 11698 18640 11704 18692
rect 11756 18680 11762 18692
rect 12161 18683 12219 18689
rect 12161 18680 12173 18683
rect 11756 18652 12173 18680
rect 11756 18640 11762 18652
rect 12161 18649 12173 18652
rect 12207 18649 12219 18683
rect 12161 18643 12219 18649
rect 14550 18640 14556 18692
rect 14608 18680 14614 18692
rect 15948 18680 15976 18711
rect 16114 18708 16120 18720
rect 16172 18708 16178 18760
rect 17126 18748 17132 18760
rect 17087 18720 17132 18748
rect 17126 18708 17132 18720
rect 17184 18708 17190 18760
rect 17402 18748 17408 18760
rect 17363 18720 17408 18748
rect 17402 18708 17408 18720
rect 17460 18708 17466 18760
rect 18322 18748 18328 18760
rect 18283 18720 18328 18748
rect 18322 18708 18328 18720
rect 18380 18708 18386 18760
rect 18598 18748 18604 18760
rect 18559 18720 18604 18748
rect 18598 18708 18604 18720
rect 18656 18708 18662 18760
rect 18708 18748 18736 18856
rect 22066 18856 23848 18884
rect 21542 18776 21548 18828
rect 21600 18816 21606 18828
rect 21637 18819 21695 18825
rect 21637 18816 21649 18819
rect 21600 18788 21649 18816
rect 21600 18776 21606 18788
rect 21637 18785 21649 18788
rect 21683 18785 21695 18819
rect 21637 18779 21695 18785
rect 21818 18776 21824 18828
rect 21876 18816 21882 18828
rect 21913 18819 21971 18825
rect 21913 18816 21925 18819
rect 21876 18788 21925 18816
rect 21876 18776 21882 18788
rect 21913 18785 21925 18788
rect 21959 18816 21971 18819
rect 22066 18816 22094 18856
rect 23842 18844 23848 18856
rect 23900 18844 23906 18896
rect 25961 18887 26019 18893
rect 25961 18853 25973 18887
rect 26007 18884 26019 18887
rect 26234 18884 26240 18896
rect 26007 18856 26240 18884
rect 26007 18853 26019 18856
rect 25961 18847 26019 18853
rect 26234 18844 26240 18856
rect 26292 18844 26298 18896
rect 27448 18816 27476 18924
rect 21959 18788 22094 18816
rect 22848 18788 27476 18816
rect 21959 18785 21971 18788
rect 21913 18779 21971 18785
rect 22848 18748 22876 18788
rect 34606 18776 34612 18828
rect 34664 18816 34670 18828
rect 34793 18819 34851 18825
rect 34793 18816 34805 18819
rect 34664 18788 34805 18816
rect 34664 18776 34670 18788
rect 34793 18785 34805 18788
rect 34839 18816 34851 18819
rect 34974 18816 34980 18828
rect 34839 18788 34980 18816
rect 34839 18785 34851 18788
rect 34793 18779 34851 18785
rect 34974 18776 34980 18788
rect 35032 18776 35038 18828
rect 35250 18816 35256 18828
rect 35211 18788 35256 18816
rect 35250 18776 35256 18788
rect 35308 18776 35314 18828
rect 36832 18788 37504 18816
rect 23014 18748 23020 18760
rect 18708 18720 22876 18748
rect 22975 18720 23020 18748
rect 23014 18708 23020 18720
rect 23072 18708 23078 18760
rect 24854 18708 24860 18760
rect 24912 18748 24918 18760
rect 25682 18748 25688 18760
rect 24912 18720 25688 18748
rect 24912 18708 24918 18720
rect 25682 18708 25688 18720
rect 25740 18708 25746 18760
rect 26145 18751 26203 18757
rect 26145 18748 26157 18751
rect 26068 18720 26157 18748
rect 16758 18680 16764 18692
rect 14608 18652 16764 18680
rect 14608 18640 14614 18652
rect 16758 18640 16764 18652
rect 16816 18640 16822 18692
rect 17494 18640 17500 18692
rect 17552 18680 17558 18692
rect 19426 18680 19432 18692
rect 17552 18652 19432 18680
rect 17552 18640 17558 18652
rect 19426 18640 19432 18652
rect 19484 18640 19490 18692
rect 25958 18640 25964 18692
rect 26016 18680 26022 18692
rect 26068 18680 26096 18720
rect 26145 18717 26157 18720
rect 26191 18717 26203 18751
rect 26145 18711 26203 18717
rect 26418 18708 26424 18760
rect 26476 18748 26482 18760
rect 26789 18751 26847 18757
rect 26789 18748 26801 18751
rect 26476 18720 26801 18748
rect 26476 18708 26482 18720
rect 26789 18717 26801 18720
rect 26835 18717 26847 18751
rect 26970 18748 26976 18760
rect 26931 18720 26976 18748
rect 26789 18711 26847 18717
rect 26970 18708 26976 18720
rect 27028 18708 27034 18760
rect 28350 18748 28356 18760
rect 28311 18720 28356 18748
rect 28350 18708 28356 18720
rect 28408 18708 28414 18760
rect 31205 18751 31263 18757
rect 31205 18748 31217 18751
rect 29932 18720 31217 18748
rect 26016 18652 26096 18680
rect 28537 18683 28595 18689
rect 26016 18640 26022 18652
rect 28537 18649 28549 18683
rect 28583 18680 28595 18683
rect 29454 18680 29460 18692
rect 28583 18652 29460 18680
rect 28583 18649 28595 18652
rect 28537 18643 28595 18649
rect 29454 18640 29460 18652
rect 29512 18640 29518 18692
rect 29546 18640 29552 18692
rect 29604 18680 29610 18692
rect 29932 18689 29960 18720
rect 31205 18717 31217 18720
rect 31251 18717 31263 18751
rect 31205 18711 31263 18717
rect 31294 18708 31300 18760
rect 31352 18748 31358 18760
rect 31461 18751 31519 18757
rect 31461 18748 31473 18751
rect 31352 18720 31473 18748
rect 31352 18708 31358 18720
rect 31461 18717 31473 18720
rect 31507 18717 31519 18751
rect 31461 18711 31519 18717
rect 34698 18708 34704 18760
rect 34756 18748 34762 18760
rect 34882 18748 34888 18760
rect 34756 18720 34888 18748
rect 34756 18708 34762 18720
rect 34882 18708 34888 18720
rect 34940 18708 34946 18760
rect 36832 18757 36860 18788
rect 36817 18751 36875 18757
rect 36817 18717 36829 18751
rect 36863 18717 36875 18751
rect 36817 18711 36875 18717
rect 29917 18683 29975 18689
rect 29917 18680 29929 18683
rect 29604 18652 29929 18680
rect 29604 18640 29610 18652
rect 29917 18649 29929 18652
rect 29963 18649 29975 18683
rect 29917 18643 29975 18649
rect 30101 18683 30159 18689
rect 30101 18649 30113 18683
rect 30147 18680 30159 18683
rect 30558 18680 30564 18692
rect 30147 18652 30564 18680
rect 30147 18649 30159 18652
rect 30101 18643 30159 18649
rect 30558 18640 30564 18652
rect 30616 18640 30622 18692
rect 34422 18640 34428 18692
rect 34480 18680 34486 18692
rect 36832 18680 36860 18711
rect 36906 18708 36912 18760
rect 36964 18748 36970 18760
rect 37476 18757 37504 18788
rect 37461 18751 37519 18757
rect 36964 18720 37009 18748
rect 36964 18708 36970 18720
rect 37461 18717 37473 18751
rect 37507 18717 37519 18751
rect 37461 18711 37519 18717
rect 37645 18751 37703 18757
rect 37645 18717 37657 18751
rect 37691 18717 37703 18751
rect 37752 18748 37780 18924
rect 43254 18884 43260 18896
rect 41386 18856 43260 18884
rect 38289 18751 38347 18757
rect 38289 18748 38301 18751
rect 37752 18720 38301 18748
rect 37645 18711 37703 18717
rect 38289 18717 38301 18720
rect 38335 18748 38347 18751
rect 41386 18748 41414 18856
rect 43254 18844 43260 18856
rect 43312 18844 43318 18896
rect 42702 18816 42708 18828
rect 42663 18788 42708 18816
rect 42702 18776 42708 18788
rect 42760 18776 42766 18828
rect 44174 18816 44180 18828
rect 44135 18788 44180 18816
rect 44174 18776 44180 18788
rect 44232 18776 44238 18828
rect 38335 18720 41414 18748
rect 38335 18717 38347 18720
rect 38289 18711 38347 18717
rect 34480 18652 36860 18680
rect 36924 18680 36952 18708
rect 37660 18680 37688 18711
rect 36924 18652 37688 18680
rect 34480 18640 34486 18652
rect 43438 18640 43444 18692
rect 43496 18680 43502 18692
rect 43993 18683 44051 18689
rect 43993 18680 44005 18683
rect 43496 18652 44005 18680
rect 43496 18640 43502 18652
rect 43993 18649 44005 18652
rect 44039 18649 44051 18683
rect 43993 18643 44051 18649
rect 14093 18615 14151 18621
rect 14093 18581 14105 18615
rect 14139 18612 14151 18615
rect 14734 18612 14740 18624
rect 14139 18584 14740 18612
rect 14139 18581 14151 18584
rect 14093 18575 14151 18581
rect 14734 18572 14740 18584
rect 14792 18572 14798 18624
rect 16022 18612 16028 18624
rect 15983 18584 16028 18612
rect 16022 18572 16028 18584
rect 16080 18572 16086 18624
rect 17586 18612 17592 18624
rect 17547 18584 17592 18612
rect 17586 18572 17592 18584
rect 17644 18572 17650 18624
rect 18046 18612 18052 18624
rect 18007 18584 18052 18612
rect 18046 18572 18052 18584
rect 18104 18572 18110 18624
rect 23201 18615 23259 18621
rect 23201 18581 23213 18615
rect 23247 18612 23259 18615
rect 25130 18612 25136 18624
rect 23247 18584 25136 18612
rect 23247 18581 23259 18584
rect 23201 18575 23259 18581
rect 25130 18572 25136 18584
rect 25188 18572 25194 18624
rect 26145 18615 26203 18621
rect 26145 18581 26157 18615
rect 26191 18612 26203 18615
rect 27062 18612 27068 18624
rect 26191 18584 27068 18612
rect 26191 18581 26203 18584
rect 26145 18575 26203 18581
rect 27062 18572 27068 18584
rect 27120 18572 27126 18624
rect 27798 18612 27804 18624
rect 27759 18584 27804 18612
rect 27798 18572 27804 18584
rect 27856 18572 27862 18624
rect 32582 18612 32588 18624
rect 32543 18584 32588 18612
rect 32582 18572 32588 18584
rect 32640 18572 32646 18624
rect 35710 18572 35716 18624
rect 35768 18612 35774 18624
rect 36633 18615 36691 18621
rect 36633 18612 36645 18615
rect 35768 18584 36645 18612
rect 35768 18572 35774 18584
rect 36633 18581 36645 18584
rect 36679 18581 36691 18615
rect 36633 18575 36691 18581
rect 37458 18572 37464 18624
rect 37516 18612 37522 18624
rect 37553 18615 37611 18621
rect 37553 18612 37565 18615
rect 37516 18584 37565 18612
rect 37516 18572 37522 18584
rect 37553 18581 37565 18584
rect 37599 18581 37611 18615
rect 38378 18612 38384 18624
rect 38339 18584 38384 18612
rect 37553 18575 37611 18581
rect 38378 18572 38384 18584
rect 38436 18572 38442 18624
rect 1104 18522 44896 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 44896 18522
rect 1104 18448 44896 18470
rect 6270 18368 6276 18420
rect 6328 18408 6334 18420
rect 6822 18408 6828 18420
rect 6328 18380 6828 18408
rect 6328 18368 6334 18380
rect 6822 18368 6828 18380
rect 6880 18408 6886 18420
rect 43438 18408 43444 18420
rect 6880 18380 41414 18408
rect 43399 18380 43444 18408
rect 6880 18368 6886 18380
rect 16022 18340 16028 18352
rect 13832 18312 16028 18340
rect 2038 18272 2044 18284
rect 1999 18244 2044 18272
rect 2038 18232 2044 18244
rect 2096 18232 2102 18284
rect 13832 18281 13860 18312
rect 16022 18300 16028 18312
rect 16080 18300 16086 18352
rect 16758 18300 16764 18352
rect 16816 18349 16822 18352
rect 16816 18343 16879 18349
rect 16816 18309 16833 18343
rect 16867 18309 16879 18343
rect 17034 18340 17040 18352
rect 16995 18312 17040 18340
rect 16816 18303 16879 18309
rect 16816 18300 16822 18303
rect 17034 18300 17040 18312
rect 17092 18300 17098 18352
rect 17586 18300 17592 18352
rect 17644 18340 17650 18352
rect 18509 18343 18567 18349
rect 18509 18340 18521 18343
rect 17644 18312 18521 18340
rect 17644 18300 17650 18312
rect 18509 18309 18521 18312
rect 18555 18309 18567 18343
rect 18509 18303 18567 18309
rect 19426 18300 19432 18352
rect 19484 18340 19490 18352
rect 23474 18340 23480 18352
rect 19484 18312 20484 18340
rect 19484 18300 19490 18312
rect 13817 18275 13875 18281
rect 13817 18241 13829 18275
rect 13863 18241 13875 18275
rect 13817 18235 13875 18241
rect 14001 18275 14059 18281
rect 14001 18241 14013 18275
rect 14047 18272 14059 18275
rect 14458 18272 14464 18284
rect 14047 18244 14464 18272
rect 14047 18241 14059 18244
rect 14001 18235 14059 18241
rect 14458 18232 14464 18244
rect 14516 18232 14522 18284
rect 14550 18232 14556 18284
rect 14608 18272 14614 18284
rect 14645 18275 14703 18281
rect 14645 18272 14657 18275
rect 14608 18244 14657 18272
rect 14608 18232 14614 18244
rect 14645 18241 14657 18244
rect 14691 18241 14703 18275
rect 14645 18235 14703 18241
rect 14734 18232 14740 18284
rect 14792 18272 14798 18284
rect 16117 18275 16175 18281
rect 16117 18272 16129 18275
rect 14792 18244 16129 18272
rect 14792 18232 14798 18244
rect 16117 18241 16129 18244
rect 16163 18272 16175 18275
rect 16942 18272 16948 18284
rect 16163 18244 16948 18272
rect 16163 18241 16175 18244
rect 16117 18235 16175 18241
rect 16942 18232 16948 18244
rect 17000 18232 17006 18284
rect 17678 18232 17684 18284
rect 17736 18272 17742 18284
rect 17773 18275 17831 18281
rect 17773 18272 17785 18275
rect 17736 18244 17785 18272
rect 17736 18232 17742 18244
rect 17773 18241 17785 18244
rect 17819 18241 17831 18275
rect 17773 18235 17831 18241
rect 17957 18275 18015 18281
rect 17957 18241 17969 18275
rect 18003 18272 18015 18275
rect 18138 18272 18144 18284
rect 18003 18244 18144 18272
rect 18003 18241 18015 18244
rect 17957 18235 18015 18241
rect 18138 18232 18144 18244
rect 18196 18232 18202 18284
rect 18690 18272 18696 18284
rect 18651 18244 18696 18272
rect 18690 18232 18696 18244
rect 18748 18232 18754 18284
rect 20456 18281 20484 18312
rect 23032 18312 23480 18340
rect 19613 18275 19671 18281
rect 19613 18272 19625 18275
rect 18984 18244 19625 18272
rect 2225 18207 2283 18213
rect 2225 18173 2237 18207
rect 2271 18204 2283 18207
rect 2866 18204 2872 18216
rect 2271 18176 2872 18204
rect 2271 18173 2283 18176
rect 2225 18167 2283 18173
rect 2866 18164 2872 18176
rect 2924 18164 2930 18216
rect 2958 18164 2964 18216
rect 3016 18204 3022 18216
rect 15841 18207 15899 18213
rect 3016 18176 3061 18204
rect 3016 18164 3022 18176
rect 15841 18173 15853 18207
rect 15887 18204 15899 18207
rect 16022 18204 16028 18216
rect 15887 18176 16028 18204
rect 15887 18173 15899 18176
rect 15841 18167 15899 18173
rect 16022 18164 16028 18176
rect 16080 18204 16086 18216
rect 18049 18207 18107 18213
rect 16080 18176 18000 18204
rect 16080 18164 16086 18176
rect 14001 18139 14059 18145
rect 14001 18105 14013 18139
rect 14047 18136 14059 18139
rect 15286 18136 15292 18148
rect 14047 18108 15292 18136
rect 14047 18105 14059 18108
rect 14001 18099 14059 18105
rect 15286 18096 15292 18108
rect 15344 18096 15350 18148
rect 17034 18096 17040 18148
rect 17092 18136 17098 18148
rect 17972 18136 18000 18176
rect 18049 18173 18061 18207
rect 18095 18204 18107 18207
rect 18322 18204 18328 18216
rect 18095 18176 18328 18204
rect 18095 18173 18107 18176
rect 18049 18167 18107 18173
rect 18322 18164 18328 18176
rect 18380 18204 18386 18216
rect 18877 18207 18935 18213
rect 18877 18204 18889 18207
rect 18380 18176 18889 18204
rect 18380 18164 18386 18176
rect 18877 18173 18889 18176
rect 18923 18173 18935 18207
rect 18877 18167 18935 18173
rect 18984 18136 19012 18244
rect 19613 18241 19625 18244
rect 19659 18272 19671 18275
rect 20257 18275 20315 18281
rect 20257 18272 20269 18275
rect 19659 18244 20269 18272
rect 19659 18241 19671 18244
rect 19613 18235 19671 18241
rect 20257 18241 20269 18244
rect 20303 18241 20315 18275
rect 20257 18235 20315 18241
rect 20441 18275 20499 18281
rect 20441 18241 20453 18275
rect 20487 18272 20499 18275
rect 21082 18272 21088 18284
rect 20487 18244 21088 18272
rect 20487 18241 20499 18244
rect 20441 18235 20499 18241
rect 19337 18207 19395 18213
rect 19337 18204 19349 18207
rect 17092 18108 17708 18136
rect 17972 18108 19012 18136
rect 19076 18176 19349 18204
rect 17092 18096 17098 18108
rect 14458 18068 14464 18080
rect 14419 18040 14464 18068
rect 14458 18028 14464 18040
rect 14516 18028 14522 18080
rect 16666 18068 16672 18080
rect 16627 18040 16672 18068
rect 16666 18028 16672 18040
rect 16724 18028 16730 18080
rect 16850 18028 16856 18080
rect 16908 18077 16914 18080
rect 16908 18068 16920 18077
rect 17586 18068 17592 18080
rect 16908 18040 16953 18068
rect 17547 18040 17592 18068
rect 16908 18031 16920 18040
rect 16908 18028 16914 18031
rect 17586 18028 17592 18040
rect 17644 18028 17650 18080
rect 17680 18068 17708 18108
rect 19076 18068 19104 18176
rect 19337 18173 19349 18176
rect 19383 18173 19395 18207
rect 19337 18167 19395 18173
rect 19426 18164 19432 18216
rect 19484 18204 19490 18216
rect 19521 18207 19579 18213
rect 19521 18204 19533 18207
rect 19484 18176 19533 18204
rect 19484 18164 19490 18176
rect 19521 18173 19533 18176
rect 19567 18173 19579 18207
rect 20272 18204 20300 18235
rect 21082 18232 21088 18244
rect 21140 18232 21146 18284
rect 21542 18232 21548 18284
rect 21600 18272 21606 18284
rect 23032 18281 23060 18312
rect 23474 18300 23480 18312
rect 23532 18300 23538 18352
rect 25130 18349 25136 18352
rect 25124 18340 25136 18349
rect 25091 18312 25136 18340
rect 25124 18303 25136 18312
rect 25130 18300 25136 18303
rect 25188 18300 25194 18352
rect 26234 18300 26240 18352
rect 26292 18340 26298 18352
rect 27525 18343 27583 18349
rect 27525 18340 27537 18343
rect 26292 18312 27537 18340
rect 26292 18300 26298 18312
rect 27525 18309 27537 18312
rect 27571 18309 27583 18343
rect 27525 18303 27583 18309
rect 27798 18300 27804 18352
rect 27856 18340 27862 18352
rect 28620 18343 28678 18349
rect 28620 18340 28632 18343
rect 27856 18312 28632 18340
rect 27856 18300 27862 18312
rect 28620 18309 28632 18312
rect 28666 18340 28678 18343
rect 34422 18340 34428 18352
rect 28666 18312 34428 18340
rect 28666 18309 28678 18312
rect 28620 18303 28678 18309
rect 34422 18300 34428 18312
rect 34480 18300 34486 18352
rect 34882 18340 34888 18352
rect 34843 18312 34888 18340
rect 34882 18300 34888 18312
rect 34940 18300 34946 18352
rect 35710 18300 35716 18352
rect 35768 18340 35774 18352
rect 38378 18340 38384 18352
rect 35768 18312 37320 18340
rect 38339 18312 38384 18340
rect 35768 18300 35774 18312
rect 22097 18275 22155 18281
rect 22097 18272 22109 18275
rect 21600 18244 22109 18272
rect 21600 18232 21606 18244
rect 22097 18241 22109 18244
rect 22143 18241 22155 18275
rect 22097 18235 22155 18241
rect 23017 18275 23075 18281
rect 23017 18241 23029 18275
rect 23063 18241 23075 18275
rect 23017 18235 23075 18241
rect 23106 18232 23112 18284
rect 23164 18272 23170 18284
rect 23273 18275 23331 18281
rect 23273 18272 23285 18275
rect 23164 18244 23285 18272
rect 23164 18232 23170 18244
rect 23273 18241 23285 18244
rect 23319 18241 23331 18275
rect 23273 18235 23331 18241
rect 23566 18232 23572 18284
rect 23624 18272 23630 18284
rect 24857 18275 24915 18281
rect 24857 18272 24869 18275
rect 23624 18244 24869 18272
rect 23624 18232 23630 18244
rect 24857 18241 24869 18244
rect 24903 18241 24915 18275
rect 24857 18235 24915 18241
rect 25682 18232 25688 18284
rect 25740 18272 25746 18284
rect 26050 18272 26056 18284
rect 25740 18244 26056 18272
rect 25740 18232 25746 18244
rect 26050 18232 26056 18244
rect 26108 18272 26114 18284
rect 26108 18244 26372 18272
rect 26108 18232 26114 18244
rect 20901 18207 20959 18213
rect 20901 18204 20913 18207
rect 20272 18176 20913 18204
rect 19521 18167 19579 18173
rect 20901 18173 20913 18176
rect 20947 18173 20959 18207
rect 20901 18167 20959 18173
rect 21821 18207 21879 18213
rect 21821 18173 21833 18207
rect 21867 18173 21879 18207
rect 26344 18204 26372 18244
rect 26418 18232 26424 18284
rect 26476 18272 26482 18284
rect 27157 18275 27215 18281
rect 27157 18272 27169 18275
rect 26476 18244 27169 18272
rect 26476 18232 26482 18244
rect 27157 18241 27169 18244
rect 27203 18241 27215 18275
rect 30190 18272 30196 18284
rect 30151 18244 30196 18272
rect 27157 18235 27215 18241
rect 30190 18232 30196 18244
rect 30248 18232 30254 18284
rect 32582 18232 32588 18284
rect 32640 18272 32646 18284
rect 32953 18275 33011 18281
rect 32953 18272 32965 18275
rect 32640 18244 32965 18272
rect 32640 18232 32646 18244
rect 32953 18241 32965 18244
rect 32999 18241 33011 18275
rect 32953 18235 33011 18241
rect 33045 18275 33103 18281
rect 33045 18241 33057 18275
rect 33091 18241 33103 18275
rect 33045 18235 33103 18241
rect 26970 18204 26976 18216
rect 26344 18176 26976 18204
rect 21821 18167 21879 18173
rect 20441 18139 20499 18145
rect 20441 18105 20453 18139
rect 20487 18136 20499 18139
rect 21836 18136 21864 18167
rect 26970 18164 26976 18176
rect 27028 18164 27034 18216
rect 28353 18207 28411 18213
rect 28353 18173 28365 18207
rect 28399 18173 28411 18207
rect 30466 18204 30472 18216
rect 30427 18176 30472 18204
rect 28353 18167 28411 18173
rect 26234 18136 26240 18148
rect 20487 18108 21864 18136
rect 26195 18108 26240 18136
rect 20487 18105 20499 18108
rect 20441 18099 20499 18105
rect 26234 18096 26240 18108
rect 26292 18096 26298 18148
rect 19426 18068 19432 18080
rect 17680 18040 19104 18068
rect 19387 18040 19432 18068
rect 19426 18028 19432 18040
rect 19484 18028 19490 18080
rect 21269 18071 21327 18077
rect 21269 18037 21281 18071
rect 21315 18068 21327 18071
rect 21913 18071 21971 18077
rect 21913 18068 21925 18071
rect 21315 18040 21925 18068
rect 21315 18037 21327 18040
rect 21269 18031 21327 18037
rect 21913 18037 21925 18040
rect 21959 18037 21971 18071
rect 21913 18031 21971 18037
rect 22281 18071 22339 18077
rect 22281 18037 22293 18071
rect 22327 18068 22339 18071
rect 23750 18068 23756 18080
rect 22327 18040 23756 18068
rect 22327 18037 22339 18040
rect 22281 18031 22339 18037
rect 23750 18028 23756 18040
rect 23808 18028 23814 18080
rect 24397 18071 24455 18077
rect 24397 18037 24409 18071
rect 24443 18068 24455 18071
rect 26418 18068 26424 18080
rect 24443 18040 26424 18068
rect 24443 18037 24455 18040
rect 24397 18031 24455 18037
rect 26418 18028 26424 18040
rect 26476 18028 26482 18080
rect 27433 18071 27491 18077
rect 27433 18037 27445 18071
rect 27479 18068 27491 18071
rect 27706 18068 27712 18080
rect 27479 18040 27712 18068
rect 27479 18037 27491 18040
rect 27433 18031 27491 18037
rect 27706 18028 27712 18040
rect 27764 18028 27770 18080
rect 28368 18068 28396 18167
rect 30466 18164 30472 18176
rect 30524 18164 30530 18216
rect 33060 18204 33088 18235
rect 33134 18232 33140 18284
rect 33192 18272 33198 18284
rect 34514 18272 34520 18284
rect 33192 18244 33237 18272
rect 34475 18244 34520 18272
rect 33192 18232 33198 18244
rect 34514 18232 34520 18244
rect 34572 18232 34578 18284
rect 34698 18281 34704 18284
rect 34665 18275 34704 18281
rect 34665 18241 34677 18275
rect 34665 18235 34704 18241
rect 34698 18232 34704 18235
rect 34756 18232 34762 18284
rect 34793 18275 34851 18281
rect 34793 18241 34805 18275
rect 34839 18241 34851 18275
rect 34793 18235 34851 18241
rect 33226 18204 33232 18216
rect 31726 18176 33232 18204
rect 31726 18136 31754 18176
rect 33226 18164 33232 18176
rect 33284 18164 33290 18216
rect 33321 18207 33379 18213
rect 33321 18173 33333 18207
rect 33367 18204 33379 18207
rect 34808 18204 34836 18235
rect 34974 18232 34980 18284
rect 35032 18281 35038 18284
rect 35032 18272 35040 18281
rect 35802 18272 35808 18284
rect 35032 18244 35077 18272
rect 35176 18244 35808 18272
rect 35032 18235 35040 18244
rect 35032 18232 35038 18235
rect 35176 18204 35204 18244
rect 35802 18232 35808 18244
rect 35860 18232 35866 18284
rect 35986 18272 35992 18284
rect 35947 18244 35992 18272
rect 35986 18232 35992 18244
rect 36044 18232 36050 18284
rect 37292 18281 37320 18312
rect 38378 18300 38384 18312
rect 38436 18300 38442 18352
rect 41386 18340 41414 18380
rect 43438 18368 43444 18380
rect 43496 18368 43502 18420
rect 41386 18312 43392 18340
rect 43364 18284 43392 18312
rect 37277 18275 37335 18281
rect 37277 18241 37289 18275
rect 37323 18241 37335 18275
rect 37458 18272 37464 18284
rect 37419 18244 37464 18272
rect 37277 18235 37335 18241
rect 37458 18232 37464 18244
rect 37516 18232 37522 18284
rect 43346 18272 43352 18284
rect 43307 18244 43352 18272
rect 43346 18232 43352 18244
rect 43404 18232 43410 18284
rect 33367 18176 35204 18204
rect 33367 18173 33379 18176
rect 33321 18167 33379 18173
rect 35250 18164 35256 18216
rect 35308 18204 35314 18216
rect 35897 18207 35955 18213
rect 35897 18204 35909 18207
rect 35308 18176 35909 18204
rect 35308 18164 35314 18176
rect 35897 18173 35909 18176
rect 35943 18173 35955 18207
rect 35897 18167 35955 18173
rect 38197 18207 38255 18213
rect 38197 18173 38209 18207
rect 38243 18204 38255 18207
rect 38746 18204 38752 18216
rect 38243 18176 38752 18204
rect 38243 18173 38255 18176
rect 38197 18167 38255 18173
rect 38746 18164 38752 18176
rect 38804 18164 38810 18216
rect 39942 18204 39948 18216
rect 39903 18176 39948 18204
rect 39942 18164 39948 18176
rect 40000 18164 40006 18216
rect 29288 18108 31754 18136
rect 28534 18068 28540 18080
rect 28368 18040 28540 18068
rect 28534 18028 28540 18040
rect 28592 18028 28598 18080
rect 28626 18028 28632 18080
rect 28684 18068 28690 18080
rect 29288 18068 29316 18108
rect 28684 18040 29316 18068
rect 29733 18071 29791 18077
rect 28684 18028 28690 18040
rect 29733 18037 29745 18071
rect 29779 18068 29791 18071
rect 30285 18071 30343 18077
rect 30285 18068 30297 18071
rect 29779 18040 30297 18068
rect 29779 18037 29791 18040
rect 29733 18031 29791 18037
rect 30285 18037 30297 18040
rect 30331 18037 30343 18071
rect 30285 18031 30343 18037
rect 30377 18071 30435 18077
rect 30377 18037 30389 18071
rect 30423 18068 30435 18071
rect 30650 18068 30656 18080
rect 30423 18040 30656 18068
rect 30423 18037 30435 18040
rect 30377 18031 30435 18037
rect 30650 18028 30656 18040
rect 30708 18028 30714 18080
rect 35161 18071 35219 18077
rect 35161 18037 35173 18071
rect 35207 18068 35219 18071
rect 35342 18068 35348 18080
rect 35207 18040 35348 18068
rect 35207 18037 35219 18040
rect 35161 18031 35219 18037
rect 35342 18028 35348 18040
rect 35400 18028 35406 18080
rect 36265 18071 36323 18077
rect 36265 18037 36277 18071
rect 36311 18068 36323 18071
rect 37274 18068 37280 18080
rect 36311 18040 37280 18068
rect 36311 18037 36323 18040
rect 36265 18031 36323 18037
rect 37274 18028 37280 18040
rect 37332 18028 37338 18080
rect 37458 18068 37464 18080
rect 37419 18040 37464 18068
rect 37458 18028 37464 18040
rect 37516 18028 37522 18080
rect 1104 17978 44896 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 44896 17978
rect 1104 17904 44896 17926
rect 2866 17864 2872 17876
rect 2827 17836 2872 17864
rect 2866 17824 2872 17836
rect 2924 17824 2930 17876
rect 16942 17824 16948 17876
rect 17000 17864 17006 17876
rect 17589 17867 17647 17873
rect 17589 17864 17601 17867
rect 17000 17836 17601 17864
rect 17000 17824 17006 17836
rect 17589 17833 17601 17836
rect 17635 17833 17647 17867
rect 17589 17827 17647 17833
rect 22189 17867 22247 17873
rect 22189 17833 22201 17867
rect 22235 17864 22247 17867
rect 23290 17864 23296 17876
rect 22235 17836 23296 17864
rect 22235 17833 22247 17836
rect 22189 17827 22247 17833
rect 23290 17824 23296 17836
rect 23348 17824 23354 17876
rect 26237 17867 26295 17873
rect 26237 17833 26249 17867
rect 26283 17864 26295 17867
rect 26418 17864 26424 17876
rect 26283 17836 26424 17864
rect 26283 17833 26295 17836
rect 26237 17827 26295 17833
rect 26418 17824 26424 17836
rect 26476 17864 26482 17876
rect 26789 17867 26847 17873
rect 26789 17864 26801 17867
rect 26476 17836 26801 17864
rect 26476 17824 26482 17836
rect 26789 17833 26801 17836
rect 26835 17833 26847 17867
rect 27893 17867 27951 17873
rect 27893 17864 27905 17867
rect 26789 17827 26847 17833
rect 27080 17836 27905 17864
rect 17310 17796 17316 17808
rect 15488 17768 17316 17796
rect 15488 17737 15516 17768
rect 17310 17756 17316 17768
rect 17368 17756 17374 17808
rect 25869 17799 25927 17805
rect 25869 17765 25881 17799
rect 25915 17796 25927 17799
rect 26694 17796 26700 17808
rect 25915 17768 26700 17796
rect 25915 17765 25927 17768
rect 25869 17759 25927 17765
rect 26694 17756 26700 17768
rect 26752 17756 26758 17808
rect 15473 17731 15531 17737
rect 15473 17697 15485 17731
rect 15519 17697 15531 17731
rect 15473 17691 15531 17697
rect 15562 17688 15568 17740
rect 15620 17728 15626 17740
rect 15620 17700 16252 17728
rect 15620 17688 15626 17700
rect 1762 17620 1768 17672
rect 1820 17660 1826 17672
rect 1857 17663 1915 17669
rect 1857 17660 1869 17663
rect 1820 17632 1869 17660
rect 1820 17620 1826 17632
rect 1857 17629 1869 17632
rect 1903 17629 1915 17663
rect 1857 17623 1915 17629
rect 2961 17663 3019 17669
rect 2961 17629 2973 17663
rect 3007 17660 3019 17663
rect 11698 17660 11704 17672
rect 3007 17632 11704 17660
rect 3007 17629 3019 17632
rect 2961 17623 3019 17629
rect 11698 17620 11704 17632
rect 11756 17620 11762 17672
rect 16224 17669 16252 17700
rect 17126 17688 17132 17740
rect 17184 17728 17190 17740
rect 17862 17728 17868 17740
rect 17184 17700 17868 17728
rect 17184 17688 17190 17700
rect 17862 17688 17868 17700
rect 17920 17688 17926 17740
rect 26234 17728 26240 17740
rect 26195 17700 26240 17728
rect 26234 17688 26240 17700
rect 26292 17688 26298 17740
rect 26881 17731 26939 17737
rect 26881 17697 26893 17731
rect 26927 17728 26939 17731
rect 26970 17728 26976 17740
rect 26927 17700 26976 17728
rect 26927 17697 26939 17700
rect 26881 17691 26939 17697
rect 26970 17688 26976 17700
rect 27028 17688 27034 17740
rect 15933 17663 15991 17669
rect 15933 17629 15945 17663
rect 15979 17629 15991 17663
rect 15933 17623 15991 17629
rect 16209 17663 16267 17669
rect 16209 17629 16221 17663
rect 16255 17660 16267 17663
rect 17034 17660 17040 17672
rect 16255 17632 17040 17660
rect 16255 17629 16267 17632
rect 16209 17623 16267 17629
rect 15194 17592 15200 17604
rect 15252 17601 15258 17604
rect 15164 17564 15200 17592
rect 15194 17552 15200 17564
rect 15252 17555 15264 17601
rect 15252 17552 15258 17555
rect 14093 17527 14151 17533
rect 14093 17493 14105 17527
rect 14139 17524 14151 17527
rect 15948 17524 15976 17623
rect 17034 17620 17040 17632
rect 17092 17620 17098 17672
rect 17494 17620 17500 17672
rect 17552 17660 17558 17672
rect 17589 17663 17647 17669
rect 17589 17660 17601 17663
rect 17552 17632 17601 17660
rect 17552 17620 17558 17632
rect 17589 17629 17601 17632
rect 17635 17629 17647 17663
rect 17589 17623 17647 17629
rect 17681 17663 17739 17669
rect 17681 17629 17693 17663
rect 17727 17629 17739 17663
rect 17681 17623 17739 17629
rect 19245 17663 19303 17669
rect 19245 17629 19257 17663
rect 19291 17660 19303 17663
rect 19426 17660 19432 17672
rect 19291 17632 19432 17660
rect 19291 17629 19303 17632
rect 19245 17623 19303 17629
rect 17402 17524 17408 17536
rect 14139 17496 17408 17524
rect 14139 17493 14151 17496
rect 14093 17487 14151 17493
rect 17402 17484 17408 17496
rect 17460 17524 17466 17536
rect 17696 17524 17724 17623
rect 19426 17620 19432 17632
rect 19484 17620 19490 17672
rect 19521 17663 19579 17669
rect 19521 17629 19533 17663
rect 19567 17629 19579 17663
rect 19521 17623 19579 17629
rect 19705 17663 19763 17669
rect 19705 17629 19717 17663
rect 19751 17660 19763 17663
rect 20346 17660 20352 17672
rect 19751 17632 20352 17660
rect 19751 17629 19763 17632
rect 19705 17623 19763 17629
rect 19536 17592 19564 17623
rect 20346 17620 20352 17632
rect 20404 17620 20410 17672
rect 20809 17663 20867 17669
rect 20809 17629 20821 17663
rect 20855 17660 20867 17663
rect 23474 17660 23480 17672
rect 20855 17632 23480 17660
rect 20855 17629 20867 17632
rect 20809 17623 20867 17629
rect 23474 17620 23480 17632
rect 23532 17620 23538 17672
rect 26050 17660 26056 17672
rect 26011 17632 26056 17660
rect 26050 17620 26056 17632
rect 26108 17620 26114 17672
rect 26252 17660 26280 17688
rect 26789 17663 26847 17669
rect 26789 17660 26801 17663
rect 26252 17632 26801 17660
rect 26789 17629 26801 17632
rect 26835 17629 26847 17663
rect 26789 17623 26847 17629
rect 21054 17595 21112 17601
rect 21054 17592 21066 17595
rect 19536 17564 21066 17592
rect 21054 17561 21066 17564
rect 21100 17561 21112 17595
rect 21054 17555 21112 17561
rect 24854 17552 24860 17604
rect 24912 17592 24918 17604
rect 25958 17592 25964 17604
rect 24912 17564 25964 17592
rect 24912 17552 24918 17564
rect 25958 17552 25964 17564
rect 26016 17592 26022 17604
rect 26329 17595 26387 17601
rect 26329 17592 26341 17595
rect 26016 17564 26341 17592
rect 26016 17552 26022 17564
rect 26329 17561 26341 17564
rect 26375 17592 26387 17595
rect 27080 17592 27108 17836
rect 27893 17833 27905 17836
rect 27939 17833 27951 17867
rect 27893 17827 27951 17833
rect 30466 17824 30472 17876
rect 30524 17864 30530 17876
rect 30929 17867 30987 17873
rect 30929 17864 30941 17867
rect 30524 17836 30941 17864
rect 30524 17824 30530 17836
rect 30929 17833 30941 17836
rect 30975 17833 30987 17867
rect 33134 17864 33140 17876
rect 30929 17827 30987 17833
rect 31726 17836 33140 17864
rect 28534 17756 28540 17808
rect 28592 17756 28598 17808
rect 28552 17728 28580 17756
rect 29546 17728 29552 17740
rect 28552 17700 29552 17728
rect 29546 17688 29552 17700
rect 29604 17688 29610 17740
rect 31726 17728 31754 17836
rect 33134 17824 33140 17836
rect 33192 17824 33198 17876
rect 34698 17824 34704 17876
rect 34756 17864 34762 17876
rect 35710 17864 35716 17876
rect 34756 17836 35716 17864
rect 34756 17824 34762 17836
rect 35710 17824 35716 17836
rect 35768 17824 35774 17876
rect 35986 17824 35992 17876
rect 36044 17864 36050 17876
rect 36173 17867 36231 17873
rect 36173 17864 36185 17867
rect 36044 17836 36185 17864
rect 36044 17824 36050 17836
rect 36173 17833 36185 17836
rect 36219 17833 36231 17867
rect 43622 17864 43628 17876
rect 36173 17827 36231 17833
rect 42444 17836 43628 17864
rect 32217 17799 32275 17805
rect 32217 17765 32229 17799
rect 32263 17796 32275 17799
rect 33318 17796 33324 17808
rect 32263 17768 33324 17796
rect 32263 17765 32275 17768
rect 32217 17759 32275 17765
rect 30576 17700 31754 17728
rect 27706 17620 27712 17672
rect 27764 17660 27770 17672
rect 28537 17663 28595 17669
rect 28537 17660 28549 17663
rect 27764 17632 28549 17660
rect 27764 17620 27770 17632
rect 28537 17629 28549 17632
rect 28583 17660 28595 17663
rect 28626 17660 28632 17672
rect 28583 17632 28632 17660
rect 28583 17629 28595 17632
rect 28537 17623 28595 17629
rect 28626 17620 28632 17632
rect 28684 17620 28690 17672
rect 28721 17663 28779 17669
rect 28721 17629 28733 17663
rect 28767 17660 28779 17663
rect 30576 17660 30604 17700
rect 32033 17663 32091 17669
rect 32033 17660 32045 17663
rect 28767 17632 30604 17660
rect 31726 17632 32045 17660
rect 28767 17629 28779 17632
rect 28721 17623 28779 17629
rect 28074 17592 28080 17604
rect 26375 17564 27108 17592
rect 27172 17564 27844 17592
rect 28035 17564 28080 17592
rect 26375 17561 26387 17564
rect 26329 17555 26387 17561
rect 17460 17496 17724 17524
rect 17957 17527 18015 17533
rect 17460 17484 17466 17496
rect 17957 17493 17969 17527
rect 18003 17524 18015 17527
rect 19337 17527 19395 17533
rect 19337 17524 19349 17527
rect 18003 17496 19349 17524
rect 18003 17493 18015 17496
rect 17957 17487 18015 17493
rect 19337 17493 19349 17496
rect 19383 17524 19395 17527
rect 19426 17524 19432 17536
rect 19383 17496 19432 17524
rect 19383 17493 19395 17496
rect 19337 17487 19395 17493
rect 19426 17484 19432 17496
rect 19484 17484 19490 17536
rect 27172 17533 27200 17564
rect 27157 17527 27215 17533
rect 27157 17493 27169 17527
rect 27203 17493 27215 17527
rect 27157 17487 27215 17493
rect 27246 17484 27252 17536
rect 27304 17524 27310 17536
rect 27709 17527 27767 17533
rect 27709 17524 27721 17527
rect 27304 17496 27721 17524
rect 27304 17484 27310 17496
rect 27709 17493 27721 17496
rect 27755 17493 27767 17527
rect 27816 17524 27844 17564
rect 28074 17552 28080 17564
rect 28132 17552 28138 17604
rect 28736 17592 28764 17623
rect 28644 17564 28764 17592
rect 27877 17527 27935 17533
rect 27877 17524 27889 17527
rect 27816 17496 27889 17524
rect 27709 17487 27767 17493
rect 27877 17493 27889 17496
rect 27923 17524 27935 17527
rect 28644 17524 28672 17564
rect 29454 17552 29460 17604
rect 29512 17592 29518 17604
rect 29794 17595 29852 17601
rect 29794 17592 29806 17595
rect 29512 17564 29806 17592
rect 29512 17552 29518 17564
rect 29794 17561 29806 17564
rect 29840 17561 29852 17595
rect 29794 17555 29852 17561
rect 30558 17552 30564 17604
rect 30616 17592 30622 17604
rect 31726 17592 31754 17632
rect 32033 17629 32045 17632
rect 32079 17629 32091 17663
rect 32033 17623 32091 17629
rect 30616 17564 31754 17592
rect 30616 17552 30622 17564
rect 27923 17496 28672 17524
rect 28721 17527 28779 17533
rect 27923 17493 27935 17496
rect 27877 17487 27935 17493
rect 28721 17493 28733 17527
rect 28767 17524 28779 17527
rect 28810 17524 28816 17536
rect 28767 17496 28816 17524
rect 28767 17493 28779 17496
rect 28721 17487 28779 17493
rect 28810 17484 28816 17496
rect 28868 17484 28874 17536
rect 31018 17484 31024 17536
rect 31076 17524 31082 17536
rect 32232 17524 32260 17759
rect 33318 17756 33324 17768
rect 33376 17756 33382 17808
rect 34532 17768 35480 17796
rect 34532 17740 34560 17768
rect 32582 17688 32588 17740
rect 32640 17728 32646 17740
rect 32769 17731 32827 17737
rect 32769 17728 32781 17731
rect 32640 17700 32781 17728
rect 32640 17688 32646 17700
rect 32769 17697 32781 17700
rect 32815 17697 32827 17731
rect 32769 17691 32827 17697
rect 32953 17731 33011 17737
rect 32953 17697 32965 17731
rect 32999 17728 33011 17731
rect 34514 17728 34520 17740
rect 32999 17700 34520 17728
rect 32999 17697 33011 17700
rect 32953 17691 33011 17697
rect 34514 17688 34520 17700
rect 34572 17688 34578 17740
rect 34790 17728 34796 17740
rect 34751 17700 34796 17728
rect 34790 17688 34796 17700
rect 34848 17688 34854 17740
rect 33226 17660 33232 17672
rect 33187 17632 33232 17660
rect 33226 17620 33232 17632
rect 33284 17620 33290 17672
rect 34606 17620 34612 17672
rect 34664 17660 34670 17672
rect 34882 17660 34888 17672
rect 34664 17632 34888 17660
rect 34664 17620 34670 17632
rect 34882 17620 34888 17632
rect 34940 17620 34946 17672
rect 35253 17663 35311 17669
rect 35253 17629 35265 17663
rect 35299 17660 35311 17663
rect 35342 17660 35348 17672
rect 35299 17632 35348 17660
rect 35299 17629 35311 17632
rect 35253 17623 35311 17629
rect 35342 17620 35348 17632
rect 35400 17620 35406 17672
rect 33134 17592 33140 17604
rect 33095 17564 33140 17592
rect 33134 17552 33140 17564
rect 33192 17552 33198 17604
rect 35161 17595 35219 17601
rect 35161 17561 35173 17595
rect 35207 17561 35219 17595
rect 35452 17592 35480 17768
rect 35728 17728 35756 17824
rect 36909 17731 36967 17737
rect 36909 17728 36921 17731
rect 35728 17700 36921 17728
rect 35728 17669 35756 17700
rect 36909 17697 36921 17700
rect 36955 17697 36967 17731
rect 36909 17691 36967 17697
rect 37369 17731 37427 17737
rect 37369 17697 37381 17731
rect 37415 17728 37427 17731
rect 38102 17728 38108 17740
rect 37415 17700 38108 17728
rect 37415 17697 37427 17700
rect 37369 17691 37427 17697
rect 38102 17688 38108 17700
rect 38160 17688 38166 17740
rect 42337 17731 42395 17737
rect 42337 17697 42349 17731
rect 42383 17728 42395 17731
rect 42444 17728 42472 17836
rect 43622 17824 43628 17836
rect 43680 17824 43686 17876
rect 42610 17756 42616 17808
rect 42668 17796 42674 17808
rect 42668 17768 43116 17796
rect 42668 17756 42674 17768
rect 42383 17700 42472 17728
rect 42521 17731 42579 17737
rect 42383 17697 42395 17700
rect 42337 17691 42395 17697
rect 42521 17697 42533 17731
rect 42567 17728 42579 17731
rect 42978 17728 42984 17740
rect 42567 17700 42984 17728
rect 42567 17697 42579 17700
rect 42521 17691 42579 17697
rect 42978 17688 42984 17700
rect 43036 17688 43042 17740
rect 43088 17737 43116 17768
rect 43073 17731 43131 17737
rect 43073 17697 43085 17731
rect 43119 17697 43131 17731
rect 43073 17691 43131 17697
rect 35713 17663 35771 17669
rect 35713 17629 35725 17663
rect 35759 17629 35771 17663
rect 35713 17623 35771 17629
rect 35802 17620 35808 17672
rect 35860 17660 35866 17672
rect 35989 17663 36047 17669
rect 35860 17632 35905 17660
rect 35860 17620 35866 17632
rect 35989 17629 36001 17663
rect 36035 17629 36047 17663
rect 36998 17660 37004 17672
rect 36959 17632 37004 17660
rect 35989 17623 36047 17629
rect 36004 17592 36032 17623
rect 36998 17620 37004 17632
rect 37056 17620 37062 17672
rect 35452 17564 36032 17592
rect 35161 17555 35219 17561
rect 31076 17496 32260 17524
rect 35176 17524 35204 17555
rect 35728 17536 35756 17564
rect 42978 17552 42984 17604
rect 43036 17592 43042 17604
rect 43162 17592 43168 17604
rect 43036 17564 43168 17592
rect 43036 17552 43042 17564
rect 43162 17552 43168 17564
rect 43220 17552 43226 17604
rect 35342 17524 35348 17536
rect 35176 17496 35348 17524
rect 31076 17484 31082 17496
rect 35342 17484 35348 17496
rect 35400 17484 35406 17536
rect 35710 17484 35716 17536
rect 35768 17484 35774 17536
rect 1104 17434 44896 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 44896 17434
rect 1104 17360 44896 17382
rect 15194 17280 15200 17332
rect 15252 17320 15258 17332
rect 15289 17323 15347 17329
rect 15289 17320 15301 17323
rect 15252 17292 15301 17320
rect 15252 17280 15258 17292
rect 15289 17289 15301 17292
rect 15335 17289 15347 17323
rect 15289 17283 15347 17289
rect 16960 17292 17264 17320
rect 14737 17255 14795 17261
rect 14737 17221 14749 17255
rect 14783 17252 14795 17255
rect 16960 17252 16988 17292
rect 14783 17224 16988 17252
rect 17037 17255 17095 17261
rect 14783 17221 14795 17224
rect 14737 17215 14795 17221
rect 17037 17221 17049 17255
rect 17083 17252 17095 17255
rect 17083 17224 17172 17252
rect 17083 17221 17095 17224
rect 17037 17215 17095 17221
rect 17144 17196 17172 17224
rect 1762 17184 1768 17196
rect 1723 17156 1768 17184
rect 1762 17144 1768 17156
rect 1820 17144 1826 17196
rect 14458 17144 14464 17196
rect 14516 17184 14522 17196
rect 14645 17187 14703 17193
rect 14645 17184 14657 17187
rect 14516 17156 14657 17184
rect 14516 17144 14522 17156
rect 14645 17153 14657 17156
rect 14691 17153 14703 17187
rect 14645 17147 14703 17153
rect 14829 17187 14887 17193
rect 14829 17153 14841 17187
rect 14875 17184 14887 17187
rect 15562 17184 15568 17196
rect 14875 17156 15568 17184
rect 14875 17153 14887 17156
rect 14829 17147 14887 17153
rect 1946 17116 1952 17128
rect 1907 17088 1952 17116
rect 1946 17076 1952 17088
rect 2004 17076 2010 17128
rect 2774 17116 2780 17128
rect 2735 17088 2780 17116
rect 2774 17076 2780 17088
rect 2832 17076 2838 17128
rect 14660 17048 14688 17147
rect 15562 17144 15568 17156
rect 15620 17144 15626 17196
rect 15657 17187 15715 17193
rect 15657 17153 15669 17187
rect 15703 17153 15715 17187
rect 15657 17147 15715 17153
rect 15749 17187 15807 17193
rect 15749 17153 15761 17187
rect 15795 17153 15807 17187
rect 15749 17147 15807 17153
rect 15933 17187 15991 17193
rect 15933 17153 15945 17187
rect 15979 17184 15991 17187
rect 16206 17184 16212 17196
rect 15979 17156 16212 17184
rect 15979 17153 15991 17156
rect 15933 17147 15991 17153
rect 15672 17048 15700 17147
rect 15764 17116 15792 17147
rect 16206 17144 16212 17156
rect 16264 17144 16270 17196
rect 16758 17144 16764 17196
rect 16816 17184 16822 17196
rect 16853 17187 16911 17193
rect 16853 17184 16865 17187
rect 16816 17156 16865 17184
rect 16816 17144 16822 17156
rect 16853 17153 16865 17156
rect 16899 17153 16911 17187
rect 16853 17147 16911 17153
rect 16942 17144 16948 17196
rect 17000 17184 17006 17196
rect 17000 17156 17045 17184
rect 17000 17144 17006 17156
rect 17126 17144 17132 17196
rect 17184 17144 17190 17196
rect 17236 17193 17264 17292
rect 17402 17280 17408 17332
rect 17460 17320 17466 17332
rect 20622 17320 20628 17332
rect 17460 17292 20628 17320
rect 17460 17280 17466 17292
rect 20622 17280 20628 17292
rect 20680 17280 20686 17332
rect 23290 17280 23296 17332
rect 23348 17320 23354 17332
rect 24854 17320 24860 17332
rect 23348 17292 24716 17320
rect 24815 17292 24860 17320
rect 23348 17280 23354 17292
rect 23750 17261 23756 17264
rect 23744 17252 23756 17261
rect 19444 17224 20484 17252
rect 23711 17224 23756 17252
rect 19444 17196 19472 17224
rect 17221 17187 17279 17193
rect 17221 17153 17233 17187
rect 17267 17153 17279 17187
rect 17221 17147 17279 17153
rect 17494 17144 17500 17196
rect 17552 17184 17558 17196
rect 17681 17187 17739 17193
rect 17681 17184 17693 17187
rect 17552 17156 17693 17184
rect 17552 17144 17558 17156
rect 17681 17153 17693 17156
rect 17727 17153 17739 17187
rect 17681 17147 17739 17153
rect 17773 17187 17831 17193
rect 17773 17153 17785 17187
rect 17819 17184 17831 17187
rect 19426 17184 19432 17196
rect 17819 17156 18276 17184
rect 19387 17156 19432 17184
rect 17819 17153 17831 17156
rect 17773 17147 17831 17153
rect 17788 17116 17816 17147
rect 15764 17088 16712 17116
rect 16684 17057 16712 17088
rect 16776 17088 17816 17116
rect 14660 17020 15700 17048
rect 16669 17051 16727 17057
rect 16669 17017 16681 17051
rect 16715 17017 16727 17051
rect 16669 17011 16727 17017
rect 15286 16940 15292 16992
rect 15344 16980 15350 16992
rect 16776 16980 16804 17088
rect 17862 17076 17868 17128
rect 17920 17116 17926 17128
rect 18141 17119 18199 17125
rect 18141 17116 18153 17119
rect 17920 17088 18153 17116
rect 17920 17076 17926 17088
rect 18141 17085 18153 17088
rect 18187 17085 18199 17119
rect 18248 17116 18276 17156
rect 19426 17144 19432 17156
rect 19484 17144 19490 17196
rect 19610 17184 19616 17196
rect 19571 17156 19616 17184
rect 19610 17144 19616 17156
rect 19668 17184 19674 17196
rect 20070 17184 20076 17196
rect 19668 17156 20076 17184
rect 19668 17144 19674 17156
rect 20070 17144 20076 17156
rect 20128 17144 20134 17196
rect 20456 17193 20484 17224
rect 23744 17215 23756 17224
rect 23750 17212 23756 17215
rect 23808 17212 23814 17264
rect 20441 17187 20499 17193
rect 20441 17153 20453 17187
rect 20487 17184 20499 17187
rect 20530 17184 20536 17196
rect 20487 17156 20536 17184
rect 20487 17153 20499 17156
rect 20441 17147 20499 17153
rect 20530 17144 20536 17156
rect 20588 17144 20594 17196
rect 21818 17184 21824 17196
rect 21779 17156 21824 17184
rect 21818 17144 21824 17156
rect 21876 17144 21882 17196
rect 22005 17187 22063 17193
rect 22005 17153 22017 17187
rect 22051 17184 22063 17187
rect 22738 17184 22744 17196
rect 22051 17156 22744 17184
rect 22051 17153 22063 17156
rect 22005 17147 22063 17153
rect 22738 17144 22744 17156
rect 22796 17144 22802 17196
rect 19337 17119 19395 17125
rect 19337 17116 19349 17119
rect 18248 17088 19349 17116
rect 18141 17079 18199 17085
rect 19337 17085 19349 17088
rect 19383 17116 19395 17119
rect 19518 17116 19524 17128
rect 19383 17088 19524 17116
rect 19383 17085 19395 17088
rect 19337 17079 19395 17085
rect 19518 17076 19524 17088
rect 19576 17116 19582 17128
rect 20257 17119 20315 17125
rect 20257 17116 20269 17119
rect 19576 17088 20269 17116
rect 19576 17076 19582 17088
rect 20257 17085 20269 17088
rect 20303 17085 20315 17119
rect 20257 17079 20315 17085
rect 20346 17076 20352 17128
rect 20404 17116 20410 17128
rect 23290 17116 23296 17128
rect 20404 17088 23296 17116
rect 20404 17076 20410 17088
rect 23290 17076 23296 17088
rect 23348 17076 23354 17128
rect 23474 17116 23480 17128
rect 23387 17088 23480 17116
rect 23474 17076 23480 17088
rect 23532 17076 23538 17128
rect 24688 17116 24716 17292
rect 24854 17280 24860 17292
rect 24912 17280 24918 17332
rect 29638 17320 29644 17332
rect 25332 17292 29644 17320
rect 25332 17264 25360 17292
rect 29638 17280 29644 17292
rect 29696 17280 29702 17332
rect 29917 17323 29975 17329
rect 29917 17289 29929 17323
rect 29963 17320 29975 17323
rect 30190 17320 30196 17332
rect 29963 17292 30196 17320
rect 29963 17289 29975 17292
rect 29917 17283 29975 17289
rect 30190 17280 30196 17292
rect 30248 17280 30254 17332
rect 30558 17320 30564 17332
rect 30519 17292 30564 17320
rect 30558 17280 30564 17292
rect 30616 17280 30622 17332
rect 25314 17252 25320 17264
rect 25275 17224 25320 17252
rect 25314 17212 25320 17224
rect 25372 17212 25378 17264
rect 25501 17255 25559 17261
rect 25501 17221 25513 17255
rect 25547 17252 25559 17255
rect 27614 17252 27620 17264
rect 25547 17224 27620 17252
rect 25547 17221 25559 17224
rect 25501 17215 25559 17221
rect 27614 17212 27620 17224
rect 27672 17212 27678 17264
rect 29454 17212 29460 17264
rect 29512 17252 29518 17264
rect 34882 17252 34888 17264
rect 29512 17224 34888 17252
rect 29512 17212 29518 17224
rect 34882 17212 34888 17224
rect 34940 17212 34946 17264
rect 35710 17212 35716 17264
rect 35768 17252 35774 17264
rect 35805 17255 35863 17261
rect 35805 17252 35817 17255
rect 35768 17224 35817 17252
rect 35768 17212 35774 17224
rect 35805 17221 35817 17224
rect 35851 17221 35863 17255
rect 35805 17215 35863 17221
rect 24762 17144 24768 17196
rect 24820 17184 24826 17196
rect 26053 17187 26111 17193
rect 26053 17184 26065 17187
rect 24820 17156 26065 17184
rect 24820 17144 24826 17156
rect 26053 17153 26065 17156
rect 26099 17153 26111 17187
rect 27157 17187 27215 17193
rect 27157 17184 27169 17187
rect 26053 17147 26111 17153
rect 26160 17156 27169 17184
rect 26160 17116 26188 17156
rect 27157 17153 27169 17156
rect 27203 17184 27215 17187
rect 28074 17184 28080 17196
rect 27203 17156 28080 17184
rect 27203 17153 27215 17156
rect 27157 17147 27215 17153
rect 28074 17144 28080 17156
rect 28132 17144 28138 17196
rect 28810 17193 28816 17196
rect 28804 17184 28816 17193
rect 28771 17156 28816 17184
rect 28804 17147 28816 17156
rect 28810 17144 28816 17147
rect 28868 17144 28874 17196
rect 29730 17144 29736 17196
rect 29788 17184 29794 17196
rect 30469 17187 30527 17193
rect 30469 17184 30481 17187
rect 29788 17156 30481 17184
rect 29788 17144 29794 17156
rect 30469 17153 30481 17156
rect 30515 17153 30527 17187
rect 32858 17184 32864 17196
rect 32819 17156 32864 17184
rect 30469 17147 30527 17153
rect 32858 17144 32864 17156
rect 32916 17144 32922 17196
rect 33042 17184 33048 17196
rect 33003 17156 33048 17184
rect 33042 17144 33048 17156
rect 33100 17144 33106 17196
rect 36998 17184 37004 17196
rect 36280 17156 37004 17184
rect 27062 17116 27068 17128
rect 24688 17088 26188 17116
rect 27023 17088 27068 17116
rect 27062 17076 27068 17088
rect 27120 17076 27126 17128
rect 28534 17116 28540 17128
rect 28495 17088 28540 17116
rect 28534 17076 28540 17088
rect 28592 17076 28598 17128
rect 36280 17125 36308 17156
rect 36998 17144 37004 17156
rect 37056 17184 37062 17196
rect 37277 17187 37335 17193
rect 37277 17184 37289 17187
rect 37056 17156 37289 17184
rect 37056 17144 37062 17156
rect 37277 17153 37289 17156
rect 37323 17153 37335 17187
rect 37458 17184 37464 17196
rect 37419 17156 37464 17184
rect 37277 17147 37335 17153
rect 37458 17144 37464 17156
rect 37516 17144 37522 17196
rect 42978 17144 42984 17196
rect 43036 17184 43042 17196
rect 43349 17187 43407 17193
rect 43349 17184 43361 17187
rect 43036 17156 43361 17184
rect 43036 17144 43042 17156
rect 43349 17153 43361 17156
rect 43395 17153 43407 17187
rect 43349 17147 43407 17153
rect 36265 17119 36323 17125
rect 36265 17085 36277 17119
rect 36311 17085 36323 17119
rect 36265 17079 36323 17085
rect 19797 17051 19855 17057
rect 19797 17017 19809 17051
rect 19843 17048 19855 17051
rect 21174 17048 21180 17060
rect 19843 17020 21180 17048
rect 19843 17017 19855 17020
rect 19797 17011 19855 17017
rect 21174 17008 21180 17020
rect 21232 17008 21238 17060
rect 15344 16952 16804 16980
rect 15344 16940 15350 16952
rect 16942 16940 16948 16992
rect 17000 16980 17006 16992
rect 17957 16983 18015 16989
rect 17957 16980 17969 16983
rect 17000 16952 17969 16980
rect 17000 16940 17006 16952
rect 17957 16949 17969 16952
rect 18003 16949 18015 16983
rect 17957 16943 18015 16949
rect 20254 16940 20260 16992
rect 20312 16980 20318 16992
rect 20625 16983 20683 16989
rect 20625 16980 20637 16983
rect 20312 16952 20637 16980
rect 20312 16940 20318 16952
rect 20625 16949 20637 16952
rect 20671 16949 20683 16983
rect 22002 16980 22008 16992
rect 21963 16952 22008 16980
rect 20625 16943 20683 16949
rect 22002 16940 22008 16952
rect 22060 16940 22066 16992
rect 23492 16980 23520 17076
rect 26237 17051 26295 17057
rect 26237 17017 26249 17051
rect 26283 17048 26295 17051
rect 26326 17048 26332 17060
rect 26283 17020 26332 17048
rect 26283 17017 26295 17020
rect 26237 17011 26295 17017
rect 26326 17008 26332 17020
rect 26384 17008 26390 17060
rect 27525 17051 27583 17057
rect 27525 17017 27537 17051
rect 27571 17048 27583 17051
rect 27614 17048 27620 17060
rect 27571 17020 27620 17048
rect 27571 17017 27583 17020
rect 27525 17011 27583 17017
rect 27614 17008 27620 17020
rect 27672 17008 27678 17060
rect 35894 17008 35900 17060
rect 35952 17048 35958 17060
rect 36081 17051 36139 17057
rect 36081 17048 36093 17051
rect 35952 17020 36093 17048
rect 35952 17008 35958 17020
rect 36081 17017 36093 17020
rect 36127 17017 36139 17051
rect 36081 17011 36139 17017
rect 23842 16980 23848 16992
rect 23492 16952 23848 16980
rect 23842 16940 23848 16952
rect 23900 16940 23906 16992
rect 32953 16983 33011 16989
rect 32953 16949 32965 16983
rect 32999 16980 33011 16983
rect 33778 16980 33784 16992
rect 32999 16952 33784 16980
rect 32999 16949 33011 16952
rect 32953 16943 33011 16949
rect 33778 16940 33784 16952
rect 33836 16940 33842 16992
rect 37645 16983 37703 16989
rect 37645 16949 37657 16983
rect 37691 16980 37703 16983
rect 38930 16980 38936 16992
rect 37691 16952 38936 16980
rect 37691 16949 37703 16952
rect 37645 16943 37703 16949
rect 38930 16940 38936 16952
rect 38988 16940 38994 16992
rect 43441 16983 43499 16989
rect 43441 16949 43453 16983
rect 43487 16980 43499 16983
rect 43990 16980 43996 16992
rect 43487 16952 43996 16980
rect 43487 16949 43499 16952
rect 43441 16943 43499 16949
rect 43990 16940 43996 16952
rect 44048 16940 44054 16992
rect 44174 16980 44180 16992
rect 44135 16952 44180 16980
rect 44174 16940 44180 16952
rect 44232 16940 44238 16992
rect 1104 16890 44896 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 44896 16890
rect 1104 16816 44896 16838
rect 1946 16736 1952 16788
rect 2004 16776 2010 16788
rect 2317 16779 2375 16785
rect 2317 16776 2329 16779
rect 2004 16748 2329 16776
rect 2004 16736 2010 16748
rect 2317 16745 2329 16748
rect 2363 16745 2375 16779
rect 15746 16776 15752 16788
rect 15707 16748 15752 16776
rect 2317 16739 2375 16745
rect 15746 16736 15752 16748
rect 15804 16736 15810 16788
rect 16022 16736 16028 16788
rect 16080 16776 16086 16788
rect 16666 16776 16672 16788
rect 16080 16748 16672 16776
rect 16080 16736 16086 16748
rect 16666 16736 16672 16748
rect 16724 16776 16730 16788
rect 17494 16776 17500 16788
rect 16724 16748 17500 16776
rect 16724 16736 16730 16748
rect 17494 16736 17500 16748
rect 17552 16736 17558 16788
rect 23106 16776 23112 16788
rect 23067 16748 23112 16776
rect 23106 16736 23112 16748
rect 23164 16736 23170 16788
rect 15838 16708 15844 16720
rect 15396 16680 15844 16708
rect 6178 16640 6184 16652
rect 2424 16612 6184 16640
rect 1670 16532 1676 16584
rect 1728 16572 1734 16584
rect 2424 16581 2452 16612
rect 6178 16600 6184 16612
rect 6236 16600 6242 16652
rect 15286 16640 15292 16652
rect 15247 16612 15292 16640
rect 15286 16600 15292 16612
rect 15344 16600 15350 16652
rect 15396 16649 15424 16680
rect 15838 16668 15844 16680
rect 15896 16668 15902 16720
rect 20806 16708 20812 16720
rect 20767 16680 20812 16708
rect 20806 16668 20812 16680
rect 20864 16668 20870 16720
rect 22738 16708 22744 16720
rect 22699 16680 22744 16708
rect 22738 16668 22744 16680
rect 22796 16668 22802 16720
rect 23290 16668 23296 16720
rect 23348 16708 23354 16720
rect 32401 16711 32459 16717
rect 23348 16680 24900 16708
rect 23348 16668 23354 16680
rect 15381 16643 15439 16649
rect 15381 16609 15393 16643
rect 15427 16609 15439 16643
rect 15381 16603 15439 16609
rect 15473 16643 15531 16649
rect 15473 16609 15485 16643
rect 15519 16640 15531 16643
rect 15930 16640 15936 16652
rect 15519 16612 15936 16640
rect 15519 16609 15531 16612
rect 15473 16603 15531 16609
rect 15930 16600 15936 16612
rect 15988 16600 15994 16652
rect 17310 16640 17316 16652
rect 16224 16612 17080 16640
rect 17271 16612 17316 16640
rect 1765 16575 1823 16581
rect 1765 16572 1777 16575
rect 1728 16544 1777 16572
rect 1728 16532 1734 16544
rect 1765 16541 1777 16544
rect 1811 16541 1823 16575
rect 1765 16535 1823 16541
rect 2409 16575 2467 16581
rect 2409 16541 2421 16575
rect 2455 16574 2467 16575
rect 13449 16575 13507 16581
rect 2455 16546 2489 16574
rect 2455 16541 2467 16546
rect 2409 16535 2467 16541
rect 13449 16541 13461 16575
rect 13495 16572 13507 16575
rect 15565 16575 15623 16581
rect 13495 16544 15148 16572
rect 13495 16541 13507 16544
rect 13449 16535 13507 16541
rect 12894 16396 12900 16448
rect 12952 16436 12958 16448
rect 13265 16439 13323 16445
rect 13265 16436 13277 16439
rect 12952 16408 13277 16436
rect 12952 16396 12958 16408
rect 13265 16405 13277 16408
rect 13311 16405 13323 16439
rect 15120 16436 15148 16544
rect 15565 16541 15577 16575
rect 15611 16572 15623 16575
rect 16022 16572 16028 16584
rect 15611 16544 16028 16572
rect 15611 16541 15623 16544
rect 15565 16535 15623 16541
rect 16022 16532 16028 16544
rect 16080 16532 16086 16584
rect 16224 16581 16252 16612
rect 16209 16575 16267 16581
rect 16209 16541 16221 16575
rect 16255 16541 16267 16575
rect 16209 16535 16267 16541
rect 16393 16575 16451 16581
rect 16393 16541 16405 16575
rect 16439 16541 16451 16575
rect 16393 16535 16451 16541
rect 16485 16575 16543 16581
rect 16485 16541 16497 16575
rect 16531 16541 16543 16575
rect 16485 16535 16543 16541
rect 16577 16575 16635 16581
rect 16577 16541 16589 16575
rect 16623 16572 16635 16575
rect 16666 16572 16672 16584
rect 16623 16544 16672 16572
rect 16623 16541 16635 16544
rect 16577 16535 16635 16541
rect 15746 16464 15752 16516
rect 15804 16504 15810 16516
rect 16408 16504 16436 16535
rect 15804 16476 16436 16504
rect 16500 16504 16528 16535
rect 16666 16532 16672 16544
rect 16724 16532 16730 16584
rect 16942 16572 16948 16584
rect 16776 16544 16948 16572
rect 16776 16504 16804 16544
rect 16942 16532 16948 16544
rect 17000 16532 17006 16584
rect 17052 16572 17080 16612
rect 17310 16600 17316 16612
rect 17368 16600 17374 16652
rect 19518 16640 19524 16652
rect 19479 16612 19524 16640
rect 19518 16600 19524 16612
rect 19576 16600 19582 16652
rect 20990 16600 20996 16652
rect 21048 16640 21054 16652
rect 21453 16643 21511 16649
rect 21453 16640 21465 16643
rect 21048 16612 21465 16640
rect 21048 16600 21054 16612
rect 21453 16609 21465 16612
rect 21499 16640 21511 16643
rect 23934 16640 23940 16652
rect 21499 16612 23940 16640
rect 21499 16609 21511 16612
rect 21453 16603 21511 16609
rect 23934 16600 23940 16612
rect 23992 16600 23998 16652
rect 24762 16640 24768 16652
rect 24044 16612 24768 16640
rect 17402 16572 17408 16584
rect 17052 16544 17408 16572
rect 17402 16532 17408 16544
rect 17460 16532 17466 16584
rect 19242 16572 19248 16584
rect 19203 16544 19248 16572
rect 19242 16532 19248 16544
rect 19300 16532 19306 16584
rect 21634 16572 21640 16584
rect 21595 16544 21640 16572
rect 21634 16532 21640 16544
rect 21692 16532 21698 16584
rect 16500 16476 16804 16504
rect 16853 16507 16911 16513
rect 15804 16464 15810 16476
rect 16853 16473 16865 16507
rect 16899 16504 16911 16507
rect 17558 16507 17616 16513
rect 17558 16504 17570 16507
rect 16899 16476 17570 16504
rect 16899 16473 16911 16476
rect 16853 16467 16911 16473
rect 17558 16473 17570 16476
rect 17604 16473 17616 16507
rect 17558 16467 17616 16473
rect 17678 16464 17684 16516
rect 17736 16504 17742 16516
rect 19610 16504 19616 16516
rect 17736 16476 19616 16504
rect 17736 16464 17742 16476
rect 19610 16464 19616 16476
rect 19668 16504 19674 16516
rect 20533 16507 20591 16513
rect 20533 16504 20545 16507
rect 19668 16476 20545 16504
rect 19668 16464 19674 16476
rect 20533 16473 20545 16476
rect 20579 16473 20591 16507
rect 20533 16467 20591 16473
rect 22186 16464 22192 16516
rect 22244 16504 22250 16516
rect 23109 16507 23167 16513
rect 23109 16504 23121 16507
rect 22244 16476 23121 16504
rect 22244 16464 22250 16476
rect 23109 16473 23121 16476
rect 23155 16473 23167 16507
rect 24044 16504 24072 16612
rect 24762 16600 24768 16612
rect 24820 16600 24826 16652
rect 24872 16649 24900 16680
rect 32401 16677 32413 16711
rect 32447 16708 32459 16711
rect 33042 16708 33048 16720
rect 32447 16680 33048 16708
rect 32447 16677 32459 16680
rect 32401 16671 32459 16677
rect 33042 16668 33048 16680
rect 33100 16668 33106 16720
rect 37093 16711 37151 16717
rect 33888 16680 35020 16708
rect 24857 16643 24915 16649
rect 24857 16609 24869 16643
rect 24903 16609 24915 16643
rect 31018 16640 31024 16652
rect 30979 16612 31024 16640
rect 24857 16603 24915 16609
rect 31018 16600 31024 16612
rect 31076 16600 31082 16652
rect 33778 16640 33784 16652
rect 33739 16612 33784 16640
rect 33778 16600 33784 16612
rect 33836 16600 33842 16652
rect 33888 16649 33916 16680
rect 33873 16643 33931 16649
rect 33873 16609 33885 16643
rect 33919 16609 33931 16643
rect 34054 16640 34060 16652
rect 34015 16612 34060 16640
rect 33873 16603 33931 16609
rect 34054 16600 34060 16612
rect 34112 16600 34118 16652
rect 34992 16649 35020 16680
rect 37093 16677 37105 16711
rect 37139 16677 37151 16711
rect 37093 16671 37151 16677
rect 34977 16643 35035 16649
rect 34977 16609 34989 16643
rect 35023 16640 35035 16643
rect 35342 16640 35348 16652
rect 35023 16612 35348 16640
rect 35023 16609 35035 16612
rect 34977 16603 35035 16609
rect 35342 16600 35348 16612
rect 35400 16600 35406 16652
rect 37108 16640 37136 16671
rect 37458 16640 37464 16652
rect 37108 16612 37464 16640
rect 37458 16600 37464 16612
rect 37516 16640 37522 16652
rect 37645 16643 37703 16649
rect 37645 16640 37657 16643
rect 37516 16612 37657 16640
rect 37516 16600 37522 16612
rect 37645 16609 37657 16612
rect 37691 16609 37703 16643
rect 43990 16640 43996 16652
rect 43951 16612 43996 16640
rect 37645 16603 37703 16609
rect 43990 16600 43996 16612
rect 44048 16600 44054 16652
rect 44174 16640 44180 16652
rect 44135 16612 44180 16640
rect 44174 16600 44180 16612
rect 44232 16600 44238 16652
rect 34888 16584 34940 16590
rect 24394 16572 24400 16584
rect 24355 16544 24400 16572
rect 24394 16532 24400 16544
rect 24452 16532 24458 16584
rect 24673 16575 24731 16581
rect 24673 16541 24685 16575
rect 24719 16572 24731 16575
rect 24946 16572 24952 16584
rect 24719 16544 24952 16572
rect 24719 16541 24731 16544
rect 24673 16535 24731 16541
rect 24946 16532 24952 16544
rect 25004 16532 25010 16584
rect 30742 16532 30748 16584
rect 30800 16572 30806 16584
rect 31277 16575 31335 16581
rect 31277 16572 31289 16575
rect 30800 16544 31289 16572
rect 30800 16532 30806 16544
rect 31277 16541 31289 16544
rect 31323 16541 31335 16575
rect 31277 16535 31335 16541
rect 36725 16575 36783 16581
rect 36725 16541 36737 16575
rect 36771 16572 36783 16575
rect 36998 16572 37004 16584
rect 36771 16544 37004 16572
rect 36771 16541 36783 16544
rect 36725 16535 36783 16541
rect 36998 16532 37004 16544
rect 37056 16532 37062 16584
rect 37918 16572 37924 16584
rect 37879 16544 37924 16572
rect 37918 16532 37924 16544
rect 37976 16532 37982 16584
rect 42334 16572 42340 16584
rect 42295 16544 42340 16572
rect 42334 16532 42340 16544
rect 42392 16532 42398 16584
rect 34888 16526 34940 16532
rect 23109 16467 23167 16473
rect 23308 16476 24072 16504
rect 18046 16436 18052 16448
rect 15120 16408 18052 16436
rect 13265 16399 13323 16405
rect 18046 16396 18052 16408
rect 18104 16396 18110 16448
rect 18690 16436 18696 16448
rect 18603 16408 18696 16436
rect 18690 16396 18696 16408
rect 18748 16436 18754 16448
rect 19242 16436 19248 16448
rect 18748 16408 19248 16436
rect 18748 16396 18754 16408
rect 19242 16396 19248 16408
rect 19300 16396 19306 16448
rect 20993 16439 21051 16445
rect 20993 16405 21005 16439
rect 21039 16436 21051 16439
rect 21082 16436 21088 16448
rect 21039 16408 21088 16436
rect 21039 16405 21051 16408
rect 20993 16399 21051 16405
rect 21082 16396 21088 16408
rect 21140 16396 21146 16448
rect 23308 16445 23336 16476
rect 32950 16464 32956 16516
rect 33008 16504 33014 16516
rect 35802 16504 35808 16516
rect 33008 16476 34836 16504
rect 35763 16476 35808 16504
rect 33008 16464 33014 16476
rect 23293 16439 23351 16445
rect 23293 16405 23305 16439
rect 23339 16405 23351 16439
rect 23293 16399 23351 16405
rect 23474 16396 23480 16448
rect 23532 16436 23538 16448
rect 24489 16439 24547 16445
rect 24489 16436 24501 16439
rect 23532 16408 24501 16436
rect 23532 16396 23538 16408
rect 24489 16405 24501 16408
rect 24535 16405 24547 16439
rect 24489 16399 24547 16405
rect 33226 16396 33232 16448
rect 33284 16436 33290 16448
rect 33413 16439 33471 16445
rect 33413 16436 33425 16439
rect 33284 16408 33425 16436
rect 33284 16396 33290 16408
rect 33413 16405 33425 16408
rect 33459 16405 33471 16439
rect 34808 16436 34836 16476
rect 35802 16464 35808 16476
rect 35860 16464 35866 16516
rect 40126 16504 40132 16516
rect 37108 16476 40132 16504
rect 37108 16436 37136 16476
rect 40126 16464 40132 16476
rect 40184 16464 40190 16516
rect 34808 16408 37136 16436
rect 37185 16439 37243 16445
rect 33413 16399 33471 16405
rect 37185 16405 37197 16439
rect 37231 16436 37243 16439
rect 37274 16436 37280 16448
rect 37231 16408 37280 16436
rect 37231 16405 37243 16408
rect 37185 16399 37243 16405
rect 37274 16396 37280 16408
rect 37332 16396 37338 16448
rect 1104 16346 44896 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 44896 16346
rect 1104 16272 44896 16294
rect 15654 16192 15660 16244
rect 15712 16232 15718 16244
rect 17678 16232 17684 16244
rect 15712 16204 17684 16232
rect 15712 16192 15718 16204
rect 17678 16192 17684 16204
rect 17736 16192 17742 16244
rect 17862 16232 17868 16244
rect 17823 16204 17868 16232
rect 17862 16192 17868 16204
rect 17920 16192 17926 16244
rect 22281 16235 22339 16241
rect 20456 16204 21588 16232
rect 16758 16124 16764 16176
rect 16816 16164 16822 16176
rect 19521 16167 19579 16173
rect 16816 16136 16905 16164
rect 16816 16124 16822 16136
rect 1670 16096 1676 16108
rect 1631 16068 1676 16096
rect 1670 16056 1676 16068
rect 1728 16056 1734 16108
rect 12894 16096 12900 16108
rect 12855 16068 12900 16096
rect 12894 16056 12900 16068
rect 12952 16056 12958 16108
rect 15286 16056 15292 16108
rect 15344 16096 15350 16108
rect 15749 16099 15807 16105
rect 15749 16096 15761 16099
rect 15344 16068 15761 16096
rect 15344 16056 15350 16068
rect 15749 16065 15761 16068
rect 15795 16065 15807 16099
rect 15749 16059 15807 16065
rect 15933 16099 15991 16105
rect 15933 16065 15945 16099
rect 15979 16096 15991 16099
rect 16022 16096 16028 16108
rect 15979 16068 16028 16096
rect 15979 16065 15991 16068
rect 15933 16059 15991 16065
rect 16022 16056 16028 16068
rect 16080 16056 16086 16108
rect 16877 16105 16905 16136
rect 19521 16133 19533 16167
rect 19567 16133 19579 16167
rect 19521 16127 19579 16133
rect 16877 16099 16957 16105
rect 16877 16068 16911 16099
rect 16899 16065 16911 16068
rect 16945 16065 16957 16099
rect 16899 16059 16957 16065
rect 17037 16099 17095 16105
rect 17037 16065 17049 16099
rect 17083 16065 17095 16099
rect 17037 16059 17095 16065
rect 1857 16031 1915 16037
rect 1857 15997 1869 16031
rect 1903 16028 1915 16031
rect 2222 16028 2228 16040
rect 1903 16000 2228 16028
rect 1903 15997 1915 16000
rect 1857 15991 1915 15997
rect 2222 15988 2228 16000
rect 2280 15988 2286 16040
rect 2774 16028 2780 16040
rect 2735 16000 2780 16028
rect 2774 15988 2780 16000
rect 2832 15988 2838 16040
rect 13081 16031 13139 16037
rect 13081 15997 13093 16031
rect 13127 16028 13139 16031
rect 13170 16028 13176 16040
rect 13127 16000 13176 16028
rect 13127 15997 13139 16000
rect 13081 15991 13139 15997
rect 13170 15988 13176 16000
rect 13228 15988 13234 16040
rect 14734 16028 14740 16040
rect 14695 16000 14740 16028
rect 14734 15988 14740 16000
rect 14792 15988 14798 16040
rect 15654 16028 15660 16040
rect 15615 16000 15660 16028
rect 15654 15988 15660 16000
rect 15712 15988 15718 16040
rect 15838 16028 15844 16040
rect 15799 16000 15844 16028
rect 15838 15988 15844 16000
rect 15896 15988 15902 16040
rect 16666 15988 16672 16040
rect 16724 16028 16730 16040
rect 17052 16028 17080 16059
rect 17126 16056 17132 16108
rect 17184 16099 17190 16108
rect 17313 16099 17371 16105
rect 17184 16071 17226 16099
rect 17184 16056 17190 16071
rect 17313 16065 17325 16099
rect 17359 16096 17371 16099
rect 17402 16096 17408 16108
rect 17359 16068 17408 16096
rect 17359 16065 17371 16068
rect 17313 16059 17371 16065
rect 17402 16056 17408 16068
rect 17460 16056 17466 16108
rect 17586 16056 17592 16108
rect 17644 16096 17650 16108
rect 17865 16099 17923 16105
rect 17865 16096 17877 16099
rect 17644 16068 17877 16096
rect 17644 16056 17650 16068
rect 17865 16065 17877 16068
rect 17911 16065 17923 16099
rect 17865 16059 17923 16065
rect 18141 16099 18199 16105
rect 18141 16065 18153 16099
rect 18187 16096 18199 16099
rect 18506 16096 18512 16108
rect 18187 16068 18512 16096
rect 18187 16065 18199 16068
rect 18141 16059 18199 16065
rect 16724 16000 17080 16028
rect 16724 15988 16730 16000
rect 16942 15960 16948 15972
rect 16132 15932 16948 15960
rect 3418 15852 3424 15904
rect 3476 15892 3482 15904
rect 12526 15892 12532 15904
rect 3476 15864 12532 15892
rect 3476 15852 3482 15864
rect 12526 15852 12532 15864
rect 12584 15852 12590 15904
rect 16132 15901 16160 15932
rect 16942 15920 16948 15932
rect 17000 15920 17006 15972
rect 16117 15895 16175 15901
rect 16117 15861 16129 15895
rect 16163 15861 16175 15895
rect 16117 15855 16175 15861
rect 16574 15852 16580 15904
rect 16632 15892 16638 15904
rect 16669 15895 16727 15901
rect 16669 15892 16681 15895
rect 16632 15864 16681 15892
rect 16632 15852 16638 15864
rect 16669 15861 16681 15864
rect 16715 15861 16727 15895
rect 16669 15855 16727 15861
rect 16758 15852 16764 15904
rect 16816 15892 16822 15904
rect 18156 15892 18184 16059
rect 18506 16056 18512 16068
rect 18564 16056 18570 16108
rect 19334 15960 19340 15972
rect 19295 15932 19340 15960
rect 19334 15920 19340 15932
rect 19392 15920 19398 15972
rect 19536 15960 19564 16127
rect 20254 16096 20260 16108
rect 20215 16068 20260 16096
rect 20254 16056 20260 16068
rect 20312 16056 20318 16108
rect 20456 16105 20484 16204
rect 21560 16176 21588 16204
rect 22281 16201 22293 16235
rect 22327 16232 22339 16235
rect 22370 16232 22376 16244
rect 22327 16204 22376 16232
rect 22327 16201 22339 16204
rect 22281 16195 22339 16201
rect 22370 16192 22376 16204
rect 22428 16192 22434 16244
rect 23477 16235 23535 16241
rect 23477 16201 23489 16235
rect 23523 16232 23535 16235
rect 32950 16232 32956 16244
rect 23523 16204 32956 16232
rect 23523 16201 23535 16204
rect 23477 16195 23535 16201
rect 32950 16192 32956 16204
rect 33008 16192 33014 16244
rect 33226 16232 33232 16244
rect 33187 16204 33232 16232
rect 33226 16192 33232 16204
rect 33284 16192 33290 16244
rect 33873 16235 33931 16241
rect 33873 16201 33885 16235
rect 33919 16232 33931 16235
rect 34882 16232 34888 16244
rect 33919 16204 34888 16232
rect 33919 16201 33931 16204
rect 33873 16195 33931 16201
rect 34882 16192 34888 16204
rect 34940 16192 34946 16244
rect 21542 16124 21548 16176
rect 21600 16164 21606 16176
rect 23293 16167 23351 16173
rect 21600 16136 22140 16164
rect 21600 16124 21606 16136
rect 20441 16099 20499 16105
rect 20441 16065 20453 16099
rect 20487 16065 20499 16099
rect 20806 16096 20812 16108
rect 20441 16059 20499 16065
rect 20548 16068 20812 16096
rect 20165 16031 20223 16037
rect 20165 15997 20177 16031
rect 20211 16028 20223 16031
rect 20548 16028 20576 16068
rect 20806 16056 20812 16068
rect 20864 16056 20870 16108
rect 21821 16099 21879 16105
rect 21821 16065 21833 16099
rect 21867 16096 21879 16099
rect 22002 16096 22008 16108
rect 21867 16068 22008 16096
rect 21867 16065 21879 16068
rect 21821 16059 21879 16065
rect 22002 16056 22008 16068
rect 22060 16056 22066 16108
rect 22112 16105 22140 16136
rect 23293 16133 23305 16167
rect 23339 16164 23351 16167
rect 26510 16164 26516 16176
rect 23339 16136 26516 16164
rect 23339 16133 23351 16136
rect 23293 16127 23351 16133
rect 26510 16124 26516 16136
rect 26568 16124 26574 16176
rect 27614 16124 27620 16176
rect 27672 16164 27678 16176
rect 28804 16167 28862 16173
rect 28804 16164 28816 16167
rect 27672 16136 28816 16164
rect 27672 16124 27678 16136
rect 28804 16133 28816 16136
rect 28850 16164 28862 16167
rect 32858 16164 32864 16176
rect 28850 16136 32864 16164
rect 28850 16133 28862 16136
rect 28804 16127 28862 16133
rect 32858 16124 32864 16136
rect 32916 16124 32922 16176
rect 33042 16164 33048 16176
rect 33003 16136 33048 16164
rect 33042 16124 33048 16136
rect 33100 16124 33106 16176
rect 22097 16099 22155 16105
rect 22097 16065 22109 16099
rect 22143 16065 22155 16099
rect 24193 16099 24251 16105
rect 24193 16096 24205 16099
rect 22097 16059 22155 16065
rect 23124 16068 24205 16096
rect 20211 16000 20576 16028
rect 20625 16031 20683 16037
rect 20211 15997 20223 16000
rect 20165 15991 20223 15997
rect 20625 15997 20637 16031
rect 20671 16028 20683 16031
rect 23124 16028 23152 16068
rect 24193 16065 24205 16068
rect 24239 16065 24251 16099
rect 24193 16059 24251 16065
rect 26973 16099 27031 16105
rect 26973 16065 26985 16099
rect 27019 16065 27031 16099
rect 26973 16059 27031 16065
rect 20671 16000 23152 16028
rect 20671 15997 20683 16000
rect 20625 15991 20683 15997
rect 23842 15988 23848 16040
rect 23900 16028 23906 16040
rect 23937 16031 23995 16037
rect 23937 16028 23949 16031
rect 23900 16000 23949 16028
rect 23900 15988 23906 16000
rect 23937 15997 23949 16000
rect 23983 15997 23995 16031
rect 23937 15991 23995 15997
rect 20990 15960 20996 15972
rect 19536 15932 20996 15960
rect 20990 15920 20996 15932
rect 21048 15920 21054 15972
rect 21082 15920 21088 15972
rect 21140 15960 21146 15972
rect 22925 15963 22983 15969
rect 22925 15960 22937 15963
rect 21140 15932 22937 15960
rect 21140 15920 21146 15932
rect 22925 15929 22937 15932
rect 22971 15929 22983 15963
rect 22925 15923 22983 15929
rect 25317 15963 25375 15969
rect 25317 15929 25329 15963
rect 25363 15960 25375 15963
rect 26234 15960 26240 15972
rect 25363 15932 26240 15960
rect 25363 15929 25375 15932
rect 25317 15923 25375 15929
rect 26234 15920 26240 15932
rect 26292 15960 26298 15972
rect 26988 15960 27016 16059
rect 27062 16056 27068 16108
rect 27120 16096 27126 16108
rect 27157 16099 27215 16105
rect 27157 16096 27169 16099
rect 27120 16068 27169 16096
rect 27120 16056 27126 16068
rect 27157 16065 27169 16068
rect 27203 16096 27215 16099
rect 27246 16096 27252 16108
rect 27203 16068 27252 16096
rect 27203 16065 27215 16068
rect 27157 16059 27215 16065
rect 27246 16056 27252 16068
rect 27304 16056 27310 16108
rect 27801 16099 27859 16105
rect 27801 16065 27813 16099
rect 27847 16065 27859 16099
rect 28534 16096 28540 16108
rect 28495 16068 28540 16096
rect 27801 16059 27859 16065
rect 26292 15932 27016 15960
rect 26292 15920 26298 15932
rect 16816 15864 18184 15892
rect 16816 15852 16822 15864
rect 21634 15852 21640 15904
rect 21692 15892 21698 15904
rect 21913 15895 21971 15901
rect 21913 15892 21925 15895
rect 21692 15864 21925 15892
rect 21692 15852 21698 15864
rect 21913 15861 21925 15864
rect 21959 15861 21971 15895
rect 21913 15855 21971 15861
rect 22554 15852 22560 15904
rect 22612 15892 22618 15904
rect 23293 15895 23351 15901
rect 23293 15892 23305 15895
rect 22612 15864 23305 15892
rect 22612 15852 22618 15864
rect 23293 15861 23305 15864
rect 23339 15892 23351 15895
rect 23474 15892 23480 15904
rect 23339 15864 23480 15892
rect 23339 15861 23351 15864
rect 23293 15855 23351 15861
rect 23474 15852 23480 15864
rect 23532 15852 23538 15904
rect 27062 15852 27068 15904
rect 27120 15892 27126 15904
rect 27157 15895 27215 15901
rect 27157 15892 27169 15895
rect 27120 15864 27169 15892
rect 27120 15852 27126 15864
rect 27157 15861 27169 15864
rect 27203 15861 27215 15895
rect 27614 15892 27620 15904
rect 27575 15864 27620 15892
rect 27157 15855 27215 15861
rect 27614 15852 27620 15864
rect 27672 15852 27678 15904
rect 27816 15892 27844 16059
rect 28534 16056 28540 16068
rect 28592 16056 28598 16108
rect 33244 16096 33272 16192
rect 37366 16124 37372 16176
rect 37424 16164 37430 16176
rect 37424 16136 37780 16164
rect 37424 16124 37430 16136
rect 33689 16099 33747 16105
rect 33689 16096 33701 16099
rect 33244 16068 33701 16096
rect 33689 16065 33701 16068
rect 33735 16065 33747 16099
rect 33689 16059 33747 16065
rect 33778 16056 33784 16108
rect 33836 16096 33842 16108
rect 33873 16099 33931 16105
rect 33873 16096 33885 16099
rect 33836 16068 33885 16096
rect 33836 16056 33842 16068
rect 33873 16065 33885 16068
rect 33919 16065 33931 16099
rect 33873 16059 33931 16065
rect 35802 16056 35808 16108
rect 35860 16096 35866 16108
rect 37752 16105 37780 16136
rect 36541 16099 36599 16105
rect 36541 16096 36553 16099
rect 35860 16068 36553 16096
rect 35860 16056 35866 16068
rect 36541 16065 36553 16068
rect 36587 16065 36599 16099
rect 36541 16059 36599 16065
rect 36725 16099 36783 16105
rect 36725 16065 36737 16099
rect 36771 16096 36783 16099
rect 37737 16099 37795 16105
rect 36771 16068 37596 16096
rect 36771 16065 36783 16068
rect 36725 16059 36783 16065
rect 36262 15988 36268 16040
rect 36320 16028 36326 16040
rect 36740 16028 36768 16059
rect 36320 16000 36768 16028
rect 36320 15988 36326 16000
rect 37568 15969 37596 16068
rect 37737 16065 37749 16099
rect 37783 16065 37795 16099
rect 38102 16096 38108 16108
rect 38063 16068 38108 16096
rect 37737 16059 37795 16065
rect 38102 16056 38108 16068
rect 38160 16056 38166 16108
rect 43254 16056 43260 16108
rect 43312 16096 43318 16108
rect 43349 16099 43407 16105
rect 43349 16096 43361 16099
rect 43312 16068 43361 16096
rect 43312 16056 43318 16068
rect 43349 16065 43361 16068
rect 43395 16065 43407 16099
rect 43349 16059 43407 16065
rect 37553 15963 37611 15969
rect 37553 15929 37565 15963
rect 37599 15929 37611 15963
rect 37553 15923 37611 15929
rect 29546 15892 29552 15904
rect 27816 15864 29552 15892
rect 29546 15852 29552 15864
rect 29604 15852 29610 15904
rect 29914 15892 29920 15904
rect 29875 15864 29920 15892
rect 29914 15852 29920 15864
rect 29972 15852 29978 15904
rect 36725 15895 36783 15901
rect 36725 15861 36737 15895
rect 36771 15892 36783 15895
rect 37458 15892 37464 15904
rect 36771 15864 37464 15892
rect 36771 15861 36783 15864
rect 36725 15855 36783 15861
rect 37458 15852 37464 15864
rect 37516 15852 37522 15904
rect 37918 15892 37924 15904
rect 37879 15864 37924 15892
rect 37918 15852 37924 15864
rect 37976 15852 37982 15904
rect 42702 15892 42708 15904
rect 42663 15864 42708 15892
rect 42702 15852 42708 15864
rect 42760 15852 42766 15904
rect 43438 15892 43444 15904
rect 43399 15864 43444 15892
rect 43438 15852 43444 15864
rect 43496 15852 43502 15904
rect 44174 15892 44180 15904
rect 44135 15864 44180 15892
rect 44174 15852 44180 15864
rect 44232 15852 44238 15904
rect 1104 15802 44896 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 44896 15802
rect 1104 15728 44896 15750
rect 2222 15688 2228 15700
rect 2183 15660 2228 15688
rect 2222 15648 2228 15660
rect 2280 15648 2286 15700
rect 13170 15688 13176 15700
rect 13131 15660 13176 15688
rect 13170 15648 13176 15660
rect 13228 15648 13234 15700
rect 15289 15691 15347 15697
rect 15289 15657 15301 15691
rect 15335 15688 15347 15691
rect 15654 15688 15660 15700
rect 15335 15660 15660 15688
rect 15335 15657 15347 15660
rect 15289 15651 15347 15657
rect 15654 15648 15660 15660
rect 15712 15648 15718 15700
rect 15930 15648 15936 15700
rect 15988 15688 15994 15700
rect 16666 15688 16672 15700
rect 15988 15660 16672 15688
rect 15988 15648 15994 15660
rect 16666 15648 16672 15660
rect 16724 15688 16730 15700
rect 17221 15691 17279 15697
rect 17221 15688 17233 15691
rect 16724 15660 17233 15688
rect 16724 15648 16730 15660
rect 17221 15657 17233 15660
rect 17267 15657 17279 15691
rect 17221 15651 17279 15657
rect 19705 15691 19763 15697
rect 19705 15657 19717 15691
rect 19751 15688 19763 15691
rect 19978 15688 19984 15700
rect 19751 15660 19984 15688
rect 19751 15657 19763 15660
rect 19705 15651 19763 15657
rect 19978 15648 19984 15660
rect 20036 15648 20042 15700
rect 20533 15691 20591 15697
rect 20533 15657 20545 15691
rect 20579 15688 20591 15691
rect 20806 15688 20812 15700
rect 20579 15660 20812 15688
rect 20579 15657 20591 15660
rect 20533 15651 20591 15657
rect 20806 15648 20812 15660
rect 20864 15648 20870 15700
rect 21174 15688 21180 15700
rect 21135 15660 21180 15688
rect 21174 15648 21180 15660
rect 21232 15648 21238 15700
rect 22186 15688 22192 15700
rect 22147 15660 22192 15688
rect 22186 15648 22192 15660
rect 22244 15648 22250 15700
rect 22554 15688 22560 15700
rect 22515 15660 22560 15688
rect 22554 15648 22560 15660
rect 22612 15648 22618 15700
rect 22738 15648 22744 15700
rect 22796 15688 22802 15700
rect 26510 15688 26516 15700
rect 22796 15660 23152 15688
rect 26471 15660 26516 15688
rect 22796 15648 22802 15660
rect 17310 15620 17316 15632
rect 16684 15592 17316 15620
rect 16684 15564 16712 15592
rect 17310 15580 17316 15592
rect 17368 15580 17374 15632
rect 21818 15580 21824 15632
rect 21876 15620 21882 15632
rect 23124 15629 23152 15660
rect 26510 15648 26516 15660
rect 26568 15648 26574 15700
rect 23109 15623 23167 15629
rect 21876 15592 23060 15620
rect 21876 15580 21882 15592
rect 16666 15512 16672 15564
rect 16724 15552 16730 15564
rect 21082 15552 21088 15564
rect 16724 15524 16817 15552
rect 21043 15524 21088 15552
rect 16724 15512 16730 15524
rect 21082 15512 21088 15524
rect 21140 15512 21146 15564
rect 21542 15552 21548 15564
rect 21376 15524 21548 15552
rect 2317 15487 2375 15493
rect 2317 15453 2329 15487
rect 2363 15484 2375 15487
rect 2406 15484 2412 15496
rect 2363 15456 2412 15484
rect 2363 15453 2375 15456
rect 2317 15447 2375 15453
rect 2406 15444 2412 15456
rect 2464 15484 2470 15496
rect 3418 15484 3424 15496
rect 2464 15456 3424 15484
rect 2464 15444 2470 15456
rect 3418 15444 3424 15456
rect 3476 15444 3482 15496
rect 13265 15487 13323 15493
rect 13265 15453 13277 15487
rect 13311 15484 13323 15487
rect 13538 15484 13544 15496
rect 13311 15456 13544 15484
rect 13311 15453 13323 15456
rect 13265 15447 13323 15453
rect 13538 15444 13544 15456
rect 13596 15444 13602 15496
rect 16413 15487 16471 15493
rect 16413 15453 16425 15487
rect 16459 15484 16471 15487
rect 16574 15484 16580 15496
rect 16459 15456 16580 15484
rect 16459 15453 16471 15456
rect 16413 15447 16471 15453
rect 16574 15444 16580 15456
rect 16632 15444 16638 15496
rect 17313 15487 17371 15493
rect 17313 15453 17325 15487
rect 17359 15484 17371 15487
rect 17586 15484 17592 15496
rect 17359 15456 17592 15484
rect 17359 15453 17371 15456
rect 17313 15447 17371 15453
rect 17586 15444 17592 15456
rect 17644 15444 17650 15496
rect 19242 15444 19248 15496
rect 19300 15484 19306 15496
rect 20349 15487 20407 15493
rect 20349 15484 20361 15487
rect 19300 15456 20361 15484
rect 19300 15444 19306 15456
rect 20349 15453 20361 15456
rect 20395 15453 20407 15487
rect 20530 15484 20536 15496
rect 20491 15456 20536 15484
rect 20349 15447 20407 15453
rect 20530 15444 20536 15456
rect 20588 15444 20594 15496
rect 21376 15493 21404 15524
rect 21542 15512 21548 15524
rect 21600 15512 21606 15564
rect 22922 15552 22928 15564
rect 22204 15524 22928 15552
rect 22204 15493 22232 15524
rect 22922 15512 22928 15524
rect 22980 15512 22986 15564
rect 21361 15487 21419 15493
rect 21361 15453 21373 15487
rect 21407 15453 21419 15487
rect 21361 15447 21419 15453
rect 22189 15487 22247 15493
rect 22189 15453 22201 15487
rect 22235 15453 22247 15487
rect 22189 15447 22247 15453
rect 22278 15444 22284 15496
rect 22336 15484 22342 15496
rect 23032 15493 23060 15592
rect 23109 15589 23121 15623
rect 23155 15589 23167 15623
rect 36078 15620 36084 15632
rect 36039 15592 36084 15620
rect 23109 15583 23167 15589
rect 36078 15580 36084 15592
rect 36136 15580 36142 15632
rect 23290 15552 23296 15564
rect 23251 15524 23296 15552
rect 23290 15512 23296 15524
rect 23348 15512 23354 15564
rect 36280 15524 37322 15552
rect 23017 15487 23075 15493
rect 22336 15456 22381 15484
rect 22336 15444 22342 15456
rect 23017 15453 23029 15487
rect 23063 15453 23075 15487
rect 23017 15447 23075 15453
rect 24397 15487 24455 15493
rect 24397 15453 24409 15487
rect 24443 15484 24455 15487
rect 27893 15487 27951 15493
rect 27893 15484 27905 15487
rect 24443 15456 27905 15484
rect 24443 15453 24455 15456
rect 24397 15447 24455 15453
rect 27540 15428 27568 15456
rect 27893 15453 27905 15456
rect 27939 15453 27951 15487
rect 29638 15484 29644 15496
rect 29599 15456 29644 15484
rect 27893 15447 27951 15453
rect 29638 15444 29644 15456
rect 29696 15444 29702 15496
rect 30929 15487 30987 15493
rect 30929 15453 30941 15487
rect 30975 15484 30987 15487
rect 31018 15484 31024 15496
rect 30975 15456 31024 15484
rect 30975 15453 30987 15456
rect 30929 15447 30987 15453
rect 31018 15444 31024 15456
rect 31076 15444 31082 15496
rect 31202 15493 31208 15496
rect 31196 15484 31208 15493
rect 31163 15456 31208 15484
rect 31196 15447 31208 15456
rect 31202 15444 31208 15447
rect 31260 15444 31266 15496
rect 32769 15487 32827 15493
rect 32769 15484 32781 15487
rect 32324 15456 32781 15484
rect 19797 15419 19855 15425
rect 19797 15416 19809 15419
rect 19260 15388 19809 15416
rect 19260 15360 19288 15388
rect 19797 15385 19809 15388
rect 19843 15385 19855 15419
rect 19797 15379 19855 15385
rect 21545 15419 21603 15425
rect 21545 15385 21557 15419
rect 21591 15416 21603 15419
rect 24642 15419 24700 15425
rect 24642 15416 24654 15419
rect 21591 15388 24654 15416
rect 21591 15385 21603 15388
rect 21545 15379 21603 15385
rect 24642 15385 24654 15388
rect 24688 15385 24700 15419
rect 24642 15379 24700 15385
rect 27522 15376 27528 15428
rect 27580 15376 27586 15428
rect 27614 15376 27620 15428
rect 27672 15425 27678 15428
rect 27672 15416 27684 15425
rect 27672 15388 27717 15416
rect 27672 15379 27684 15388
rect 27672 15376 27678 15379
rect 32324 15360 32352 15456
rect 32769 15453 32781 15456
rect 32815 15453 32827 15487
rect 32950 15484 32956 15496
rect 32911 15456 32956 15484
rect 32769 15447 32827 15453
rect 32950 15444 32956 15456
rect 33008 15444 33014 15496
rect 33226 15444 33232 15496
rect 33284 15484 33290 15496
rect 33597 15487 33655 15493
rect 33597 15484 33609 15487
rect 33284 15456 33609 15484
rect 33284 15444 33290 15456
rect 33597 15453 33609 15456
rect 33643 15453 33655 15487
rect 33597 15447 33655 15453
rect 33781 15487 33839 15493
rect 33781 15453 33793 15487
rect 33827 15453 33839 15487
rect 33781 15447 33839 15453
rect 33796 15416 33824 15447
rect 35802 15444 35808 15496
rect 35860 15484 35866 15496
rect 36280 15493 36308 15524
rect 36081 15487 36139 15493
rect 36081 15484 36093 15487
rect 35860 15456 36093 15484
rect 35860 15444 35866 15456
rect 36081 15453 36093 15456
rect 36127 15453 36139 15487
rect 36081 15447 36139 15453
rect 36265 15487 36323 15493
rect 36265 15453 36277 15487
rect 36311 15453 36323 15487
rect 36265 15447 36323 15453
rect 36357 15487 36415 15493
rect 36357 15453 36369 15487
rect 36403 15484 36415 15487
rect 37294 15484 37322 15524
rect 37366 15512 37372 15564
rect 37424 15552 37430 15564
rect 37645 15555 37703 15561
rect 37645 15552 37657 15555
rect 37424 15524 37657 15552
rect 37424 15512 37430 15524
rect 37645 15521 37657 15524
rect 37691 15521 37703 15555
rect 42610 15552 42616 15564
rect 42571 15524 42616 15552
rect 37645 15515 37703 15521
rect 42610 15512 42616 15524
rect 42668 15512 42674 15564
rect 44174 15552 44180 15564
rect 44135 15524 44180 15552
rect 44174 15512 44180 15524
rect 44232 15512 44238 15564
rect 37734 15484 37740 15496
rect 36403 15456 37228 15484
rect 37294 15456 37740 15484
rect 36403 15453 36415 15456
rect 36357 15447 36415 15453
rect 37200 15425 37228 15456
rect 37734 15444 37740 15456
rect 37792 15484 37798 15496
rect 37921 15487 37979 15493
rect 37921 15484 37933 15487
rect 37792 15456 37933 15484
rect 37792 15444 37798 15456
rect 37921 15453 37933 15456
rect 37967 15453 37979 15487
rect 38930 15484 38936 15496
rect 38891 15456 38936 15484
rect 37921 15447 37979 15453
rect 38930 15444 38936 15456
rect 38988 15444 38994 15496
rect 33152 15388 33824 15416
rect 37001 15419 37059 15425
rect 33152 15360 33180 15388
rect 37001 15385 37013 15419
rect 37047 15385 37059 15419
rect 37001 15379 37059 15385
rect 37185 15419 37243 15425
rect 37185 15385 37197 15419
rect 37231 15416 37243 15419
rect 37274 15416 37280 15428
rect 37231 15388 37280 15416
rect 37231 15385 37243 15388
rect 37185 15379 37243 15385
rect 19242 15308 19248 15360
rect 19300 15308 19306 15360
rect 23293 15351 23351 15357
rect 23293 15317 23305 15351
rect 23339 15348 23351 15351
rect 24394 15348 24400 15360
rect 23339 15320 24400 15348
rect 23339 15317 23351 15320
rect 23293 15311 23351 15317
rect 24394 15308 24400 15320
rect 24452 15308 24458 15360
rect 25777 15351 25835 15357
rect 25777 15317 25789 15351
rect 25823 15348 25835 15351
rect 25958 15348 25964 15360
rect 25823 15320 25964 15348
rect 25823 15317 25835 15320
rect 25777 15311 25835 15317
rect 25958 15308 25964 15320
rect 26016 15308 26022 15360
rect 29730 15348 29736 15360
rect 29691 15320 29736 15348
rect 29730 15308 29736 15320
rect 29788 15308 29794 15360
rect 32306 15348 32312 15360
rect 32267 15320 32312 15348
rect 32306 15308 32312 15320
rect 32364 15308 32370 15360
rect 33134 15348 33140 15360
rect 33095 15320 33140 15348
rect 33134 15308 33140 15320
rect 33192 15308 33198 15360
rect 33594 15308 33600 15360
rect 33652 15348 33658 15360
rect 33689 15351 33747 15357
rect 33689 15348 33701 15351
rect 33652 15320 33701 15348
rect 33652 15308 33658 15320
rect 33689 15317 33701 15320
rect 33735 15317 33747 15351
rect 36814 15348 36820 15360
rect 36775 15320 36820 15348
rect 33689 15311 33747 15317
rect 36814 15308 36820 15320
rect 36872 15308 36878 15360
rect 37016 15348 37044 15379
rect 37274 15376 37280 15388
rect 37332 15376 37338 15428
rect 43990 15416 43996 15428
rect 43951 15388 43996 15416
rect 43990 15376 43996 15388
rect 44048 15376 44054 15428
rect 37366 15348 37372 15360
rect 37016 15320 37372 15348
rect 37366 15308 37372 15320
rect 37424 15308 37430 15360
rect 39022 15348 39028 15360
rect 38983 15320 39028 15348
rect 39022 15308 39028 15320
rect 39080 15308 39086 15360
rect 1104 15258 44896 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 44896 15258
rect 1104 15184 44896 15206
rect 15838 15104 15844 15156
rect 15896 15144 15902 15156
rect 17497 15147 17555 15153
rect 17497 15144 17509 15147
rect 15896 15116 17509 15144
rect 15896 15104 15902 15116
rect 17497 15113 17509 15116
rect 17543 15113 17555 15147
rect 17497 15107 17555 15113
rect 17665 15147 17723 15153
rect 17665 15113 17677 15147
rect 17711 15144 17723 15147
rect 18138 15144 18144 15156
rect 17711 15116 18144 15144
rect 17711 15113 17723 15116
rect 17665 15107 17723 15113
rect 18138 15104 18144 15116
rect 18196 15104 18202 15156
rect 23658 15104 23664 15156
rect 23716 15144 23722 15156
rect 25501 15147 25559 15153
rect 25501 15144 25513 15147
rect 23716 15116 25513 15144
rect 23716 15104 23722 15116
rect 25501 15113 25513 15116
rect 25547 15113 25559 15147
rect 25501 15107 25559 15113
rect 25884 15116 27292 15144
rect 17865 15079 17923 15085
rect 17865 15045 17877 15079
rect 17911 15076 17923 15079
rect 19058 15076 19064 15088
rect 17911 15048 19064 15076
rect 17911 15045 17923 15048
rect 17865 15039 17923 15045
rect 19058 15036 19064 15048
rect 19116 15036 19122 15088
rect 21174 15076 21180 15088
rect 21008 15048 21180 15076
rect 13357 15011 13415 15017
rect 13357 14977 13369 15011
rect 13403 15008 13415 15011
rect 13538 15008 13544 15020
rect 13403 14980 13544 15008
rect 13403 14977 13415 14980
rect 13357 14971 13415 14977
rect 13538 14968 13544 14980
rect 13596 14968 13602 15020
rect 18506 15008 18512 15020
rect 18467 14980 18512 15008
rect 18506 14968 18512 14980
rect 18564 14968 18570 15020
rect 19521 15011 19579 15017
rect 19521 14977 19533 15011
rect 19567 15008 19579 15011
rect 19978 15008 19984 15020
rect 19567 14980 19984 15008
rect 19567 14977 19579 14980
rect 19521 14971 19579 14977
rect 19978 14968 19984 14980
rect 20036 14968 20042 15020
rect 20809 15011 20867 15017
rect 20809 14977 20821 15011
rect 20855 15008 20867 15011
rect 20898 15008 20904 15020
rect 20855 14980 20904 15008
rect 20855 14977 20867 14980
rect 20809 14971 20867 14977
rect 20898 14968 20904 14980
rect 20956 14968 20962 15020
rect 21008 15017 21036 15048
rect 21174 15036 21180 15048
rect 21232 15076 21238 15088
rect 22738 15076 22744 15088
rect 21232 15048 22744 15076
rect 21232 15036 21238 15048
rect 22738 15036 22744 15048
rect 22796 15036 22802 15088
rect 22922 15036 22928 15088
rect 22980 15076 22986 15088
rect 23293 15079 23351 15085
rect 23293 15076 23305 15079
rect 22980 15048 23305 15076
rect 22980 15036 22986 15048
rect 23293 15045 23305 15048
rect 23339 15045 23351 15079
rect 23934 15076 23940 15088
rect 23895 15048 23940 15076
rect 23293 15039 23351 15045
rect 23934 15036 23940 15048
rect 23992 15036 23998 15088
rect 25409 15079 25467 15085
rect 25409 15045 25421 15079
rect 25455 15076 25467 15079
rect 25774 15076 25780 15088
rect 25455 15048 25780 15076
rect 25455 15045 25467 15048
rect 25409 15039 25467 15045
rect 25774 15036 25780 15048
rect 25832 15036 25838 15088
rect 20993 15011 21051 15017
rect 20993 14977 21005 15011
rect 21039 14977 21051 15011
rect 20993 14971 21051 14977
rect 21821 15011 21879 15017
rect 21821 14977 21833 15011
rect 21867 15008 21879 15011
rect 22186 15008 22192 15020
rect 21867 14980 22192 15008
rect 21867 14977 21879 14980
rect 21821 14971 21879 14977
rect 22186 14968 22192 14980
rect 22244 14968 22250 15020
rect 22756 15008 22784 15036
rect 23109 15011 23167 15017
rect 23109 15008 23121 15011
rect 22756 14980 23121 15008
rect 23109 14977 23121 14980
rect 23155 14977 23167 15011
rect 23109 14971 23167 14977
rect 24210 14968 24216 15020
rect 24268 15008 24274 15020
rect 25884 15008 25912 15116
rect 25958 15036 25964 15088
rect 26016 15076 26022 15088
rect 27264 15076 27292 15116
rect 29546 15104 29552 15156
rect 29604 15144 29610 15156
rect 30561 15147 30619 15153
rect 30561 15144 30573 15147
rect 29604 15116 30573 15144
rect 29604 15104 29610 15116
rect 30561 15113 30573 15116
rect 30607 15113 30619 15147
rect 35345 15147 35403 15153
rect 30561 15107 30619 15113
rect 30668 15116 34192 15144
rect 30668 15076 30696 15116
rect 26016 15048 27200 15076
rect 27264 15048 30696 15076
rect 30745 15079 30803 15085
rect 26016 15036 26022 15048
rect 26234 15008 26240 15020
rect 24268 14980 25912 15008
rect 26195 14980 26240 15008
rect 24268 14968 24274 14980
rect 26234 14968 26240 14980
rect 26292 14968 26298 15020
rect 26421 15011 26479 15017
rect 26421 14977 26433 15011
rect 26467 15008 26479 15011
rect 26970 15008 26976 15020
rect 26467 14980 26976 15008
rect 26467 14977 26479 14980
rect 26421 14971 26479 14977
rect 26970 14968 26976 14980
rect 27028 14968 27034 15020
rect 27172 15017 27200 15048
rect 30745 15045 30757 15079
rect 30791 15076 30803 15079
rect 30834 15076 30840 15088
rect 30791 15048 30840 15076
rect 30791 15045 30803 15048
rect 30745 15039 30803 15045
rect 30834 15036 30840 15048
rect 30892 15036 30898 15088
rect 33226 15076 33232 15088
rect 32232 15048 33232 15076
rect 27157 15011 27215 15017
rect 27157 14977 27169 15011
rect 27203 14977 27215 15011
rect 27157 14971 27215 14977
rect 27430 14968 27436 15020
rect 27488 15008 27494 15020
rect 32232 15017 32260 15048
rect 33226 15036 33232 15048
rect 33284 15036 33290 15088
rect 28077 15011 28135 15017
rect 28077 15008 28089 15011
rect 27488 14980 28089 15008
rect 27488 14968 27494 14980
rect 28077 14977 28089 14980
rect 28123 14977 28135 15011
rect 28988 15011 29046 15017
rect 28988 15008 29000 15011
rect 28077 14971 28135 14977
rect 28368 14980 29000 15008
rect 18693 14943 18751 14949
rect 18693 14909 18705 14943
rect 18739 14909 18751 14943
rect 18693 14903 18751 14909
rect 18708 14872 18736 14903
rect 18782 14900 18788 14952
rect 18840 14940 18846 14952
rect 19245 14943 19303 14949
rect 19245 14940 19257 14943
rect 18840 14912 19257 14940
rect 18840 14900 18846 14912
rect 19245 14909 19257 14912
rect 19291 14940 19303 14943
rect 22097 14943 22155 14949
rect 22097 14940 22109 14943
rect 19291 14912 22109 14940
rect 19291 14909 19303 14912
rect 19245 14903 19303 14909
rect 22097 14909 22109 14912
rect 22143 14940 22155 14943
rect 23290 14940 23296 14952
rect 22143 14912 23296 14940
rect 22143 14909 22155 14912
rect 22097 14903 22155 14909
rect 23290 14900 23296 14912
rect 23348 14900 23354 14952
rect 27062 14940 27068 14952
rect 27023 14912 27068 14940
rect 27062 14900 27068 14912
rect 27120 14900 27126 14952
rect 18708 14844 22094 14872
rect 13449 14807 13507 14813
rect 13449 14773 13461 14807
rect 13495 14804 13507 14807
rect 14274 14804 14280 14816
rect 13495 14776 14280 14804
rect 13495 14773 13507 14776
rect 13449 14767 13507 14773
rect 14274 14764 14280 14776
rect 14332 14764 14338 14816
rect 17681 14807 17739 14813
rect 17681 14773 17693 14807
rect 17727 14804 17739 14807
rect 18046 14804 18052 14816
rect 17727 14776 18052 14804
rect 17727 14773 17739 14776
rect 17681 14767 17739 14773
rect 18046 14764 18052 14776
rect 18104 14764 18110 14816
rect 18325 14807 18383 14813
rect 18325 14773 18337 14807
rect 18371 14804 18383 14807
rect 19242 14804 19248 14816
rect 18371 14776 19248 14804
rect 18371 14773 18383 14776
rect 18325 14767 18383 14773
rect 19242 14764 19248 14776
rect 19300 14764 19306 14816
rect 19337 14807 19395 14813
rect 19337 14773 19349 14807
rect 19383 14804 19395 14807
rect 19426 14804 19432 14816
rect 19383 14776 19432 14804
rect 19383 14773 19395 14776
rect 19337 14767 19395 14773
rect 19426 14764 19432 14776
rect 19484 14764 19490 14816
rect 19702 14804 19708 14816
rect 19663 14776 19708 14804
rect 19702 14764 19708 14776
rect 19760 14764 19766 14816
rect 20901 14807 20959 14813
rect 20901 14773 20913 14807
rect 20947 14804 20959 14807
rect 21082 14804 21088 14816
rect 20947 14776 21088 14804
rect 20947 14773 20959 14776
rect 20901 14767 20959 14773
rect 21082 14764 21088 14776
rect 21140 14764 21146 14816
rect 22066 14804 22094 14844
rect 22830 14832 22836 14884
rect 22888 14872 22894 14884
rect 23842 14872 23848 14884
rect 22888 14844 23848 14872
rect 22888 14832 22894 14844
rect 23842 14832 23848 14844
rect 23900 14872 23906 14884
rect 24121 14875 24179 14881
rect 24121 14872 24133 14875
rect 23900 14844 24133 14872
rect 23900 14832 23906 14844
rect 24121 14841 24133 14844
rect 24167 14841 24179 14875
rect 26418 14872 26424 14884
rect 24121 14835 24179 14841
rect 25424 14844 26424 14872
rect 25424 14804 25452 14844
rect 26418 14832 26424 14844
rect 26476 14832 26482 14884
rect 28261 14875 28319 14881
rect 28261 14841 28273 14875
rect 28307 14872 28319 14875
rect 28368 14872 28396 14980
rect 28988 14977 29000 14980
rect 29034 15008 29046 15011
rect 32217 15011 32275 15017
rect 29034 14980 31754 15008
rect 29034 14977 29046 14980
rect 28988 14971 29046 14977
rect 28442 14900 28448 14952
rect 28500 14940 28506 14952
rect 28721 14943 28779 14949
rect 28721 14940 28733 14943
rect 28500 14912 28733 14940
rect 28500 14900 28506 14912
rect 28721 14909 28733 14912
rect 28767 14909 28779 14943
rect 28721 14903 28779 14909
rect 28307 14844 28396 14872
rect 28307 14841 28319 14844
rect 28261 14835 28319 14841
rect 30190 14832 30196 14884
rect 30248 14872 30254 14884
rect 31113 14875 31171 14881
rect 31113 14872 31125 14875
rect 30248 14844 31125 14872
rect 30248 14832 30254 14844
rect 31113 14841 31125 14844
rect 31159 14841 31171 14875
rect 31726 14872 31754 14980
rect 32217 14977 32229 15011
rect 32263 14977 32275 15011
rect 32217 14971 32275 14977
rect 32401 15011 32459 15017
rect 32401 14977 32413 15011
rect 32447 14977 32459 15011
rect 32401 14971 32459 14977
rect 32677 15011 32735 15017
rect 32677 14977 32689 15011
rect 32723 15008 32735 15011
rect 33134 15008 33140 15020
rect 32723 14980 33140 15008
rect 32723 14977 32735 14980
rect 32677 14971 32735 14977
rect 32416 14940 32444 14971
rect 33134 14968 33140 14980
rect 33192 14968 33198 15020
rect 33594 15008 33600 15020
rect 33555 14980 33600 15008
rect 33594 14968 33600 14980
rect 33652 14968 33658 15020
rect 33873 15011 33931 15017
rect 33873 14977 33885 15011
rect 33919 15008 33931 15011
rect 34054 15008 34060 15020
rect 33919 14980 34060 15008
rect 33919 14977 33931 14980
rect 33873 14971 33931 14977
rect 33888 14940 33916 14971
rect 34054 14968 34060 14980
rect 34112 14968 34118 15020
rect 32416 14912 33916 14940
rect 32214 14872 32220 14884
rect 31726 14844 32220 14872
rect 31113 14835 31171 14841
rect 32214 14832 32220 14844
rect 32272 14872 32278 14884
rect 32950 14872 32956 14884
rect 32272 14844 32956 14872
rect 32272 14832 32278 14844
rect 32950 14832 32956 14844
rect 33008 14832 33014 14884
rect 34164 14872 34192 15116
rect 35345 15113 35357 15147
rect 35391 15144 35403 15147
rect 39485 15147 39543 15153
rect 39485 15144 39497 15147
rect 35391 15116 39497 15144
rect 35391 15113 35403 15116
rect 35345 15107 35403 15113
rect 39485 15113 39497 15116
rect 39531 15113 39543 15147
rect 39485 15107 39543 15113
rect 43441 15147 43499 15153
rect 43441 15113 43453 15147
rect 43487 15144 43499 15147
rect 43990 15144 43996 15156
rect 43487 15116 43996 15144
rect 43487 15113 43499 15116
rect 43441 15107 43499 15113
rect 43990 15104 43996 15116
rect 44048 15104 44054 15156
rect 36078 15036 36084 15088
rect 36136 15076 36142 15088
rect 36567 15079 36625 15085
rect 36567 15076 36579 15079
rect 36136 15048 36579 15076
rect 36136 15036 36142 15048
rect 36567 15045 36579 15048
rect 36613 15045 36625 15079
rect 36567 15039 36625 15045
rect 37274 15036 37280 15088
rect 37332 15076 37338 15088
rect 39117 15079 39175 15085
rect 39117 15076 39129 15079
rect 37332 15048 39129 15076
rect 37332 15036 37338 15048
rect 39117 15045 39129 15048
rect 39163 15045 39175 15079
rect 39117 15039 39175 15045
rect 35253 15011 35311 15017
rect 35253 14977 35265 15011
rect 35299 15008 35311 15011
rect 35986 15008 35992 15020
rect 35299 14980 35992 15008
rect 35299 14977 35311 14980
rect 35253 14971 35311 14977
rect 35986 14968 35992 14980
rect 36044 14968 36050 15020
rect 36262 15008 36268 15020
rect 36223 14980 36268 15008
rect 36262 14968 36268 14980
rect 36320 14968 36326 15020
rect 36357 15011 36415 15017
rect 36357 14977 36369 15011
rect 36403 14977 36415 15011
rect 36357 14971 36415 14977
rect 34241 14943 34299 14949
rect 34241 14909 34253 14943
rect 34287 14940 34299 14943
rect 35526 14940 35532 14952
rect 34287 14912 35532 14940
rect 34287 14909 34299 14912
rect 34241 14903 34299 14909
rect 35526 14900 35532 14912
rect 35584 14900 35590 14952
rect 36372 14940 36400 14971
rect 36446 14968 36452 15020
rect 36504 15008 36510 15020
rect 36725 15011 36783 15017
rect 36504 14980 36549 15008
rect 36504 14968 36510 14980
rect 36725 14977 36737 15011
rect 36771 15008 36783 15011
rect 36814 15008 36820 15020
rect 36771 14980 36820 15008
rect 36771 14977 36783 14980
rect 36725 14971 36783 14977
rect 36814 14968 36820 14980
rect 36872 14968 36878 15020
rect 37458 14968 37464 15020
rect 37516 15008 37522 15020
rect 38841 15011 38899 15017
rect 38841 15008 38853 15011
rect 37516 14980 38853 15008
rect 37516 14968 37522 14980
rect 38841 14977 38853 14980
rect 38887 14977 38899 15011
rect 38841 14971 38899 14977
rect 38930 14968 38936 15020
rect 38988 15008 38994 15020
rect 39209 15011 39267 15017
rect 38988 14980 39033 15008
rect 38988 14968 38994 14980
rect 39209 14977 39221 15011
rect 39255 14977 39267 15011
rect 39209 14971 39267 14977
rect 39306 15011 39364 15017
rect 39306 14977 39318 15011
rect 39352 14977 39364 15011
rect 39306 14971 39364 14977
rect 43349 15011 43407 15017
rect 43349 14977 43361 15011
rect 43395 15008 43407 15011
rect 43898 15008 43904 15020
rect 43395 14980 43904 15008
rect 43395 14977 43407 14980
rect 43349 14971 43407 14977
rect 36372 14912 37320 14940
rect 36538 14872 36544 14884
rect 34164 14844 36544 14872
rect 36538 14832 36544 14844
rect 36596 14832 36602 14884
rect 37292 14872 37320 14912
rect 37366 14900 37372 14952
rect 37424 14940 37430 14952
rect 37553 14943 37611 14949
rect 37553 14940 37565 14943
rect 37424 14912 37565 14940
rect 37424 14900 37430 14912
rect 37553 14909 37565 14912
rect 37599 14909 37611 14943
rect 37553 14903 37611 14909
rect 37829 14943 37887 14949
rect 37829 14909 37841 14943
rect 37875 14909 37887 14943
rect 37829 14903 37887 14909
rect 37458 14872 37464 14884
rect 37292 14844 37464 14872
rect 37458 14832 37464 14844
rect 37516 14832 37522 14884
rect 37642 14832 37648 14884
rect 37700 14872 37706 14884
rect 37844 14872 37872 14903
rect 37918 14900 37924 14952
rect 37976 14940 37982 14952
rect 38378 14940 38384 14952
rect 37976 14912 38384 14940
rect 37976 14900 37982 14912
rect 38378 14900 38384 14912
rect 38436 14940 38442 14952
rect 39224 14940 39252 14971
rect 38436 14912 39252 14940
rect 38436 14900 38442 14912
rect 39316 14872 39344 14971
rect 43898 14968 43904 14980
rect 43956 14968 43962 15020
rect 37700 14844 39344 14872
rect 37700 14832 37706 14844
rect 22066 14776 25452 14804
rect 26329 14807 26387 14813
rect 26329 14773 26341 14807
rect 26375 14804 26387 14807
rect 26970 14804 26976 14816
rect 26375 14776 26976 14804
rect 26375 14773 26387 14776
rect 26329 14767 26387 14773
rect 26970 14764 26976 14776
rect 27028 14764 27034 14816
rect 27525 14807 27583 14813
rect 27525 14773 27537 14807
rect 27571 14804 27583 14807
rect 28350 14804 28356 14816
rect 27571 14776 28356 14804
rect 27571 14773 27583 14776
rect 27525 14767 27583 14773
rect 28350 14764 28356 14776
rect 28408 14764 28414 14816
rect 30006 14764 30012 14816
rect 30064 14804 30070 14816
rect 30101 14807 30159 14813
rect 30101 14804 30113 14807
rect 30064 14776 30113 14804
rect 30064 14764 30070 14776
rect 30101 14773 30113 14776
rect 30147 14773 30159 14807
rect 30101 14767 30159 14773
rect 30650 14764 30656 14816
rect 30708 14804 30714 14816
rect 30745 14807 30803 14813
rect 30745 14804 30757 14807
rect 30708 14776 30757 14804
rect 30708 14764 30714 14776
rect 30745 14773 30757 14776
rect 30791 14773 30803 14807
rect 32398 14804 32404 14816
rect 32359 14776 32404 14804
rect 30745 14767 30803 14773
rect 32398 14764 32404 14776
rect 32456 14764 32462 14816
rect 34422 14764 34428 14816
rect 34480 14804 34486 14816
rect 34885 14807 34943 14813
rect 34885 14804 34897 14807
rect 34480 14776 34897 14804
rect 34480 14764 34486 14776
rect 34885 14773 34897 14776
rect 34931 14773 34943 14807
rect 34885 14767 34943 14773
rect 35342 14764 35348 14816
rect 35400 14804 35406 14816
rect 36081 14807 36139 14813
rect 36081 14804 36093 14807
rect 35400 14776 36093 14804
rect 35400 14764 35406 14776
rect 36081 14773 36093 14776
rect 36127 14773 36139 14807
rect 36081 14767 36139 14773
rect 37274 14764 37280 14816
rect 37332 14804 37338 14816
rect 38286 14804 38292 14816
rect 37332 14776 38292 14804
rect 37332 14764 37338 14776
rect 38286 14764 38292 14776
rect 38344 14804 38350 14816
rect 38930 14804 38936 14816
rect 38344 14776 38936 14804
rect 38344 14764 38350 14776
rect 38930 14764 38936 14776
rect 38988 14764 38994 14816
rect 1104 14714 44896 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 44896 14714
rect 1104 14640 44896 14662
rect 18233 14603 18291 14609
rect 18233 14569 18245 14603
rect 18279 14600 18291 14603
rect 18506 14600 18512 14612
rect 18279 14572 18512 14600
rect 18279 14569 18291 14572
rect 18233 14563 18291 14569
rect 18506 14560 18512 14572
rect 18564 14560 18570 14612
rect 21821 14603 21879 14609
rect 21821 14569 21833 14603
rect 21867 14600 21879 14603
rect 22002 14600 22008 14612
rect 21867 14572 22008 14600
rect 21867 14569 21879 14572
rect 21821 14563 21879 14569
rect 22002 14560 22008 14572
rect 22060 14560 22066 14612
rect 22833 14603 22891 14609
rect 22833 14569 22845 14603
rect 22879 14600 22891 14603
rect 22922 14600 22928 14612
rect 22879 14572 22928 14600
rect 22879 14569 22891 14572
rect 22833 14563 22891 14569
rect 22922 14560 22928 14572
rect 22980 14560 22986 14612
rect 25961 14603 26019 14609
rect 25961 14569 25973 14603
rect 26007 14600 26019 14603
rect 26234 14600 26240 14612
rect 26007 14572 26240 14600
rect 26007 14569 26019 14572
rect 25961 14563 26019 14569
rect 26234 14560 26240 14572
rect 26292 14560 26298 14612
rect 27062 14600 27068 14612
rect 27023 14572 27068 14600
rect 27062 14560 27068 14572
rect 27120 14560 27126 14612
rect 27430 14600 27436 14612
rect 27391 14572 27436 14600
rect 27430 14560 27436 14572
rect 27488 14560 27494 14612
rect 30006 14600 30012 14612
rect 29967 14572 30012 14600
rect 30006 14560 30012 14572
rect 30064 14560 30070 14612
rect 30190 14600 30196 14612
rect 30151 14572 30196 14600
rect 30190 14560 30196 14572
rect 30248 14560 30254 14612
rect 35986 14560 35992 14612
rect 36044 14600 36050 14612
rect 36173 14603 36231 14609
rect 36173 14600 36185 14603
rect 36044 14572 36185 14600
rect 36044 14560 36050 14572
rect 36173 14569 36185 14572
rect 36219 14569 36231 14603
rect 36173 14563 36231 14569
rect 36538 14560 36544 14612
rect 36596 14600 36602 14612
rect 43898 14600 43904 14612
rect 36596 14572 43904 14600
rect 36596 14560 36602 14572
rect 43898 14560 43904 14572
rect 43956 14560 43962 14612
rect 20993 14535 21051 14541
rect 20993 14501 21005 14535
rect 21039 14532 21051 14535
rect 22186 14532 22192 14544
rect 21039 14504 22192 14532
rect 21039 14501 21051 14504
rect 20993 14495 21051 14501
rect 22186 14492 22192 14504
rect 22244 14492 22250 14544
rect 26142 14532 26148 14544
rect 26103 14504 26148 14532
rect 26142 14492 26148 14504
rect 26200 14492 26206 14544
rect 36446 14532 36452 14544
rect 33980 14504 36452 14532
rect 14274 14464 14280 14476
rect 14235 14436 14280 14464
rect 14274 14424 14280 14436
rect 14332 14424 14338 14476
rect 18782 14464 18788 14476
rect 18156 14436 18788 14464
rect 2038 14356 2044 14408
rect 2096 14396 2102 14408
rect 2133 14399 2191 14405
rect 2133 14396 2145 14399
rect 2096 14368 2145 14396
rect 2096 14356 2102 14368
rect 2133 14365 2145 14368
rect 2179 14365 2191 14399
rect 2133 14359 2191 14365
rect 3053 14399 3111 14405
rect 3053 14365 3065 14399
rect 3099 14396 3111 14399
rect 9214 14396 9220 14408
rect 3099 14368 9220 14396
rect 3099 14365 3111 14368
rect 3053 14359 3111 14365
rect 9214 14356 9220 14368
rect 9272 14356 9278 14408
rect 13998 14356 14004 14408
rect 14056 14396 14062 14408
rect 14093 14399 14151 14405
rect 14093 14396 14105 14399
rect 14056 14368 14105 14396
rect 14056 14356 14062 14368
rect 14093 14365 14105 14368
rect 14139 14365 14151 14399
rect 14093 14359 14151 14365
rect 17865 14399 17923 14405
rect 17865 14365 17877 14399
rect 17911 14365 17923 14399
rect 17865 14359 17923 14365
rect 15930 14328 15936 14340
rect 15891 14300 15936 14328
rect 15930 14288 15936 14300
rect 15988 14288 15994 14340
rect 17880 14328 17908 14359
rect 18046 14356 18052 14408
rect 18104 14396 18110 14408
rect 18156 14396 18184 14436
rect 18782 14424 18788 14436
rect 18840 14424 18846 14476
rect 22002 14424 22008 14476
rect 22060 14464 22066 14476
rect 25774 14464 25780 14476
rect 22060 14424 22094 14464
rect 25735 14436 25780 14464
rect 25774 14424 25780 14436
rect 25832 14424 25838 14476
rect 29914 14464 29920 14476
rect 29875 14436 29920 14464
rect 29914 14424 29920 14436
rect 29972 14424 29978 14476
rect 30190 14424 30196 14476
rect 30248 14464 30254 14476
rect 31205 14467 31263 14473
rect 31205 14464 31217 14467
rect 30248 14436 31217 14464
rect 30248 14424 30254 14436
rect 31205 14433 31217 14436
rect 31251 14433 31263 14467
rect 31205 14427 31263 14433
rect 31665 14467 31723 14473
rect 31665 14433 31677 14467
rect 31711 14464 31723 14467
rect 32585 14467 32643 14473
rect 32585 14464 32597 14467
rect 31711 14436 32597 14464
rect 31711 14433 31723 14436
rect 31665 14427 31723 14433
rect 32585 14433 32597 14436
rect 32631 14433 32643 14467
rect 32585 14427 32643 14433
rect 18322 14396 18328 14408
rect 18104 14368 18197 14396
rect 18283 14368 18328 14396
rect 18104 14356 18110 14368
rect 18322 14356 18328 14368
rect 18380 14356 18386 14408
rect 19334 14356 19340 14408
rect 19392 14396 19398 14408
rect 19613 14399 19671 14405
rect 19613 14396 19625 14399
rect 19392 14368 19625 14396
rect 19392 14356 19398 14368
rect 19613 14365 19625 14368
rect 19659 14365 19671 14399
rect 19613 14359 19671 14365
rect 19702 14356 19708 14408
rect 19760 14396 19766 14408
rect 19869 14399 19927 14405
rect 19869 14396 19881 14399
rect 19760 14368 19881 14396
rect 19760 14356 19766 14368
rect 19869 14365 19881 14368
rect 19915 14365 19927 14399
rect 22066 14396 22094 14424
rect 22557 14399 22615 14405
rect 22557 14396 22569 14399
rect 22066 14368 22569 14396
rect 19869 14359 19927 14365
rect 22557 14365 22569 14368
rect 22603 14365 22615 14399
rect 22557 14359 22615 14365
rect 18138 14328 18144 14340
rect 17880 14300 18144 14328
rect 18138 14288 18144 14300
rect 18196 14288 18202 14340
rect 21805 14331 21863 14337
rect 21805 14297 21817 14331
rect 21851 14328 21863 14331
rect 21910 14328 21916 14340
rect 21851 14300 21916 14328
rect 21851 14297 21863 14300
rect 21805 14291 21863 14297
rect 21910 14288 21916 14300
rect 21968 14288 21974 14340
rect 22005 14331 22063 14337
rect 22005 14297 22017 14331
rect 22051 14328 22063 14331
rect 22094 14328 22100 14340
rect 22051 14300 22100 14328
rect 22051 14297 22063 14300
rect 22005 14291 22063 14297
rect 22094 14288 22100 14300
rect 22152 14328 22158 14340
rect 22278 14328 22284 14340
rect 22152 14300 22284 14328
rect 22152 14288 22158 14300
rect 22278 14288 22284 14300
rect 22336 14288 22342 14340
rect 22572 14328 22600 14359
rect 22646 14356 22652 14408
rect 22704 14396 22710 14408
rect 23661 14399 23719 14405
rect 23661 14396 23673 14399
rect 22704 14368 23673 14396
rect 22704 14356 22710 14368
rect 23661 14365 23673 14368
rect 23707 14365 23719 14399
rect 25958 14396 25964 14408
rect 25919 14368 25964 14396
rect 23661 14359 23719 14365
rect 25958 14356 25964 14368
rect 26016 14356 26022 14408
rect 26970 14396 26976 14408
rect 26931 14368 26976 14396
rect 26970 14356 26976 14368
rect 27028 14356 27034 14408
rect 30009 14399 30067 14405
rect 30009 14365 30021 14399
rect 30055 14396 30067 14399
rect 30098 14396 30104 14408
rect 30055 14368 30104 14396
rect 30055 14365 30067 14368
rect 30009 14359 30067 14365
rect 30098 14356 30104 14368
rect 30156 14356 30162 14408
rect 31297 14399 31355 14405
rect 31297 14365 31309 14399
rect 31343 14396 31355 14399
rect 31570 14396 31576 14408
rect 31343 14368 31576 14396
rect 31343 14365 31355 14368
rect 31297 14359 31355 14365
rect 31570 14356 31576 14368
rect 31628 14356 31634 14408
rect 32398 14356 32404 14408
rect 32456 14396 32462 14408
rect 33980 14405 34008 14504
rect 36446 14492 36452 14504
rect 36504 14492 36510 14544
rect 38013 14535 38071 14541
rect 38013 14532 38025 14535
rect 36648 14504 38025 14532
rect 34164 14436 35480 14464
rect 34164 14405 34192 14436
rect 32677 14399 32735 14405
rect 32677 14396 32689 14399
rect 32456 14368 32689 14396
rect 32456 14356 32462 14368
rect 32677 14365 32689 14368
rect 32723 14365 32735 14399
rect 32677 14359 32735 14365
rect 33965 14399 34023 14405
rect 33965 14365 33977 14399
rect 34011 14365 34023 14399
rect 33965 14359 34023 14365
rect 34149 14399 34207 14405
rect 34149 14365 34161 14399
rect 34195 14365 34207 14399
rect 35342 14396 35348 14408
rect 35303 14368 35348 14396
rect 34149 14359 34207 14365
rect 35342 14356 35348 14368
rect 35400 14356 35406 14408
rect 35452 14396 35480 14436
rect 35526 14424 35532 14476
rect 35584 14464 35590 14476
rect 35584 14436 35629 14464
rect 35584 14424 35590 14436
rect 36648 14405 36676 14504
rect 38013 14501 38025 14504
rect 38059 14501 38071 14535
rect 38013 14495 38071 14501
rect 38194 14492 38200 14544
rect 38252 14532 38258 14544
rect 38565 14535 38623 14541
rect 38565 14532 38577 14535
rect 38252 14504 38577 14532
rect 38252 14492 38258 14504
rect 38565 14501 38577 14504
rect 38611 14501 38623 14535
rect 38565 14495 38623 14501
rect 36725 14467 36783 14473
rect 36725 14433 36737 14467
rect 36771 14433 36783 14467
rect 36725 14427 36783 14433
rect 36633 14399 36691 14405
rect 36633 14396 36645 14399
rect 35452 14368 36645 14396
rect 36633 14365 36645 14368
rect 36679 14365 36691 14399
rect 36740 14396 36768 14427
rect 36814 14424 36820 14476
rect 36872 14464 36878 14476
rect 37369 14467 37427 14473
rect 37369 14464 37381 14467
rect 36872 14436 37381 14464
rect 36872 14424 36878 14436
rect 37369 14433 37381 14436
rect 37415 14464 37427 14467
rect 37458 14464 37464 14476
rect 37415 14436 37464 14464
rect 37415 14433 37427 14436
rect 37369 14427 37427 14433
rect 37458 14424 37464 14436
rect 37516 14424 37522 14476
rect 37734 14464 37740 14476
rect 37695 14436 37740 14464
rect 37734 14424 37740 14436
rect 37792 14424 37798 14476
rect 37829 14467 37887 14473
rect 37829 14433 37841 14467
rect 37875 14464 37887 14467
rect 39022 14464 39028 14476
rect 37875 14436 39028 14464
rect 37875 14433 37887 14436
rect 37829 14427 37887 14433
rect 39022 14424 39028 14436
rect 39080 14424 39086 14476
rect 42337 14467 42395 14473
rect 42337 14433 42349 14467
rect 42383 14464 42395 14467
rect 42702 14464 42708 14476
rect 42383 14436 42708 14464
rect 42383 14433 42395 14436
rect 42337 14427 42395 14433
rect 42702 14424 42708 14436
rect 42760 14424 42766 14476
rect 44082 14464 44088 14476
rect 44043 14436 44088 14464
rect 44082 14424 44088 14436
rect 44140 14424 44146 14476
rect 37274 14396 37280 14408
rect 36740 14368 37280 14396
rect 36633 14359 36691 14365
rect 37274 14356 37280 14368
rect 37332 14356 37338 14408
rect 38010 14356 38016 14408
rect 38068 14396 38074 14408
rect 38465 14399 38523 14405
rect 38465 14396 38477 14399
rect 38068 14368 38477 14396
rect 38068 14356 38074 14368
rect 38465 14365 38477 14368
rect 38511 14365 38523 14399
rect 38465 14359 38523 14365
rect 38562 14356 38568 14408
rect 38620 14396 38626 14408
rect 38657 14399 38715 14405
rect 38657 14396 38669 14399
rect 38620 14368 38669 14396
rect 38620 14356 38626 14368
rect 38657 14365 38669 14368
rect 38703 14365 38715 14399
rect 38657 14359 38715 14365
rect 23477 14331 23535 14337
rect 23477 14328 23489 14331
rect 22572 14300 23489 14328
rect 23477 14297 23489 14300
rect 23523 14297 23535 14331
rect 25682 14328 25688 14340
rect 25643 14300 25688 14328
rect 23477 14291 23535 14297
rect 25682 14288 25688 14300
rect 25740 14288 25746 14340
rect 29638 14288 29644 14340
rect 29696 14328 29702 14340
rect 29733 14331 29791 14337
rect 29733 14328 29745 14331
rect 29696 14300 29745 14328
rect 29696 14288 29702 14300
rect 29733 14297 29745 14300
rect 29779 14297 29791 14331
rect 29733 14291 29791 14297
rect 34057 14331 34115 14337
rect 34057 14297 34069 14331
rect 34103 14328 34115 14331
rect 35437 14331 35495 14337
rect 35437 14328 35449 14331
rect 34103 14300 35449 14328
rect 34103 14297 34115 14300
rect 34057 14291 34115 14297
rect 35437 14297 35449 14300
rect 35483 14297 35495 14331
rect 38930 14328 38936 14340
rect 35437 14291 35495 14297
rect 38626 14300 38936 14328
rect 38626 14272 38654 14300
rect 38930 14288 38936 14300
rect 38988 14288 38994 14340
rect 42521 14331 42579 14337
rect 42521 14297 42533 14331
rect 42567 14328 42579 14331
rect 43438 14328 43444 14340
rect 42567 14300 43444 14328
rect 42567 14297 42579 14300
rect 42521 14291 42579 14297
rect 43438 14288 43444 14300
rect 43496 14288 43502 14340
rect 2222 14220 2228 14272
rect 2280 14260 2286 14272
rect 2961 14263 3019 14269
rect 2961 14260 2973 14263
rect 2280 14232 2973 14260
rect 2280 14220 2286 14232
rect 2961 14229 2973 14232
rect 3007 14229 3019 14263
rect 2961 14223 3019 14229
rect 20714 14220 20720 14272
rect 20772 14260 20778 14272
rect 21634 14260 21640 14272
rect 20772 14232 21640 14260
rect 20772 14220 20778 14232
rect 21634 14220 21640 14232
rect 21692 14220 21698 14272
rect 23290 14260 23296 14272
rect 23251 14232 23296 14260
rect 23290 14220 23296 14232
rect 23348 14220 23354 14272
rect 33502 14260 33508 14272
rect 33463 14232 33508 14260
rect 33502 14220 33508 14232
rect 33560 14220 33566 14272
rect 34330 14220 34336 14272
rect 34388 14260 34394 14272
rect 34977 14263 35035 14269
rect 34977 14260 34989 14263
rect 34388 14232 34989 14260
rect 34388 14220 34394 14232
rect 34977 14229 34989 14232
rect 35023 14229 35035 14263
rect 36538 14260 36544 14272
rect 36499 14232 36544 14260
rect 34977 14223 35035 14229
rect 36538 14220 36544 14232
rect 36596 14220 36602 14272
rect 38562 14220 38568 14272
rect 38620 14232 38654 14272
rect 38620 14220 38626 14232
rect 1104 14170 44896 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 44896 14170
rect 1104 14096 44896 14118
rect 13998 14056 14004 14068
rect 13959 14028 14004 14056
rect 13998 14016 14004 14028
rect 14056 14016 14062 14068
rect 17954 14016 17960 14068
rect 18012 14056 18018 14068
rect 20349 14059 20407 14065
rect 20349 14056 20361 14059
rect 18012 14028 20361 14056
rect 18012 14016 18018 14028
rect 20349 14025 20361 14028
rect 20395 14025 20407 14059
rect 21174 14056 21180 14068
rect 21135 14028 21180 14056
rect 20349 14019 20407 14025
rect 21174 14016 21180 14028
rect 21232 14016 21238 14068
rect 22646 14016 22652 14068
rect 22704 14056 22710 14068
rect 23569 14059 23627 14065
rect 23569 14056 23581 14059
rect 22704 14028 23581 14056
rect 22704 14016 22710 14028
rect 23569 14025 23581 14028
rect 23615 14025 23627 14059
rect 23569 14019 23627 14025
rect 25866 14016 25872 14068
rect 25924 14056 25930 14068
rect 26145 14059 26203 14065
rect 26145 14056 26157 14059
rect 25924 14028 26157 14056
rect 25924 14016 25930 14028
rect 26145 14025 26157 14028
rect 26191 14025 26203 14059
rect 29638 14056 29644 14068
rect 29599 14028 29644 14056
rect 26145 14019 26203 14025
rect 29638 14016 29644 14028
rect 29696 14016 29702 14068
rect 30098 14056 30104 14068
rect 30059 14028 30104 14056
rect 30098 14016 30104 14028
rect 30156 14016 30162 14068
rect 32309 14059 32367 14065
rect 32309 14025 32321 14059
rect 32355 14056 32367 14059
rect 33226 14056 33232 14068
rect 32355 14028 33232 14056
rect 32355 14025 32367 14028
rect 32309 14019 32367 14025
rect 33226 14016 33232 14028
rect 33284 14016 33290 14068
rect 34330 14056 34336 14068
rect 34291 14028 34336 14056
rect 34330 14016 34336 14028
rect 34388 14016 34394 14068
rect 34422 14016 34428 14068
rect 34480 14056 34486 14068
rect 34480 14028 34525 14056
rect 34480 14016 34486 14028
rect 36538 14016 36544 14068
rect 36596 14056 36602 14068
rect 37445 14059 37503 14065
rect 37445 14056 37457 14059
rect 36596 14028 37457 14056
rect 36596 14016 36602 14028
rect 37445 14025 37457 14028
rect 37491 14056 37503 14059
rect 38194 14056 38200 14068
rect 37491 14028 38200 14056
rect 37491 14025 37503 14028
rect 37445 14019 37503 14025
rect 38194 14016 38200 14028
rect 38252 14016 38258 14068
rect 38378 14016 38384 14068
rect 38436 14056 38442 14068
rect 38562 14056 38568 14068
rect 38436 14028 38568 14056
rect 38436 14016 38442 14028
rect 38562 14016 38568 14028
rect 38620 14056 38626 14068
rect 38620 14028 39620 14056
rect 38620 14016 38626 14028
rect 2222 13988 2228 14000
rect 2183 13960 2228 13988
rect 2222 13948 2228 13960
rect 2280 13948 2286 14000
rect 18046 13988 18052 14000
rect 13832 13960 18052 13988
rect 2038 13920 2044 13932
rect 1999 13892 2044 13920
rect 2038 13880 2044 13892
rect 2096 13880 2102 13932
rect 13832 13929 13860 13960
rect 18046 13948 18052 13960
rect 18104 13948 18110 14000
rect 19058 13948 19064 14000
rect 19116 13988 19122 14000
rect 20165 13991 20223 13997
rect 19116 13960 20024 13988
rect 19116 13948 19122 13960
rect 13817 13923 13875 13929
rect 13817 13889 13829 13923
rect 13863 13889 13875 13923
rect 16666 13920 16672 13932
rect 16627 13892 16672 13920
rect 13817 13883 13875 13889
rect 16666 13880 16672 13892
rect 16724 13880 16730 13932
rect 16942 13929 16948 13932
rect 16936 13883 16948 13929
rect 17000 13920 17006 13932
rect 17000 13892 17036 13920
rect 18984 13892 19380 13920
rect 16942 13880 16948 13883
rect 17000 13880 17006 13892
rect 2774 13852 2780 13864
rect 2735 13824 2780 13852
rect 2774 13812 2780 13824
rect 2832 13812 2838 13864
rect 18322 13852 18328 13864
rect 18064 13824 18328 13852
rect 18064 13793 18092 13824
rect 18322 13812 18328 13824
rect 18380 13852 18386 13864
rect 18984 13852 19012 13892
rect 18380 13824 19012 13852
rect 18380 13812 18386 13824
rect 19058 13812 19064 13864
rect 19116 13852 19122 13864
rect 19352 13861 19380 13892
rect 19426 13880 19432 13932
rect 19484 13920 19490 13932
rect 19797 13923 19855 13929
rect 19797 13920 19809 13923
rect 19484 13892 19809 13920
rect 19484 13880 19490 13892
rect 19797 13889 19809 13892
rect 19843 13889 19855 13923
rect 19996 13920 20024 13960
rect 20165 13957 20177 13991
rect 20211 13988 20223 13991
rect 20809 13991 20867 13997
rect 20809 13988 20821 13991
rect 20211 13960 20821 13988
rect 20211 13957 20223 13960
rect 20165 13951 20223 13957
rect 20809 13957 20821 13960
rect 20855 13957 20867 13991
rect 21818 13988 21824 14000
rect 20809 13951 20867 13957
rect 21008 13960 21824 13988
rect 21008 13929 21036 13960
rect 21818 13948 21824 13960
rect 21876 13948 21882 14000
rect 22830 13988 22836 14000
rect 22204 13960 22836 13988
rect 20993 13923 21051 13929
rect 20993 13920 21005 13923
rect 19996 13892 21005 13920
rect 19797 13883 19855 13889
rect 20993 13889 21005 13892
rect 21039 13889 21051 13923
rect 21266 13920 21272 13932
rect 21227 13892 21272 13920
rect 20993 13883 21051 13889
rect 21266 13880 21272 13892
rect 21324 13880 21330 13932
rect 22204 13929 22232 13960
rect 22830 13948 22836 13960
rect 22888 13948 22894 14000
rect 27709 13991 27767 13997
rect 27709 13957 27721 13991
rect 27755 13988 27767 13991
rect 29730 13988 29736 14000
rect 27755 13960 29736 13988
rect 27755 13957 27767 13960
rect 27709 13951 27767 13957
rect 29730 13948 29736 13960
rect 29788 13948 29794 14000
rect 37090 13948 37096 14000
rect 37148 13988 37154 14000
rect 37645 13991 37703 13997
rect 37645 13988 37657 13991
rect 37148 13960 37657 13988
rect 37148 13948 37154 13960
rect 37645 13957 37657 13960
rect 37691 13957 37703 13991
rect 37645 13951 37703 13957
rect 37734 13948 37740 14000
rect 37792 13988 37798 14000
rect 38470 13988 38476 14000
rect 37792 13960 38476 13988
rect 37792 13948 37798 13960
rect 38470 13948 38476 13960
rect 38528 13988 38534 14000
rect 38838 13988 38844 14000
rect 38528 13960 38654 13988
rect 38799 13960 38844 13988
rect 38528 13948 38534 13960
rect 22189 13923 22247 13929
rect 22189 13889 22201 13923
rect 22235 13889 22247 13923
rect 22189 13883 22247 13889
rect 22278 13880 22284 13932
rect 22336 13920 22342 13932
rect 22445 13923 22503 13929
rect 22445 13920 22457 13923
rect 22336 13892 22457 13920
rect 22336 13880 22342 13892
rect 22445 13889 22457 13892
rect 22491 13889 22503 13923
rect 22445 13883 22503 13889
rect 26329 13923 26387 13929
rect 26329 13889 26341 13923
rect 26375 13920 26387 13923
rect 26418 13920 26424 13932
rect 26375 13892 26424 13920
rect 26375 13889 26387 13892
rect 26329 13883 26387 13889
rect 26418 13880 26424 13892
rect 26476 13880 26482 13932
rect 27522 13880 27528 13932
rect 27580 13920 27586 13932
rect 28261 13923 28319 13929
rect 28261 13920 28273 13923
rect 27580 13892 28273 13920
rect 27580 13880 27586 13892
rect 28261 13889 28273 13892
rect 28307 13889 28319 13923
rect 28261 13883 28319 13889
rect 28350 13880 28356 13932
rect 28408 13920 28414 13932
rect 28528 13923 28586 13929
rect 28528 13920 28540 13923
rect 28408 13892 28540 13920
rect 28408 13880 28414 13892
rect 28528 13889 28540 13892
rect 28574 13920 28586 13923
rect 30190 13920 30196 13932
rect 28574 13892 30196 13920
rect 28574 13889 28586 13892
rect 28528 13883 28586 13889
rect 30190 13880 30196 13892
rect 30248 13880 30254 13932
rect 31214 13923 31272 13929
rect 31214 13920 31226 13923
rect 30300 13892 31226 13920
rect 19337 13855 19395 13861
rect 19116 13824 19161 13852
rect 19116 13812 19122 13824
rect 19337 13821 19349 13855
rect 19383 13852 19395 13855
rect 22094 13852 22100 13864
rect 19383 13824 22100 13852
rect 19383 13821 19395 13824
rect 19337 13815 19395 13821
rect 22094 13812 22100 13824
rect 22152 13812 22158 13864
rect 29270 13812 29276 13864
rect 29328 13852 29334 13864
rect 30300 13852 30328 13892
rect 31214 13889 31226 13892
rect 31260 13889 31272 13923
rect 32214 13920 32220 13932
rect 32175 13892 32220 13920
rect 31214 13883 31272 13889
rect 32214 13880 32220 13892
rect 32272 13880 32278 13932
rect 32306 13880 32312 13932
rect 32364 13920 32370 13932
rect 32401 13923 32459 13929
rect 32401 13920 32413 13923
rect 32364 13892 32413 13920
rect 32364 13880 32370 13892
rect 32401 13889 32413 13892
rect 32447 13889 32459 13923
rect 32401 13883 32459 13889
rect 35713 13923 35771 13929
rect 35713 13889 35725 13923
rect 35759 13920 35771 13923
rect 35802 13920 35808 13932
rect 35759 13892 35808 13920
rect 35759 13889 35771 13892
rect 35713 13883 35771 13889
rect 35802 13880 35808 13892
rect 35860 13920 35866 13932
rect 37366 13920 37372 13932
rect 35860 13892 37372 13920
rect 35860 13880 35866 13892
rect 37366 13880 37372 13892
rect 37424 13920 37430 13932
rect 38197 13923 38255 13929
rect 38197 13920 38209 13923
rect 37424 13892 38209 13920
rect 37424 13880 37430 13892
rect 38197 13889 38209 13892
rect 38243 13889 38255 13923
rect 38626 13920 38654 13960
rect 38838 13948 38844 13960
rect 38896 13948 38902 14000
rect 39592 13929 39620 14028
rect 39117 13923 39175 13929
rect 39117 13920 39129 13923
rect 38626 13892 39129 13920
rect 38197 13883 38255 13889
rect 39117 13889 39129 13892
rect 39163 13889 39175 13923
rect 39117 13883 39175 13889
rect 39577 13923 39635 13929
rect 39577 13889 39589 13923
rect 39623 13889 39635 13923
rect 39577 13883 39635 13889
rect 39761 13923 39819 13929
rect 39761 13889 39773 13923
rect 39807 13889 39819 13923
rect 39761 13883 39819 13889
rect 43625 13923 43683 13929
rect 43625 13889 43637 13923
rect 43671 13920 43683 13923
rect 43714 13920 43720 13932
rect 43671 13892 43720 13920
rect 43671 13889 43683 13892
rect 43625 13883 43683 13889
rect 31478 13852 31484 13864
rect 29328 13824 30328 13852
rect 31439 13824 31484 13852
rect 29328 13812 29334 13824
rect 31478 13812 31484 13824
rect 31536 13812 31542 13864
rect 33502 13812 33508 13864
rect 33560 13852 33566 13864
rect 34422 13852 34428 13864
rect 33560 13824 34428 13852
rect 33560 13812 33566 13824
rect 34422 13812 34428 13824
rect 34480 13852 34486 13864
rect 34517 13855 34575 13861
rect 34517 13852 34529 13855
rect 34480 13824 34529 13852
rect 34480 13812 34486 13824
rect 34517 13821 34529 13824
rect 34563 13821 34575 13855
rect 34517 13815 34575 13821
rect 35989 13855 36047 13861
rect 35989 13821 36001 13855
rect 36035 13852 36047 13855
rect 36446 13852 36452 13864
rect 36035 13824 36452 13852
rect 36035 13821 36047 13824
rect 35989 13815 36047 13821
rect 36446 13812 36452 13824
rect 36504 13852 36510 13864
rect 37090 13852 37096 13864
rect 36504 13824 37096 13852
rect 36504 13812 36510 13824
rect 37090 13812 37096 13824
rect 37148 13812 37154 13864
rect 37550 13812 37556 13864
rect 37608 13852 37614 13864
rect 38841 13855 38899 13861
rect 38841 13852 38853 13855
rect 37608 13824 38853 13852
rect 37608 13812 37614 13824
rect 38841 13821 38853 13824
rect 38887 13852 38899 13855
rect 39132 13852 39160 13883
rect 39776 13852 39804 13883
rect 43714 13880 43720 13892
rect 43772 13880 43778 13932
rect 38887 13824 38976 13852
rect 39132 13824 39804 13852
rect 38887 13821 38899 13824
rect 38841 13815 38899 13821
rect 18049 13787 18107 13793
rect 18049 13753 18061 13787
rect 18095 13753 18107 13787
rect 18049 13747 18107 13753
rect 24578 13744 24584 13796
rect 24636 13784 24642 13796
rect 25498 13784 25504 13796
rect 24636 13756 25504 13784
rect 24636 13744 24642 13756
rect 25498 13744 25504 13756
rect 25556 13744 25562 13796
rect 27522 13784 27528 13796
rect 27483 13756 27528 13784
rect 27522 13744 27528 13756
rect 27580 13744 27586 13796
rect 19242 13676 19248 13728
rect 19300 13716 19306 13728
rect 20165 13719 20223 13725
rect 20165 13716 20177 13719
rect 19300 13688 20177 13716
rect 19300 13676 19306 13688
rect 20165 13685 20177 13688
rect 20211 13685 20223 13719
rect 20165 13679 20223 13685
rect 27798 13676 27804 13728
rect 27856 13716 27862 13728
rect 29288 13716 29316 13812
rect 33962 13716 33968 13728
rect 27856 13688 29316 13716
rect 33923 13688 33968 13716
rect 27856 13676 27862 13688
rect 33962 13676 33968 13688
rect 34020 13676 34026 13728
rect 37274 13716 37280 13728
rect 37235 13688 37280 13716
rect 37274 13676 37280 13688
rect 37332 13676 37338 13728
rect 37458 13716 37464 13728
rect 37419 13688 37464 13716
rect 37458 13676 37464 13688
rect 37516 13676 37522 13728
rect 38286 13716 38292 13728
rect 38247 13688 38292 13716
rect 38286 13676 38292 13688
rect 38344 13676 38350 13728
rect 38948 13716 38976 13824
rect 39025 13787 39083 13793
rect 39025 13753 39037 13787
rect 39071 13784 39083 13787
rect 39114 13784 39120 13796
rect 39071 13756 39120 13784
rect 39071 13753 39083 13756
rect 39025 13747 39083 13753
rect 39114 13744 39120 13756
rect 39172 13744 39178 13796
rect 39669 13719 39727 13725
rect 39669 13716 39681 13719
rect 38948 13688 39681 13716
rect 39669 13685 39681 13688
rect 39715 13685 39727 13719
rect 42794 13716 42800 13728
rect 42755 13688 42800 13716
rect 39669 13679 39727 13685
rect 42794 13676 42800 13688
rect 42852 13676 42858 13728
rect 43530 13716 43536 13728
rect 43491 13688 43536 13716
rect 43530 13676 43536 13688
rect 43588 13676 43594 13728
rect 1104 13626 44896 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 44896 13626
rect 1104 13552 44896 13574
rect 16853 13515 16911 13521
rect 16853 13481 16865 13515
rect 16899 13512 16911 13515
rect 16942 13512 16948 13524
rect 16899 13484 16948 13512
rect 16899 13481 16911 13484
rect 16853 13475 16911 13481
rect 16942 13472 16948 13484
rect 17000 13472 17006 13524
rect 18046 13512 18052 13524
rect 18007 13484 18052 13512
rect 18046 13472 18052 13484
rect 18104 13472 18110 13524
rect 18509 13515 18567 13521
rect 18509 13481 18521 13515
rect 18555 13512 18567 13515
rect 18782 13512 18788 13524
rect 18555 13484 18788 13512
rect 18555 13481 18567 13484
rect 18509 13475 18567 13481
rect 18782 13472 18788 13484
rect 18840 13472 18846 13524
rect 21361 13515 21419 13521
rect 21361 13481 21373 13515
rect 21407 13512 21419 13515
rect 22278 13512 22284 13524
rect 21407 13484 22284 13512
rect 21407 13481 21419 13484
rect 21361 13475 21419 13481
rect 22278 13472 22284 13484
rect 22336 13472 22342 13524
rect 25682 13472 25688 13524
rect 25740 13512 25746 13524
rect 25777 13515 25835 13521
rect 25777 13512 25789 13515
rect 25740 13484 25789 13512
rect 25740 13472 25746 13484
rect 25777 13481 25789 13484
rect 25823 13481 25835 13515
rect 25777 13475 25835 13481
rect 36725 13515 36783 13521
rect 36725 13481 36737 13515
rect 36771 13512 36783 13515
rect 38286 13512 38292 13524
rect 36771 13484 38292 13512
rect 36771 13481 36783 13484
rect 36725 13475 36783 13481
rect 38286 13472 38292 13484
rect 38344 13472 38350 13524
rect 38930 13512 38936 13524
rect 38891 13484 38936 13512
rect 38930 13472 38936 13484
rect 38988 13472 38994 13524
rect 17218 13404 17224 13456
rect 17276 13444 17282 13456
rect 17313 13447 17371 13453
rect 17313 13444 17325 13447
rect 17276 13416 17325 13444
rect 17276 13404 17282 13416
rect 17313 13413 17325 13416
rect 17359 13413 17371 13447
rect 19058 13444 19064 13456
rect 17313 13407 17371 13413
rect 18248 13416 19064 13444
rect 1670 13268 1676 13320
rect 1728 13308 1734 13320
rect 1765 13311 1823 13317
rect 1765 13308 1777 13311
rect 1728 13280 1777 13308
rect 1728 13268 1734 13280
rect 1765 13277 1777 13280
rect 1811 13277 1823 13311
rect 1765 13271 1823 13277
rect 16669 13311 16727 13317
rect 16669 13277 16681 13311
rect 16715 13308 16727 13311
rect 17954 13308 17960 13320
rect 16715 13280 17960 13308
rect 16715 13277 16727 13280
rect 16669 13271 16727 13277
rect 17954 13268 17960 13280
rect 18012 13268 18018 13320
rect 18248 13317 18276 13416
rect 19058 13404 19064 13416
rect 19116 13404 19122 13456
rect 21910 13404 21916 13456
rect 21968 13444 21974 13456
rect 21968 13416 22094 13444
rect 21968 13404 21974 13416
rect 18414 13376 18420 13388
rect 18375 13348 18420 13376
rect 18414 13336 18420 13348
rect 18472 13336 18478 13388
rect 21821 13379 21879 13385
rect 21821 13376 21833 13379
rect 20916 13348 21833 13376
rect 20916 13320 20944 13348
rect 21821 13345 21833 13348
rect 21867 13345 21879 13379
rect 22066 13376 22094 13416
rect 23017 13379 23075 13385
rect 23017 13376 23029 13379
rect 22066 13348 23029 13376
rect 21821 13339 21879 13345
rect 18233 13311 18291 13317
rect 18233 13277 18245 13311
rect 18279 13277 18291 13311
rect 19242 13308 19248 13320
rect 18233 13271 18291 13277
rect 18340 13280 19248 13308
rect 17497 13243 17555 13249
rect 17497 13209 17509 13243
rect 17543 13240 17555 13243
rect 18340 13240 18368 13280
rect 19242 13268 19248 13280
rect 19300 13308 19306 13320
rect 19705 13311 19763 13317
rect 19705 13308 19717 13311
rect 19300 13280 19717 13308
rect 19300 13268 19306 13280
rect 19705 13277 19717 13280
rect 19751 13277 19763 13311
rect 19705 13271 19763 13277
rect 19981 13311 20039 13317
rect 19981 13277 19993 13311
rect 20027 13308 20039 13311
rect 20898 13308 20904 13320
rect 20027 13280 20904 13308
rect 20027 13277 20039 13280
rect 19981 13271 20039 13277
rect 20898 13268 20904 13280
rect 20956 13268 20962 13320
rect 20990 13268 20996 13320
rect 21048 13308 21054 13320
rect 21085 13311 21143 13317
rect 21085 13308 21097 13311
rect 21048 13280 21097 13308
rect 21048 13268 21054 13280
rect 21085 13277 21097 13280
rect 21131 13308 21143 13311
rect 21910 13308 21916 13320
rect 21131 13280 21916 13308
rect 21131 13277 21143 13280
rect 21085 13271 21143 13277
rect 21910 13268 21916 13280
rect 21968 13308 21974 13320
rect 22112 13317 22140 13348
rect 23017 13345 23029 13348
rect 23063 13345 23075 13379
rect 23017 13339 23075 13345
rect 36541 13379 36599 13385
rect 36541 13345 36553 13379
rect 36587 13376 36599 13379
rect 38010 13376 38016 13388
rect 36587 13348 38016 13376
rect 36587 13345 36599 13348
rect 36541 13339 36599 13345
rect 38010 13336 38016 13348
rect 38068 13336 38074 13388
rect 42337 13379 42395 13385
rect 42337 13345 42349 13379
rect 42383 13376 42395 13379
rect 42794 13376 42800 13388
rect 42383 13348 42800 13376
rect 42383 13345 42395 13348
rect 42337 13339 42395 13345
rect 42794 13336 42800 13348
rect 42852 13336 42858 13388
rect 44082 13376 44088 13388
rect 44043 13348 44088 13376
rect 44082 13336 44088 13348
rect 44140 13336 44146 13388
rect 22005 13311 22063 13317
rect 22005 13308 22017 13311
rect 21968 13280 22017 13308
rect 21968 13268 21974 13280
rect 22005 13277 22017 13280
rect 22051 13277 22063 13311
rect 22005 13271 22063 13277
rect 22097 13311 22155 13317
rect 22097 13277 22109 13311
rect 22143 13277 22155 13311
rect 22097 13271 22155 13277
rect 22646 13268 22652 13320
rect 22704 13308 22710 13320
rect 22741 13311 22799 13317
rect 22741 13308 22753 13311
rect 22704 13280 22753 13308
rect 22704 13268 22710 13280
rect 22741 13277 22753 13280
rect 22787 13277 22799 13311
rect 24394 13308 24400 13320
rect 24355 13280 24400 13308
rect 22741 13271 22799 13277
rect 24394 13268 24400 13280
rect 24452 13268 24458 13320
rect 32493 13311 32551 13317
rect 32493 13277 32505 13311
rect 32539 13308 32551 13311
rect 33962 13308 33968 13320
rect 32539 13280 33968 13308
rect 32539 13277 32551 13280
rect 32493 13271 32551 13277
rect 33962 13268 33968 13280
rect 34020 13268 34026 13320
rect 36817 13311 36875 13317
rect 36817 13277 36829 13311
rect 36863 13277 36875 13311
rect 36817 13271 36875 13277
rect 18506 13240 18512 13252
rect 17543 13212 18368 13240
rect 18467 13212 18512 13240
rect 17543 13209 17555 13212
rect 17497 13203 17555 13209
rect 18506 13200 18512 13212
rect 18564 13200 18570 13252
rect 24670 13249 24676 13252
rect 21361 13243 21419 13249
rect 21361 13209 21373 13243
rect 21407 13240 21419 13243
rect 21821 13243 21879 13249
rect 21821 13240 21833 13243
rect 21407 13212 21833 13240
rect 21407 13209 21419 13212
rect 21361 13203 21419 13209
rect 21821 13209 21833 13212
rect 21867 13209 21879 13243
rect 21821 13203 21879 13209
rect 24664 13203 24676 13249
rect 24728 13240 24734 13252
rect 36832 13240 36860 13271
rect 37366 13268 37372 13320
rect 37424 13308 37430 13320
rect 37461 13311 37519 13317
rect 37461 13308 37473 13311
rect 37424 13280 37473 13308
rect 37424 13268 37430 13280
rect 37461 13277 37473 13280
rect 37507 13277 37519 13311
rect 37642 13308 37648 13320
rect 37603 13280 37648 13308
rect 37461 13271 37519 13277
rect 37642 13268 37648 13280
rect 37700 13268 37706 13320
rect 37737 13311 37795 13317
rect 37737 13277 37749 13311
rect 37783 13277 37795 13311
rect 37737 13271 37795 13277
rect 37660 13240 37688 13268
rect 24728 13212 24764 13240
rect 36832 13212 37688 13240
rect 37752 13240 37780 13271
rect 37826 13268 37832 13320
rect 37884 13308 37890 13320
rect 39114 13308 39120 13320
rect 37884 13280 37929 13308
rect 38028 13280 39120 13308
rect 37884 13268 37890 13280
rect 38028 13240 38056 13280
rect 39114 13268 39120 13280
rect 39172 13268 39178 13320
rect 37752 13212 38056 13240
rect 24670 13200 24676 13203
rect 24728 13200 24734 13212
rect 38194 13200 38200 13252
rect 38252 13240 38258 13252
rect 38562 13240 38568 13252
rect 38252 13212 38568 13240
rect 38252 13200 38258 13212
rect 38562 13200 38568 13212
rect 38620 13200 38626 13252
rect 38654 13200 38660 13252
rect 38712 13240 38718 13252
rect 38749 13243 38807 13249
rect 38749 13240 38761 13243
rect 38712 13212 38761 13240
rect 38712 13200 38718 13212
rect 38749 13209 38761 13212
rect 38795 13209 38807 13243
rect 38749 13203 38807 13209
rect 42521 13243 42579 13249
rect 42521 13209 42533 13243
rect 42567 13240 42579 13243
rect 43530 13240 43536 13252
rect 42567 13212 43536 13240
rect 42567 13209 42579 13212
rect 42521 13203 42579 13209
rect 43530 13200 43536 13212
rect 43588 13200 43594 13252
rect 21177 13175 21235 13181
rect 21177 13141 21189 13175
rect 21223 13172 21235 13175
rect 21726 13172 21732 13184
rect 21223 13144 21732 13172
rect 21223 13141 21235 13144
rect 21177 13135 21235 13141
rect 21726 13132 21732 13144
rect 21784 13132 21790 13184
rect 32674 13172 32680 13184
rect 32635 13144 32680 13172
rect 32674 13132 32680 13144
rect 32732 13132 32738 13184
rect 36078 13132 36084 13184
rect 36136 13172 36142 13184
rect 36265 13175 36323 13181
rect 36265 13172 36277 13175
rect 36136 13144 36277 13172
rect 36136 13132 36142 13144
rect 36265 13141 36277 13144
rect 36311 13141 36323 13175
rect 38102 13172 38108 13184
rect 38063 13144 38108 13172
rect 36265 13135 36323 13141
rect 38102 13132 38108 13144
rect 38160 13132 38166 13184
rect 1104 13082 44896 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 44896 13082
rect 1104 13008 44896 13030
rect 18138 12928 18144 12980
rect 18196 12968 18202 12980
rect 18325 12971 18383 12977
rect 18325 12968 18337 12971
rect 18196 12940 18337 12968
rect 18196 12928 18202 12940
rect 18325 12937 18337 12940
rect 18371 12937 18383 12971
rect 18325 12931 18383 12937
rect 19426 12928 19432 12980
rect 19484 12968 19490 12980
rect 19521 12971 19579 12977
rect 19521 12968 19533 12971
rect 19484 12940 19533 12968
rect 19484 12928 19490 12940
rect 19521 12937 19533 12940
rect 19567 12937 19579 12971
rect 19521 12931 19579 12937
rect 21269 12971 21327 12977
rect 21269 12937 21281 12971
rect 21315 12968 21327 12971
rect 23845 12971 23903 12977
rect 21315 12940 22968 12968
rect 21315 12937 21327 12940
rect 21269 12931 21327 12937
rect 18690 12900 18696 12912
rect 18651 12872 18696 12900
rect 18690 12860 18696 12872
rect 18748 12860 18754 12912
rect 20714 12900 20720 12912
rect 19720 12872 20720 12900
rect 1670 12832 1676 12844
rect 1631 12804 1676 12832
rect 1670 12792 1676 12804
rect 1728 12792 1734 12844
rect 9214 12832 9220 12844
rect 9127 12804 9220 12832
rect 9214 12792 9220 12804
rect 9272 12832 9278 12844
rect 12710 12832 12716 12844
rect 9272 12804 12716 12832
rect 9272 12792 9278 12804
rect 12710 12792 12716 12804
rect 12768 12792 12774 12844
rect 18506 12832 18512 12844
rect 18419 12804 18512 12832
rect 18506 12792 18512 12804
rect 18564 12792 18570 12844
rect 19720 12841 19748 12872
rect 20714 12860 20720 12872
rect 20772 12860 20778 12912
rect 20898 12900 20904 12912
rect 20859 12872 20904 12900
rect 20898 12860 20904 12872
rect 20956 12860 20962 12912
rect 21117 12903 21175 12909
rect 21117 12869 21129 12903
rect 21163 12900 21175 12903
rect 21821 12903 21879 12909
rect 21821 12900 21833 12903
rect 21163 12872 21833 12900
rect 21163 12869 21175 12872
rect 21117 12863 21175 12869
rect 21821 12869 21833 12872
rect 21867 12869 21879 12903
rect 21821 12863 21879 12869
rect 21910 12860 21916 12912
rect 21968 12900 21974 12912
rect 21968 12872 22324 12900
rect 21968 12860 21974 12872
rect 19705 12835 19763 12841
rect 19705 12801 19717 12835
rect 19751 12801 19763 12835
rect 19705 12795 19763 12801
rect 19886 12792 19892 12844
rect 19944 12832 19950 12844
rect 21266 12832 21272 12844
rect 19944 12804 21272 12832
rect 19944 12792 19950 12804
rect 21266 12792 21272 12804
rect 21324 12792 21330 12844
rect 22002 12832 22008 12844
rect 21963 12804 22008 12832
rect 22002 12792 22008 12804
rect 22060 12792 22066 12844
rect 22296 12841 22324 12872
rect 22940 12841 22968 12940
rect 23845 12937 23857 12971
rect 23891 12968 23903 12971
rect 24578 12968 24584 12980
rect 23891 12940 24584 12968
rect 23891 12937 23903 12940
rect 23845 12931 23903 12937
rect 24578 12928 24584 12940
rect 24636 12928 24642 12980
rect 25774 12968 25780 12980
rect 25735 12940 25780 12968
rect 25774 12928 25780 12940
rect 25832 12928 25838 12980
rect 27157 12971 27215 12977
rect 27157 12937 27169 12971
rect 27203 12968 27215 12971
rect 27430 12968 27436 12980
rect 27203 12940 27436 12968
rect 27203 12937 27215 12940
rect 27157 12931 27215 12937
rect 27430 12928 27436 12940
rect 27488 12928 27494 12980
rect 36078 12968 36084 12980
rect 36039 12940 36084 12968
rect 36078 12928 36084 12940
rect 36136 12928 36142 12980
rect 37826 12928 37832 12980
rect 37884 12968 37890 12980
rect 39117 12971 39175 12977
rect 39117 12968 39129 12971
rect 37884 12940 39129 12968
rect 37884 12928 37890 12940
rect 39117 12937 39129 12940
rect 39163 12937 39175 12971
rect 39117 12931 39175 12937
rect 27249 12903 27307 12909
rect 27249 12869 27261 12903
rect 27295 12900 27307 12903
rect 27522 12900 27528 12912
rect 27295 12872 27528 12900
rect 27295 12869 27307 12872
rect 27249 12863 27307 12869
rect 27522 12860 27528 12872
rect 27580 12900 27586 12912
rect 31021 12903 31079 12909
rect 31021 12900 31033 12903
rect 27580 12872 31033 12900
rect 27580 12860 27586 12872
rect 31021 12869 31033 12872
rect 31067 12869 31079 12903
rect 31021 12863 31079 12869
rect 31110 12860 31116 12912
rect 31168 12900 31174 12912
rect 31205 12903 31263 12909
rect 31205 12900 31217 12903
rect 31168 12872 31217 12900
rect 31168 12860 31174 12872
rect 31205 12869 31217 12872
rect 31251 12900 31263 12903
rect 31478 12900 31484 12912
rect 31251 12872 31484 12900
rect 31251 12869 31263 12872
rect 31205 12863 31263 12869
rect 31478 12860 31484 12872
rect 31536 12900 31542 12912
rect 31536 12872 33548 12900
rect 31536 12860 31542 12872
rect 33520 12844 33548 12872
rect 38654 12860 38660 12912
rect 38712 12900 38718 12912
rect 41693 12903 41751 12909
rect 38712 12872 39252 12900
rect 38712 12860 38718 12872
rect 22189 12835 22247 12841
rect 22189 12801 22201 12835
rect 22235 12801 22247 12835
rect 22189 12795 22247 12801
rect 22281 12835 22339 12841
rect 22281 12801 22293 12835
rect 22327 12801 22339 12835
rect 22281 12795 22339 12801
rect 22925 12835 22983 12841
rect 22925 12801 22937 12835
rect 22971 12801 22983 12835
rect 23658 12832 23664 12844
rect 23619 12804 23664 12832
rect 22925 12795 22983 12801
rect 1854 12764 1860 12776
rect 1815 12736 1860 12764
rect 1854 12724 1860 12736
rect 1912 12724 1918 12776
rect 2774 12764 2780 12776
rect 2735 12736 2780 12764
rect 2774 12724 2780 12736
rect 2832 12724 2838 12776
rect 18524 12696 18552 12792
rect 18690 12724 18696 12776
rect 18748 12764 18754 12776
rect 19904 12764 19932 12792
rect 18748 12736 19932 12764
rect 18748 12724 18754 12736
rect 21818 12724 21824 12776
rect 21876 12764 21882 12776
rect 22204 12764 22232 12795
rect 23658 12792 23664 12804
rect 23716 12792 23722 12844
rect 23842 12792 23848 12844
rect 23900 12832 23906 12844
rect 24653 12835 24711 12841
rect 24653 12832 24665 12835
rect 23900 12804 24665 12832
rect 23900 12792 23906 12804
rect 24653 12801 24665 12804
rect 24699 12801 24711 12835
rect 27798 12832 27804 12844
rect 27759 12804 27804 12832
rect 24653 12795 24711 12801
rect 27798 12792 27804 12804
rect 27856 12792 27862 12844
rect 27982 12832 27988 12844
rect 27943 12804 27988 12832
rect 27982 12792 27988 12804
rect 28040 12792 28046 12844
rect 28169 12835 28227 12841
rect 28169 12801 28181 12835
rect 28215 12832 28227 12835
rect 28629 12835 28687 12841
rect 28629 12832 28641 12835
rect 28215 12804 28641 12832
rect 28215 12801 28227 12804
rect 28169 12795 28227 12801
rect 28629 12801 28641 12804
rect 28675 12801 28687 12835
rect 29822 12832 29828 12844
rect 29783 12804 29828 12832
rect 28629 12795 28687 12801
rect 29822 12792 29828 12804
rect 29880 12792 29886 12844
rect 32674 12792 32680 12844
rect 32732 12832 32738 12844
rect 33238 12835 33296 12841
rect 33238 12832 33250 12835
rect 32732 12804 33250 12832
rect 32732 12792 32738 12804
rect 33238 12801 33250 12804
rect 33284 12801 33296 12835
rect 33502 12832 33508 12844
rect 33415 12804 33508 12832
rect 33238 12795 33296 12801
rect 33502 12792 33508 12804
rect 33560 12792 33566 12844
rect 35621 12835 35679 12841
rect 35621 12801 35633 12835
rect 35667 12832 35679 12835
rect 36538 12832 36544 12844
rect 35667 12804 36544 12832
rect 35667 12801 35679 12804
rect 35621 12795 35679 12801
rect 36538 12792 36544 12804
rect 36596 12792 36602 12844
rect 38010 12792 38016 12844
rect 38068 12832 38074 12844
rect 38194 12832 38200 12844
rect 38068 12804 38200 12832
rect 38068 12792 38074 12804
rect 38194 12792 38200 12804
rect 38252 12832 38258 12844
rect 39224 12841 39252 12872
rect 41693 12869 41705 12903
rect 41739 12900 41751 12903
rect 43533 12903 43591 12909
rect 43533 12900 43545 12903
rect 41739 12872 43545 12900
rect 41739 12869 41751 12872
rect 41693 12863 41751 12869
rect 43533 12869 43545 12872
rect 43579 12869 43591 12903
rect 43533 12863 43591 12869
rect 38289 12835 38347 12841
rect 38289 12832 38301 12835
rect 38252 12804 38301 12832
rect 38252 12792 38258 12804
rect 38289 12801 38301 12804
rect 38335 12832 38347 12835
rect 39025 12835 39083 12841
rect 39025 12832 39037 12835
rect 38335 12804 39037 12832
rect 38335 12801 38347 12804
rect 38289 12795 38347 12801
rect 39025 12801 39037 12804
rect 39071 12801 39083 12835
rect 39025 12795 39083 12801
rect 39209 12835 39267 12841
rect 39209 12801 39221 12835
rect 39255 12801 39267 12835
rect 39209 12795 39267 12801
rect 43625 12835 43683 12841
rect 43625 12801 43637 12835
rect 43671 12832 43683 12835
rect 43714 12832 43720 12844
rect 43671 12804 43720 12832
rect 43671 12801 43683 12804
rect 43625 12795 43683 12801
rect 43714 12792 43720 12804
rect 43772 12792 43778 12844
rect 24394 12764 24400 12776
rect 21876 12736 22232 12764
rect 24307 12736 24400 12764
rect 21876 12724 21882 12736
rect 24394 12724 24400 12736
rect 24452 12724 24458 12776
rect 34422 12724 34428 12776
rect 34480 12764 34486 12776
rect 35710 12764 35716 12776
rect 34480 12736 35716 12764
rect 34480 12724 34486 12736
rect 35710 12724 35716 12736
rect 35768 12724 35774 12776
rect 38562 12764 38568 12776
rect 38523 12736 38568 12764
rect 38562 12724 38568 12736
rect 38620 12724 38626 12776
rect 41325 12767 41383 12773
rect 41325 12733 41337 12767
rect 41371 12764 41383 12767
rect 41414 12764 41420 12776
rect 41371 12736 41420 12764
rect 41371 12733 41383 12736
rect 41325 12727 41383 12733
rect 41414 12724 41420 12736
rect 41472 12724 41478 12776
rect 41877 12767 41935 12773
rect 41877 12733 41889 12767
rect 41923 12764 41935 12767
rect 42797 12767 42855 12773
rect 42797 12764 42809 12767
rect 41923 12736 42809 12764
rect 41923 12733 41935 12736
rect 41877 12727 41935 12733
rect 42797 12733 42809 12736
rect 42843 12733 42855 12767
rect 42797 12727 42855 12733
rect 23290 12696 23296 12708
rect 18524 12668 23296 12696
rect 23290 12656 23296 12668
rect 23348 12656 23354 12708
rect 9309 12631 9367 12637
rect 9309 12597 9321 12631
rect 9355 12628 9367 12631
rect 9398 12628 9404 12640
rect 9355 12600 9404 12628
rect 9355 12597 9367 12600
rect 9309 12591 9367 12597
rect 9398 12588 9404 12600
rect 9456 12588 9462 12640
rect 21082 12628 21088 12640
rect 21043 12600 21088 12628
rect 21082 12588 21088 12600
rect 21140 12588 21146 12640
rect 22646 12588 22652 12640
rect 22704 12628 22710 12640
rect 22741 12631 22799 12637
rect 22741 12628 22753 12631
rect 22704 12600 22753 12628
rect 22704 12588 22710 12600
rect 22741 12597 22753 12600
rect 22787 12597 22799 12631
rect 24412 12628 24440 12724
rect 24762 12628 24768 12640
rect 24412 12600 24768 12628
rect 22741 12591 22799 12597
rect 24762 12588 24768 12600
rect 24820 12588 24826 12640
rect 28810 12628 28816 12640
rect 28771 12600 28816 12628
rect 28810 12588 28816 12600
rect 28868 12588 28874 12640
rect 30466 12628 30472 12640
rect 30427 12600 30472 12628
rect 30466 12588 30472 12600
rect 30524 12588 30530 12640
rect 32122 12628 32128 12640
rect 32083 12600 32128 12628
rect 32122 12588 32128 12600
rect 32180 12588 32186 12640
rect 35434 12628 35440 12640
rect 35395 12600 35440 12628
rect 35434 12588 35440 12600
rect 35492 12588 35498 12640
rect 1104 12538 44896 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 44896 12538
rect 1104 12464 44896 12486
rect 1854 12384 1860 12436
rect 1912 12424 1918 12436
rect 2225 12427 2283 12433
rect 2225 12424 2237 12427
rect 1912 12396 2237 12424
rect 1912 12384 1918 12396
rect 2225 12393 2237 12396
rect 2271 12393 2283 12427
rect 18414 12424 18420 12436
rect 18375 12396 18420 12424
rect 2225 12387 2283 12393
rect 18414 12384 18420 12396
rect 18472 12384 18478 12436
rect 21545 12427 21603 12433
rect 21545 12393 21557 12427
rect 21591 12424 21603 12427
rect 22002 12424 22008 12436
rect 21591 12396 22008 12424
rect 21591 12393 21603 12396
rect 21545 12387 21603 12393
rect 22002 12384 22008 12396
rect 22060 12384 22066 12436
rect 23842 12424 23848 12436
rect 23803 12396 23848 12424
rect 23842 12384 23848 12396
rect 23900 12384 23906 12436
rect 38930 12356 38936 12368
rect 37844 12328 38936 12356
rect 19886 12288 19892 12300
rect 19847 12260 19892 12288
rect 19886 12248 19892 12260
rect 19944 12248 19950 12300
rect 20165 12291 20223 12297
rect 20165 12257 20177 12291
rect 20211 12288 20223 12291
rect 20806 12288 20812 12300
rect 20211 12260 20812 12288
rect 20211 12257 20223 12260
rect 20165 12251 20223 12257
rect 20806 12248 20812 12260
rect 20864 12248 20870 12300
rect 24578 12288 24584 12300
rect 24539 12260 24584 12288
rect 24578 12248 24584 12260
rect 24636 12248 24642 12300
rect 32122 12248 32128 12300
rect 32180 12288 32186 12300
rect 32217 12291 32275 12297
rect 32217 12288 32229 12291
rect 32180 12260 32229 12288
rect 32180 12248 32186 12260
rect 32217 12257 32229 12260
rect 32263 12257 32275 12291
rect 32217 12251 32275 12257
rect 32306 12248 32312 12300
rect 32364 12288 32370 12300
rect 35342 12288 35348 12300
rect 32364 12260 32409 12288
rect 35303 12260 35348 12288
rect 32364 12248 32370 12260
rect 35342 12248 35348 12260
rect 35400 12288 35406 12300
rect 37844 12297 37872 12328
rect 38930 12316 38936 12328
rect 38988 12316 38994 12368
rect 36449 12291 36507 12297
rect 36449 12288 36461 12291
rect 35400 12260 36461 12288
rect 35400 12248 35406 12260
rect 36449 12257 36461 12260
rect 36495 12257 36507 12291
rect 36449 12251 36507 12257
rect 37829 12291 37887 12297
rect 37829 12257 37841 12291
rect 37875 12257 37887 12291
rect 37829 12251 37887 12257
rect 38013 12291 38071 12297
rect 38013 12257 38025 12291
rect 38059 12288 38071 12291
rect 38286 12288 38292 12300
rect 38059 12260 38292 12288
rect 38059 12257 38071 12260
rect 38013 12251 38071 12257
rect 38286 12248 38292 12260
rect 38344 12288 38350 12300
rect 42702 12288 42708 12300
rect 38344 12260 38792 12288
rect 42663 12260 42708 12288
rect 38344 12248 38350 12260
rect 2317 12223 2375 12229
rect 2317 12189 2329 12223
rect 2363 12220 2375 12223
rect 4890 12220 4896 12232
rect 2363 12192 4896 12220
rect 2363 12189 2375 12192
rect 2317 12183 2375 12189
rect 4890 12180 4896 12192
rect 4948 12180 4954 12232
rect 17862 12180 17868 12232
rect 17920 12220 17926 12232
rect 18141 12223 18199 12229
rect 18141 12220 18153 12223
rect 17920 12192 18153 12220
rect 17920 12180 17926 12192
rect 18141 12189 18153 12192
rect 18187 12189 18199 12223
rect 18141 12183 18199 12189
rect 22646 12180 22652 12232
rect 22704 12229 22710 12232
rect 22704 12220 22716 12229
rect 22704 12192 22749 12220
rect 22704 12183 22716 12192
rect 22704 12180 22710 12183
rect 22830 12180 22836 12232
rect 22888 12220 22894 12232
rect 22925 12223 22983 12229
rect 22925 12220 22937 12223
rect 22888 12192 22937 12220
rect 22888 12180 22894 12192
rect 22925 12189 22937 12192
rect 22971 12189 22983 12223
rect 23658 12220 23664 12232
rect 23619 12192 23664 12220
rect 22925 12183 22983 12189
rect 23658 12180 23664 12192
rect 23716 12180 23722 12232
rect 24765 12223 24823 12229
rect 24765 12220 24777 12223
rect 23768 12192 24777 12220
rect 18322 12112 18328 12164
rect 18380 12152 18386 12164
rect 18417 12155 18475 12161
rect 18417 12152 18429 12155
rect 18380 12124 18429 12152
rect 18380 12112 18386 12124
rect 18417 12121 18429 12124
rect 18463 12152 18475 12155
rect 21634 12152 21640 12164
rect 18463 12124 21640 12152
rect 18463 12121 18475 12124
rect 18417 12115 18475 12121
rect 21634 12112 21640 12124
rect 21692 12152 21698 12164
rect 23768 12152 23796 12192
rect 24765 12189 24777 12192
rect 24811 12189 24823 12223
rect 24765 12183 24823 12189
rect 25409 12223 25467 12229
rect 25409 12189 25421 12223
rect 25455 12220 25467 12223
rect 27249 12223 27307 12229
rect 27249 12220 27261 12223
rect 25455 12192 27261 12220
rect 25455 12189 25467 12192
rect 25409 12183 25467 12189
rect 27249 12189 27261 12192
rect 27295 12220 27307 12223
rect 27338 12220 27344 12232
rect 27295 12192 27344 12220
rect 27295 12189 27307 12192
rect 27249 12183 27307 12189
rect 25424 12152 25452 12183
rect 27338 12180 27344 12192
rect 27396 12180 27402 12232
rect 27516 12223 27574 12229
rect 27516 12220 27528 12223
rect 27448 12192 27528 12220
rect 25682 12161 25688 12164
rect 21692 12124 23796 12152
rect 24780 12124 25452 12152
rect 21692 12112 21698 12124
rect 24780 12096 24808 12124
rect 25676 12115 25688 12161
rect 25740 12152 25746 12164
rect 25740 12124 25776 12152
rect 25682 12112 25688 12115
rect 25740 12112 25746 12124
rect 18233 12087 18291 12093
rect 18233 12053 18245 12087
rect 18279 12084 18291 12087
rect 18598 12084 18604 12096
rect 18279 12056 18604 12084
rect 18279 12053 18291 12056
rect 18233 12047 18291 12053
rect 18598 12044 18604 12056
rect 18656 12044 18662 12096
rect 24762 12044 24768 12096
rect 24820 12044 24826 12096
rect 24949 12087 25007 12093
rect 24949 12053 24961 12087
rect 24995 12084 25007 12087
rect 25866 12084 25872 12096
rect 24995 12056 25872 12084
rect 24995 12053 25007 12056
rect 24949 12047 25007 12053
rect 25866 12044 25872 12056
rect 25924 12044 25930 12096
rect 26789 12087 26847 12093
rect 26789 12053 26801 12087
rect 26835 12084 26847 12087
rect 27448 12084 27476 12192
rect 27516 12189 27528 12192
rect 27562 12220 27574 12223
rect 27982 12220 27988 12232
rect 27562 12192 27988 12220
rect 27562 12189 27574 12192
rect 27516 12183 27574 12189
rect 27982 12180 27988 12192
rect 28040 12180 28046 12232
rect 28442 12180 28448 12232
rect 28500 12220 28506 12232
rect 29641 12223 29699 12229
rect 29641 12220 29653 12223
rect 28500 12192 29653 12220
rect 28500 12180 28506 12192
rect 29641 12189 29653 12192
rect 29687 12220 29699 12223
rect 31110 12220 31116 12232
rect 29687 12192 31116 12220
rect 29687 12189 29699 12192
rect 29641 12183 29699 12189
rect 31110 12180 31116 12192
rect 31168 12180 31174 12232
rect 33318 12220 33324 12232
rect 33279 12192 33324 12220
rect 33318 12180 33324 12192
rect 33376 12180 33382 12232
rect 33965 12223 34023 12229
rect 33965 12189 33977 12223
rect 34011 12220 34023 12223
rect 35161 12223 35219 12229
rect 34011 12192 34744 12220
rect 34011 12189 34023 12192
rect 33965 12183 34023 12189
rect 29908 12155 29966 12161
rect 29908 12121 29920 12155
rect 29954 12152 29966 12155
rect 30466 12152 30472 12164
rect 29954 12124 30472 12152
rect 29954 12121 29966 12124
rect 29908 12115 29966 12121
rect 30466 12112 30472 12124
rect 30524 12112 30530 12164
rect 31018 12084 31024 12096
rect 26835 12056 27476 12084
rect 30979 12056 31024 12084
rect 26835 12053 26847 12056
rect 26789 12047 26847 12053
rect 31018 12044 31024 12056
rect 31076 12044 31082 12096
rect 31202 12044 31208 12096
rect 31260 12084 31266 12096
rect 31757 12087 31815 12093
rect 31757 12084 31769 12087
rect 31260 12056 31769 12084
rect 31260 12044 31266 12056
rect 31757 12053 31769 12056
rect 31803 12053 31815 12087
rect 32122 12084 32128 12096
rect 32083 12056 32128 12084
rect 31757 12047 31815 12053
rect 32122 12044 32128 12056
rect 32180 12044 32186 12096
rect 33134 12084 33140 12096
rect 33095 12056 33140 12084
rect 33134 12044 33140 12056
rect 33192 12044 33198 12096
rect 33778 12084 33784 12096
rect 33739 12056 33784 12084
rect 33778 12044 33784 12056
rect 33836 12044 33842 12096
rect 34716 12093 34744 12192
rect 35161 12189 35173 12223
rect 35207 12220 35219 12223
rect 35434 12220 35440 12232
rect 35207 12192 35440 12220
rect 35207 12189 35219 12192
rect 35161 12183 35219 12189
rect 35434 12180 35440 12192
rect 35492 12180 35498 12232
rect 37642 12180 37648 12232
rect 37700 12220 37706 12232
rect 38764 12229 38792 12260
rect 42702 12248 42708 12260
rect 42760 12248 42766 12300
rect 38565 12223 38623 12229
rect 38565 12220 38577 12223
rect 37700 12192 38577 12220
rect 37700 12180 37706 12192
rect 38565 12189 38577 12192
rect 38611 12189 38623 12223
rect 38565 12183 38623 12189
rect 38749 12223 38807 12229
rect 38749 12189 38761 12223
rect 38795 12189 38807 12223
rect 38749 12183 38807 12189
rect 44174 12180 44180 12232
rect 44232 12220 44238 12232
rect 44232 12192 44277 12220
rect 44232 12180 44238 12192
rect 37737 12155 37795 12161
rect 37737 12121 37749 12155
rect 37783 12152 37795 12155
rect 38838 12152 38844 12164
rect 37783 12124 38844 12152
rect 37783 12121 37795 12124
rect 37737 12115 37795 12121
rect 38838 12112 38844 12124
rect 38896 12112 38902 12164
rect 43438 12112 43444 12164
rect 43496 12152 43502 12164
rect 43993 12155 44051 12161
rect 43993 12152 44005 12155
rect 43496 12124 44005 12152
rect 43496 12112 43502 12124
rect 43993 12121 44005 12124
rect 44039 12121 44051 12155
rect 43993 12115 44051 12121
rect 34701 12087 34759 12093
rect 34701 12053 34713 12087
rect 34747 12053 34759 12087
rect 34701 12047 34759 12053
rect 35069 12087 35127 12093
rect 35069 12053 35081 12087
rect 35115 12084 35127 12087
rect 35526 12084 35532 12096
rect 35115 12056 35532 12084
rect 35115 12053 35127 12056
rect 35069 12047 35127 12053
rect 35526 12044 35532 12056
rect 35584 12044 35590 12096
rect 35894 12044 35900 12096
rect 35952 12084 35958 12096
rect 36262 12084 36268 12096
rect 35952 12056 35997 12084
rect 36223 12056 36268 12084
rect 35952 12044 35958 12056
rect 36262 12044 36268 12056
rect 36320 12044 36326 12096
rect 36357 12087 36415 12093
rect 36357 12053 36369 12087
rect 36403 12084 36415 12087
rect 37369 12087 37427 12093
rect 37369 12084 37381 12087
rect 36403 12056 37381 12084
rect 36403 12053 36415 12056
rect 36357 12047 36415 12053
rect 37369 12053 37381 12056
rect 37415 12053 37427 12087
rect 37369 12047 37427 12053
rect 38286 12044 38292 12096
rect 38344 12084 38350 12096
rect 38657 12087 38715 12093
rect 38657 12084 38669 12087
rect 38344 12056 38669 12084
rect 38344 12044 38350 12056
rect 38657 12053 38669 12056
rect 38703 12053 38715 12087
rect 38657 12047 38715 12053
rect 1104 11994 44896 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 44896 11994
rect 1104 11920 44896 11942
rect 24581 11883 24639 11889
rect 24581 11849 24593 11883
rect 24627 11880 24639 11883
rect 24670 11880 24676 11892
rect 24627 11852 24676 11880
rect 24627 11849 24639 11852
rect 24581 11843 24639 11849
rect 24670 11840 24676 11852
rect 24728 11840 24734 11892
rect 25682 11880 25688 11892
rect 25643 11852 25688 11880
rect 25682 11840 25688 11852
rect 25740 11840 25746 11892
rect 29822 11880 29828 11892
rect 29783 11852 29828 11880
rect 29822 11840 29828 11852
rect 29880 11840 29886 11892
rect 30742 11840 30748 11892
rect 30800 11880 30806 11892
rect 30837 11883 30895 11889
rect 30837 11880 30849 11883
rect 30800 11852 30849 11880
rect 30800 11840 30806 11852
rect 30837 11849 30849 11852
rect 30883 11849 30895 11883
rect 31202 11880 31208 11892
rect 31163 11852 31208 11880
rect 30837 11843 30895 11849
rect 31202 11840 31208 11852
rect 31260 11840 31266 11892
rect 32122 11880 32128 11892
rect 32083 11852 32128 11880
rect 32122 11840 32128 11852
rect 32180 11840 32186 11892
rect 33318 11840 33324 11892
rect 33376 11880 33382 11892
rect 34333 11883 34391 11889
rect 34333 11880 34345 11883
rect 33376 11852 34345 11880
rect 33376 11840 33382 11852
rect 34333 11849 34345 11852
rect 34379 11849 34391 11883
rect 35526 11880 35532 11892
rect 35487 11852 35532 11880
rect 34333 11843 34391 11849
rect 35526 11840 35532 11852
rect 35584 11840 35590 11892
rect 35710 11880 35716 11892
rect 35671 11852 35716 11880
rect 35710 11840 35716 11852
rect 35768 11840 35774 11892
rect 36538 11840 36544 11892
rect 36596 11880 36602 11892
rect 37277 11883 37335 11889
rect 37277 11880 37289 11883
rect 36596 11852 37289 11880
rect 36596 11840 36602 11852
rect 37277 11849 37289 11852
rect 37323 11849 37335 11883
rect 43438 11880 43444 11892
rect 43399 11852 43444 11880
rect 37277 11843 37335 11849
rect 43438 11840 43444 11852
rect 43496 11840 43502 11892
rect 20254 11812 20260 11824
rect 20215 11784 20260 11812
rect 20254 11772 20260 11784
rect 20312 11772 20318 11824
rect 28712 11815 28770 11821
rect 28712 11781 28724 11815
rect 28758 11812 28770 11815
rect 28810 11812 28816 11824
rect 28758 11784 28816 11812
rect 28758 11781 28770 11784
rect 28712 11775 28770 11781
rect 28810 11772 28816 11784
rect 28868 11772 28874 11824
rect 33134 11772 33140 11824
rect 33192 11812 33198 11824
rect 33238 11815 33296 11821
rect 33238 11812 33250 11815
rect 33192 11784 33250 11812
rect 33192 11772 33198 11784
rect 33238 11781 33250 11784
rect 33284 11781 33296 11815
rect 33238 11775 33296 11781
rect 34793 11815 34851 11821
rect 34793 11781 34805 11815
rect 34839 11812 34851 11815
rect 35894 11812 35900 11824
rect 34839 11784 35900 11812
rect 34839 11781 34851 11784
rect 34793 11775 34851 11781
rect 35894 11772 35900 11784
rect 35952 11772 35958 11824
rect 36630 11772 36636 11824
rect 36688 11812 36694 11824
rect 37090 11812 37096 11824
rect 36688 11784 37096 11812
rect 36688 11772 36694 11784
rect 37090 11772 37096 11784
rect 37148 11812 37154 11824
rect 37369 11815 37427 11821
rect 37369 11812 37381 11815
rect 37148 11784 37381 11812
rect 37148 11772 37154 11784
rect 37369 11781 37381 11784
rect 37415 11781 37427 11815
rect 37550 11812 37556 11824
rect 37511 11784 37556 11812
rect 37369 11775 37427 11781
rect 37550 11772 37556 11784
rect 37608 11772 37614 11824
rect 38013 11815 38071 11821
rect 38013 11781 38025 11815
rect 38059 11812 38071 11815
rect 38102 11812 38108 11824
rect 38059 11784 38108 11812
rect 38059 11781 38071 11784
rect 38013 11775 38071 11781
rect 38102 11772 38108 11784
rect 38160 11772 38166 11824
rect 17212 11747 17270 11753
rect 17212 11713 17224 11747
rect 17258 11744 17270 11747
rect 17494 11744 17500 11756
rect 17258 11716 17500 11744
rect 17258 11713 17270 11716
rect 17212 11707 17270 11713
rect 17494 11704 17500 11716
rect 17552 11704 17558 11756
rect 20625 11747 20683 11753
rect 20625 11713 20637 11747
rect 20671 11744 20683 11747
rect 20806 11744 20812 11756
rect 20671 11716 20812 11744
rect 20671 11713 20683 11716
rect 20625 11707 20683 11713
rect 20806 11704 20812 11716
rect 20864 11704 20870 11756
rect 23750 11744 23756 11756
rect 23711 11716 23756 11744
rect 23750 11704 23756 11716
rect 23808 11704 23814 11756
rect 24394 11744 24400 11756
rect 24355 11716 24400 11744
rect 24394 11704 24400 11716
rect 24452 11704 24458 11756
rect 25038 11744 25044 11756
rect 24999 11716 25044 11744
rect 25038 11704 25044 11716
rect 25096 11704 25102 11756
rect 25866 11744 25872 11756
rect 25827 11716 25872 11744
rect 25866 11704 25872 11716
rect 25924 11704 25930 11756
rect 28442 11744 28448 11756
rect 28403 11716 28448 11744
rect 28442 11704 28448 11716
rect 28500 11704 28506 11756
rect 31018 11704 31024 11756
rect 31076 11744 31082 11756
rect 33502 11744 33508 11756
rect 31076 11716 31432 11744
rect 33463 11716 33508 11744
rect 31076 11704 31082 11716
rect 16666 11636 16672 11688
rect 16724 11676 16730 11688
rect 16945 11679 17003 11685
rect 16945 11676 16957 11679
rect 16724 11648 16957 11676
rect 16724 11636 16730 11648
rect 16945 11645 16957 11648
rect 16991 11645 17003 11679
rect 16945 11639 17003 11645
rect 18785 11679 18843 11685
rect 18785 11645 18797 11679
rect 18831 11645 18843 11679
rect 19058 11676 19064 11688
rect 19019 11648 19064 11676
rect 18785 11639 18843 11645
rect 16960 11540 16988 11639
rect 18325 11611 18383 11617
rect 18325 11577 18337 11611
rect 18371 11608 18383 11611
rect 18506 11608 18512 11620
rect 18371 11580 18512 11608
rect 18371 11577 18383 11580
rect 18325 11571 18383 11577
rect 18506 11568 18512 11580
rect 18564 11608 18570 11620
rect 18800 11608 18828 11639
rect 19058 11636 19064 11648
rect 19116 11636 19122 11688
rect 31294 11676 31300 11688
rect 31255 11648 31300 11676
rect 31294 11636 31300 11648
rect 31352 11636 31358 11688
rect 31404 11685 31432 11716
rect 33502 11704 33508 11716
rect 33560 11704 33566 11756
rect 34698 11744 34704 11756
rect 34659 11716 34704 11744
rect 34698 11704 34704 11716
rect 34756 11704 34762 11756
rect 35710 11747 35768 11753
rect 35710 11713 35722 11747
rect 35756 11744 35768 11747
rect 37182 11744 37188 11756
rect 35756 11716 37188 11744
rect 35756 11713 35768 11716
rect 35710 11707 35768 11713
rect 37182 11704 37188 11716
rect 37240 11704 37246 11756
rect 37279 11747 37337 11753
rect 37279 11713 37291 11747
rect 37325 11744 37337 11747
rect 38194 11744 38200 11756
rect 37325 11716 38200 11744
rect 37325 11713 37337 11716
rect 37279 11707 37337 11713
rect 37384 11688 37412 11716
rect 38194 11704 38200 11716
rect 38252 11704 38258 11756
rect 38286 11704 38292 11756
rect 38344 11744 38350 11756
rect 38344 11716 38389 11744
rect 38344 11704 38350 11716
rect 42886 11704 42892 11756
rect 42944 11744 42950 11756
rect 43349 11747 43407 11753
rect 43349 11744 43361 11747
rect 42944 11716 43361 11744
rect 42944 11704 42950 11716
rect 43349 11713 43361 11716
rect 43395 11713 43407 11747
rect 44174 11744 44180 11756
rect 44135 11716 44180 11744
rect 43349 11707 43407 11713
rect 44174 11704 44180 11716
rect 44232 11704 44238 11756
rect 31389 11679 31447 11685
rect 31389 11645 31401 11679
rect 31435 11645 31447 11679
rect 31389 11639 31447 11645
rect 34977 11679 35035 11685
rect 34977 11645 34989 11679
rect 35023 11645 35035 11679
rect 36170 11676 36176 11688
rect 36131 11648 36176 11676
rect 34977 11639 35035 11645
rect 18564 11580 18828 11608
rect 34992 11608 35020 11639
rect 36170 11636 36176 11648
rect 36228 11636 36234 11688
rect 37366 11636 37372 11688
rect 37424 11636 37430 11688
rect 35710 11608 35716 11620
rect 34992 11580 35716 11608
rect 18564 11568 18570 11580
rect 35710 11568 35716 11580
rect 35768 11568 35774 11620
rect 36262 11568 36268 11620
rect 36320 11608 36326 11620
rect 38013 11611 38071 11617
rect 38013 11608 38025 11611
rect 36320 11580 38025 11608
rect 36320 11568 36326 11580
rect 38013 11577 38025 11580
rect 38059 11577 38071 11611
rect 38013 11571 38071 11577
rect 17678 11540 17684 11552
rect 16960 11512 17684 11540
rect 17678 11500 17684 11512
rect 17736 11500 17742 11552
rect 19610 11500 19616 11552
rect 19668 11540 19674 11552
rect 20073 11543 20131 11549
rect 20073 11540 20085 11543
rect 19668 11512 20085 11540
rect 19668 11500 19674 11512
rect 20073 11509 20085 11512
rect 20119 11509 20131 11543
rect 20073 11503 20131 11509
rect 20257 11543 20315 11549
rect 20257 11509 20269 11543
rect 20303 11540 20315 11543
rect 20714 11540 20720 11552
rect 20303 11512 20720 11540
rect 20303 11509 20315 11512
rect 20257 11503 20315 11509
rect 20714 11500 20720 11512
rect 20772 11500 20778 11552
rect 23937 11543 23995 11549
rect 23937 11509 23949 11543
rect 23983 11540 23995 11543
rect 24210 11540 24216 11552
rect 23983 11512 24216 11540
rect 23983 11509 23995 11512
rect 23937 11503 23995 11509
rect 24210 11500 24216 11512
rect 24268 11500 24274 11552
rect 25225 11543 25283 11549
rect 25225 11509 25237 11543
rect 25271 11540 25283 11543
rect 25406 11540 25412 11552
rect 25271 11512 25412 11540
rect 25271 11509 25283 11512
rect 25225 11503 25283 11509
rect 25406 11500 25412 11512
rect 25464 11500 25470 11552
rect 36081 11543 36139 11549
rect 36081 11509 36093 11543
rect 36127 11540 36139 11543
rect 37826 11540 37832 11552
rect 36127 11512 37832 11540
rect 36127 11509 36139 11512
rect 36081 11503 36139 11509
rect 37826 11500 37832 11512
rect 37884 11500 37890 11552
rect 1104 11450 44896 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 44896 11450
rect 1104 11376 44896 11398
rect 18506 11336 18512 11348
rect 18467 11308 18512 11336
rect 18506 11296 18512 11308
rect 18564 11296 18570 11348
rect 18690 11336 18696 11348
rect 18651 11308 18696 11336
rect 18690 11296 18696 11308
rect 18748 11296 18754 11348
rect 21634 11336 21640 11348
rect 21595 11308 21640 11336
rect 21634 11296 21640 11308
rect 21692 11296 21698 11348
rect 23661 11339 23719 11345
rect 23661 11305 23673 11339
rect 23707 11336 23719 11339
rect 24394 11336 24400 11348
rect 23707 11308 24400 11336
rect 23707 11305 23719 11308
rect 23661 11299 23719 11305
rect 24394 11296 24400 11308
rect 24452 11296 24458 11348
rect 24765 11339 24823 11345
rect 24765 11305 24777 11339
rect 24811 11336 24823 11339
rect 25038 11336 25044 11348
rect 24811 11308 25044 11336
rect 24811 11305 24823 11308
rect 24765 11299 24823 11305
rect 25038 11296 25044 11308
rect 25096 11296 25102 11348
rect 26786 11296 26792 11348
rect 26844 11336 26850 11348
rect 27157 11339 27215 11345
rect 27157 11336 27169 11339
rect 26844 11308 27169 11336
rect 26844 11296 26850 11308
rect 27157 11305 27169 11308
rect 27203 11305 27215 11339
rect 27338 11336 27344 11348
rect 27299 11308 27344 11336
rect 27157 11299 27215 11305
rect 27338 11296 27344 11308
rect 27396 11296 27402 11348
rect 31294 11296 31300 11348
rect 31352 11336 31358 11348
rect 31849 11339 31907 11345
rect 31849 11336 31861 11339
rect 31352 11308 31861 11336
rect 31352 11296 31358 11308
rect 31849 11305 31861 11308
rect 31895 11305 31907 11339
rect 31849 11299 31907 11305
rect 34698 11296 34704 11348
rect 34756 11336 34762 11348
rect 35253 11339 35311 11345
rect 35253 11336 35265 11339
rect 34756 11308 35265 11336
rect 34756 11296 34762 11308
rect 35253 11305 35265 11308
rect 35299 11305 35311 11339
rect 35253 11299 35311 11305
rect 18230 11268 18236 11280
rect 17604 11240 18236 11268
rect 17126 11160 17132 11212
rect 17184 11200 17190 11212
rect 17604 11209 17632 11240
rect 18230 11228 18236 11240
rect 18288 11268 18294 11280
rect 19426 11268 19432 11280
rect 18288 11240 19432 11268
rect 18288 11228 18294 11240
rect 19426 11228 19432 11240
rect 19484 11228 19490 11280
rect 26697 11271 26755 11277
rect 26697 11237 26709 11271
rect 26743 11237 26755 11271
rect 26697 11231 26755 11237
rect 32033 11271 32091 11277
rect 32033 11237 32045 11271
rect 32079 11268 32091 11271
rect 32769 11271 32827 11277
rect 32769 11268 32781 11271
rect 32079 11240 32781 11268
rect 32079 11237 32091 11240
rect 32033 11231 32091 11237
rect 32769 11237 32781 11240
rect 32815 11237 32827 11271
rect 32769 11231 32827 11237
rect 17589 11203 17647 11209
rect 17589 11200 17601 11203
rect 17184 11172 17601 11200
rect 17184 11160 17190 11172
rect 17589 11169 17601 11172
rect 17635 11169 17647 11203
rect 17589 11163 17647 11169
rect 17678 11160 17684 11212
rect 17736 11200 17742 11212
rect 19334 11200 19340 11212
rect 17736 11172 19340 11200
rect 17736 11160 17742 11172
rect 19334 11160 19340 11172
rect 19392 11200 19398 11212
rect 20257 11203 20315 11209
rect 20257 11200 20269 11203
rect 19392 11172 20269 11200
rect 19392 11160 19398 11172
rect 20257 11169 20269 11172
rect 20303 11169 20315 11203
rect 20257 11163 20315 11169
rect 23293 11203 23351 11209
rect 23293 11169 23305 11203
rect 23339 11200 23351 11203
rect 23339 11172 24256 11200
rect 23339 11169 23351 11172
rect 23293 11163 23351 11169
rect 24228 11144 24256 11172
rect 2041 11135 2099 11141
rect 2041 11101 2053 11135
rect 2087 11132 2099 11135
rect 3234 11132 3240 11144
rect 2087 11104 3240 11132
rect 2087 11101 2099 11104
rect 2041 11095 2099 11101
rect 3234 11092 3240 11104
rect 3292 11092 3298 11144
rect 17770 11132 17776 11144
rect 17731 11104 17776 11132
rect 17770 11092 17776 11104
rect 17828 11092 17834 11144
rect 17862 11092 17868 11144
rect 17920 11132 17926 11144
rect 19058 11132 19064 11144
rect 17920 11104 19064 11132
rect 17920 11092 17926 11104
rect 19058 11092 19064 11104
rect 19116 11092 19122 11144
rect 19610 11132 19616 11144
rect 19571 11104 19616 11132
rect 19610 11092 19616 11104
rect 19668 11092 19674 11144
rect 23474 11132 23480 11144
rect 23435 11104 23480 11132
rect 23474 11092 23480 11104
rect 23532 11092 23538 11144
rect 24210 11092 24216 11144
rect 24268 11132 24274 11144
rect 24397 11135 24455 11141
rect 24397 11132 24409 11135
rect 24268 11104 24409 11132
rect 24268 11092 24274 11104
rect 24397 11101 24409 11104
rect 24443 11101 24455 11135
rect 24397 11095 24455 11101
rect 24581 11135 24639 11141
rect 24581 11101 24593 11135
rect 24627 11101 24639 11135
rect 24581 11095 24639 11101
rect 18322 11064 18328 11076
rect 18283 11036 18328 11064
rect 18322 11024 18328 11036
rect 18380 11024 18386 11076
rect 20502 11067 20560 11073
rect 20502 11064 20514 11067
rect 19812 11036 20514 11064
rect 17586 10996 17592 11008
rect 17547 10968 17592 10996
rect 17586 10956 17592 10968
rect 17644 10956 17650 11008
rect 17770 10956 17776 11008
rect 17828 10996 17834 11008
rect 19812 11005 19840 11036
rect 20502 11033 20514 11036
rect 20548 11033 20560 11067
rect 20502 11027 20560 11033
rect 20806 11024 20812 11076
rect 20864 11064 20870 11076
rect 24596 11064 24624 11095
rect 24762 11092 24768 11144
rect 24820 11132 24826 11144
rect 25317 11135 25375 11141
rect 25317 11132 25329 11135
rect 24820 11104 25329 11132
rect 24820 11092 24826 11104
rect 25317 11101 25329 11104
rect 25363 11101 25375 11135
rect 25317 11095 25375 11101
rect 25406 11092 25412 11144
rect 25464 11132 25470 11144
rect 25573 11135 25631 11141
rect 25573 11132 25585 11135
rect 25464 11104 25585 11132
rect 25464 11092 25470 11104
rect 25573 11101 25585 11104
rect 25619 11101 25631 11135
rect 26712 11132 26740 11231
rect 27525 11203 27583 11209
rect 27525 11169 27537 11203
rect 27571 11200 27583 11203
rect 27982 11200 27988 11212
rect 27571 11172 27988 11200
rect 27571 11169 27583 11172
rect 27525 11163 27583 11169
rect 27982 11160 27988 11172
rect 28040 11160 28046 11212
rect 36170 11200 36176 11212
rect 35728 11172 36176 11200
rect 27341 11135 27399 11141
rect 27341 11132 27353 11135
rect 26712 11104 27353 11132
rect 25573 11095 25631 11101
rect 27341 11101 27353 11104
rect 27387 11101 27399 11135
rect 28261 11135 28319 11141
rect 28261 11132 28273 11135
rect 27341 11095 27399 11101
rect 27632 11104 28273 11132
rect 27632 11076 27660 11104
rect 28261 11101 28273 11104
rect 28307 11101 28319 11135
rect 30190 11132 30196 11144
rect 30151 11104 30196 11132
rect 28261 11095 28319 11101
rect 30190 11092 30196 11104
rect 30248 11092 30254 11144
rect 33502 11092 33508 11144
rect 33560 11132 33566 11144
rect 34149 11135 34207 11141
rect 34149 11132 34161 11135
rect 33560 11104 34161 11132
rect 33560 11092 33566 11104
rect 34149 11101 34161 11104
rect 34195 11101 34207 11135
rect 34149 11095 34207 11101
rect 35342 11092 35348 11144
rect 35400 11132 35406 11144
rect 35728 11141 35756 11172
rect 36170 11160 36176 11172
rect 36228 11200 36234 11212
rect 36357 11203 36415 11209
rect 36357 11200 36369 11203
rect 36228 11172 36369 11200
rect 36228 11160 36234 11172
rect 36357 11169 36369 11172
rect 36403 11169 36415 11203
rect 43714 11200 43720 11212
rect 43675 11172 43720 11200
rect 36357 11163 36415 11169
rect 43714 11160 43720 11172
rect 43772 11160 43778 11212
rect 35437 11135 35495 11141
rect 35437 11132 35449 11135
rect 35400 11104 35449 11132
rect 35400 11092 35406 11104
rect 35437 11101 35449 11104
rect 35483 11101 35495 11135
rect 35437 11095 35495 11101
rect 35713 11135 35771 11141
rect 35713 11101 35725 11135
rect 35759 11101 35771 11135
rect 35713 11095 35771 11101
rect 35897 11135 35955 11141
rect 35897 11101 35909 11135
rect 35943 11132 35955 11135
rect 37366 11132 37372 11144
rect 35943 11104 37372 11132
rect 35943 11101 35955 11104
rect 35897 11095 35955 11101
rect 37366 11092 37372 11104
rect 37424 11092 37430 11144
rect 44174 11092 44180 11144
rect 44232 11132 44238 11144
rect 44232 11104 44277 11132
rect 44232 11092 44238 11104
rect 27614 11064 27620 11076
rect 20864 11036 24624 11064
rect 27575 11036 27620 11064
rect 20864 11024 20870 11036
rect 27614 11024 27620 11036
rect 27672 11024 27678 11076
rect 27798 11024 27804 11076
rect 27856 11064 27862 11076
rect 28077 11067 28135 11073
rect 28077 11064 28089 11067
rect 27856 11036 28089 11064
rect 27856 11024 27862 11036
rect 28077 11033 28089 11036
rect 28123 11033 28135 11067
rect 32306 11064 32312 11076
rect 32267 11036 32312 11064
rect 28077 11027 28135 11033
rect 32306 11024 32312 11036
rect 32364 11024 32370 11076
rect 33778 11024 33784 11076
rect 33836 11064 33842 11076
rect 33882 11067 33940 11073
rect 33882 11064 33894 11067
rect 33836 11036 33894 11064
rect 33836 11024 33842 11036
rect 33882 11033 33894 11036
rect 33928 11033 33940 11067
rect 33882 11027 33940 11033
rect 36541 11067 36599 11073
rect 36541 11033 36553 11067
rect 36587 11064 36599 11067
rect 36630 11064 36636 11076
rect 36587 11036 36636 11064
rect 36587 11033 36599 11036
rect 36541 11027 36599 11033
rect 36630 11024 36636 11036
rect 36688 11024 36694 11076
rect 36725 11067 36783 11073
rect 36725 11033 36737 11067
rect 36771 11064 36783 11067
rect 37642 11064 37648 11076
rect 36771 11036 37648 11064
rect 36771 11033 36783 11036
rect 36725 11027 36783 11033
rect 37642 11024 37648 11036
rect 37700 11024 37706 11076
rect 43990 11064 43996 11076
rect 43951 11036 43996 11064
rect 43990 11024 43996 11036
rect 44048 11024 44054 11076
rect 18525 10999 18583 11005
rect 18525 10996 18537 10999
rect 17828 10968 18537 10996
rect 17828 10956 17834 10968
rect 18525 10965 18537 10968
rect 18571 10965 18583 10999
rect 18525 10959 18583 10965
rect 19797 10999 19855 11005
rect 19797 10965 19809 10999
rect 19843 10965 19855 10999
rect 19797 10959 19855 10965
rect 28166 10956 28172 11008
rect 28224 10996 28230 11008
rect 28445 10999 28503 11005
rect 28445 10996 28457 10999
rect 28224 10968 28457 10996
rect 28224 10956 28230 10968
rect 28445 10965 28457 10968
rect 28491 10965 28503 10999
rect 30834 10996 30840 11008
rect 30795 10968 30840 10996
rect 28445 10959 28503 10965
rect 30834 10956 30840 10968
rect 30892 10956 30898 11008
rect 1104 10906 44896 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 44896 10906
rect 1104 10832 44896 10854
rect 17681 10795 17739 10801
rect 17681 10761 17693 10795
rect 17727 10792 17739 10795
rect 17862 10792 17868 10804
rect 17727 10764 17868 10792
rect 17727 10761 17739 10764
rect 17681 10755 17739 10761
rect 17862 10752 17868 10764
rect 17920 10752 17926 10804
rect 20254 10752 20260 10804
rect 20312 10792 20318 10804
rect 20441 10795 20499 10801
rect 20441 10792 20453 10795
rect 20312 10764 20453 10792
rect 20312 10752 20318 10764
rect 20441 10761 20453 10764
rect 20487 10761 20499 10795
rect 23658 10792 23664 10804
rect 23619 10764 23664 10792
rect 20441 10755 20499 10761
rect 23658 10752 23664 10764
rect 23716 10752 23722 10804
rect 26421 10795 26479 10801
rect 26421 10761 26433 10795
rect 26467 10792 26479 10795
rect 27338 10792 27344 10804
rect 26467 10764 27344 10792
rect 26467 10761 26479 10764
rect 26421 10755 26479 10761
rect 27338 10752 27344 10764
rect 27396 10752 27402 10804
rect 28353 10795 28411 10801
rect 28353 10761 28365 10795
rect 28399 10761 28411 10795
rect 30190 10792 30196 10804
rect 30151 10764 30196 10792
rect 28353 10755 28411 10761
rect 17497 10727 17555 10733
rect 17497 10693 17509 10727
rect 17543 10724 17555 10727
rect 17586 10724 17592 10736
rect 17543 10696 17592 10724
rect 17543 10693 17555 10696
rect 17497 10687 17555 10693
rect 17586 10684 17592 10696
rect 17644 10684 17650 10736
rect 19058 10684 19064 10736
rect 19116 10724 19122 10736
rect 28368 10724 28396 10755
rect 30190 10752 30196 10764
rect 30248 10752 30254 10804
rect 43441 10795 43499 10801
rect 43441 10761 43453 10795
rect 43487 10792 43499 10795
rect 43990 10792 43996 10804
rect 43487 10764 43996 10792
rect 43487 10761 43499 10764
rect 43441 10755 43499 10761
rect 43990 10752 43996 10764
rect 44048 10752 44054 10804
rect 29058 10727 29116 10733
rect 29058 10724 29070 10727
rect 19116 10696 24348 10724
rect 28368 10696 29070 10724
rect 19116 10684 19122 10696
rect 2590 10656 2596 10668
rect 2503 10628 2596 10656
rect 2590 10616 2596 10628
rect 2648 10656 2654 10668
rect 4982 10656 4988 10668
rect 2648 10628 4988 10656
rect 2648 10616 2654 10628
rect 4982 10616 4988 10628
rect 5040 10616 5046 10668
rect 17770 10616 17776 10668
rect 17828 10656 17834 10668
rect 18325 10659 18383 10665
rect 18325 10656 18337 10659
rect 17828 10628 18337 10656
rect 17828 10616 17834 10628
rect 18325 10625 18337 10628
rect 18371 10625 18383 10659
rect 18325 10619 18383 10625
rect 18414 10616 18420 10668
rect 18472 10656 18478 10668
rect 20732 10665 20760 10696
rect 18509 10659 18567 10665
rect 18509 10656 18521 10659
rect 18472 10628 18521 10656
rect 18472 10616 18478 10628
rect 18509 10625 18521 10628
rect 18555 10656 18567 10659
rect 20625 10659 20683 10665
rect 20625 10656 20637 10659
rect 18555 10628 20637 10656
rect 18555 10625 18567 10628
rect 18509 10619 18567 10625
rect 20625 10625 20637 10628
rect 20671 10625 20683 10659
rect 20625 10619 20683 10625
rect 20717 10659 20775 10665
rect 20717 10625 20729 10659
rect 20763 10625 20775 10659
rect 20717 10619 20775 10625
rect 18690 10588 18696 10600
rect 18603 10560 18696 10588
rect 18690 10548 18696 10560
rect 18748 10588 18754 10600
rect 18748 10560 19012 10588
rect 18748 10548 18754 10560
rect 17494 10520 17500 10532
rect 17455 10492 17500 10520
rect 17494 10480 17500 10492
rect 17552 10480 17558 10532
rect 1854 10412 1860 10464
rect 1912 10452 1918 10464
rect 1949 10455 2007 10461
rect 1949 10452 1961 10455
rect 1912 10424 1961 10452
rect 1912 10412 1918 10424
rect 1949 10421 1961 10424
rect 1995 10421 2007 10455
rect 1949 10415 2007 10421
rect 2130 10412 2136 10464
rect 2188 10452 2194 10464
rect 2501 10455 2559 10461
rect 2501 10452 2513 10455
rect 2188 10424 2513 10452
rect 2188 10412 2194 10424
rect 2501 10421 2513 10424
rect 2547 10421 2559 10455
rect 18984 10452 19012 10560
rect 20640 10520 20668 10619
rect 23106 10616 23112 10668
rect 23164 10656 23170 10668
rect 23477 10659 23535 10665
rect 23477 10656 23489 10659
rect 23164 10628 23489 10656
rect 23164 10616 23170 10628
rect 23477 10625 23489 10628
rect 23523 10625 23535 10659
rect 24210 10656 24216 10668
rect 24171 10628 24216 10656
rect 23477 10619 23535 10625
rect 24210 10616 24216 10628
rect 24268 10616 24274 10668
rect 24320 10665 24348 10696
rect 29058 10693 29070 10696
rect 29104 10693 29116 10727
rect 29058 10687 29116 10693
rect 24305 10659 24363 10665
rect 24305 10625 24317 10659
rect 24351 10625 24363 10659
rect 24305 10619 24363 10625
rect 24946 10616 24952 10668
rect 25004 10656 25010 10668
rect 25297 10659 25355 10665
rect 25297 10656 25309 10659
rect 25004 10628 25309 10656
rect 25004 10616 25010 10628
rect 25297 10625 25309 10628
rect 25343 10625 25355 10659
rect 28166 10656 28172 10668
rect 28127 10628 28172 10656
rect 25297 10619 25355 10625
rect 28166 10616 28172 10628
rect 28224 10616 28230 10668
rect 28442 10616 28448 10668
rect 28500 10656 28506 10668
rect 28813 10659 28871 10665
rect 28813 10656 28825 10659
rect 28500 10628 28825 10656
rect 28500 10616 28506 10628
rect 28813 10625 28825 10628
rect 28859 10625 28871 10659
rect 43346 10656 43352 10668
rect 43307 10628 43352 10656
rect 28813 10619 28871 10625
rect 43346 10616 43352 10628
rect 43404 10616 43410 10668
rect 44174 10656 44180 10668
rect 44135 10628 44180 10656
rect 44174 10616 44180 10628
rect 44232 10616 44238 10668
rect 20806 10588 20812 10600
rect 20767 10560 20812 10588
rect 20806 10548 20812 10560
rect 20864 10548 20870 10600
rect 20901 10591 20959 10597
rect 20901 10557 20913 10591
rect 20947 10588 20959 10591
rect 21634 10588 21640 10600
rect 20947 10560 21640 10588
rect 20947 10557 20959 10560
rect 20901 10551 20959 10557
rect 21634 10548 21640 10560
rect 21692 10548 21698 10600
rect 23293 10591 23351 10597
rect 23293 10557 23305 10591
rect 23339 10588 23351 10591
rect 24228 10588 24256 10616
rect 23339 10560 24256 10588
rect 23339 10557 23351 10560
rect 23293 10551 23351 10557
rect 24854 10548 24860 10600
rect 24912 10588 24918 10600
rect 25041 10591 25099 10597
rect 25041 10588 25053 10591
rect 24912 10560 25053 10588
rect 24912 10548 24918 10560
rect 25041 10557 25053 10560
rect 25087 10557 25099 10591
rect 25041 10551 25099 10557
rect 21910 10520 21916 10532
rect 20640 10492 21916 10520
rect 21910 10480 21916 10492
rect 21968 10480 21974 10532
rect 20806 10452 20812 10464
rect 18984 10424 20812 10452
rect 2501 10415 2559 10421
rect 20806 10412 20812 10424
rect 20864 10412 20870 10464
rect 24489 10455 24547 10461
rect 24489 10421 24501 10455
rect 24535 10452 24547 10455
rect 25406 10452 25412 10464
rect 24535 10424 25412 10452
rect 24535 10421 24547 10424
rect 24489 10415 24547 10421
rect 25406 10412 25412 10424
rect 25464 10412 25470 10464
rect 1104 10362 44896 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 44896 10362
rect 1104 10288 44896 10310
rect 17678 10248 17684 10260
rect 17328 10220 17684 10248
rect 1394 10112 1400 10124
rect 1355 10084 1400 10112
rect 1394 10072 1400 10084
rect 1452 10072 1458 10124
rect 3234 10112 3240 10124
rect 3195 10084 3240 10112
rect 3234 10072 3240 10084
rect 3292 10072 3298 10124
rect 17328 10121 17356 10220
rect 17678 10208 17684 10220
rect 17736 10208 17742 10260
rect 18690 10248 18696 10260
rect 18651 10220 18696 10248
rect 18690 10208 18696 10220
rect 18748 10208 18754 10260
rect 20714 10208 20720 10260
rect 20772 10248 20778 10260
rect 22281 10251 22339 10257
rect 22281 10248 22293 10251
rect 20772 10220 22293 10248
rect 20772 10208 20778 10220
rect 20824 10189 20852 10220
rect 22281 10217 22293 10220
rect 22327 10217 22339 10251
rect 22925 10251 22983 10257
rect 22925 10248 22937 10251
rect 22281 10211 22339 10217
rect 22388 10220 22937 10248
rect 20809 10183 20867 10189
rect 20809 10149 20821 10183
rect 20855 10149 20867 10183
rect 21910 10180 21916 10192
rect 21871 10152 21916 10180
rect 20809 10143 20867 10149
rect 21910 10140 21916 10152
rect 21968 10180 21974 10192
rect 22388 10180 22416 10220
rect 22925 10217 22937 10220
rect 22971 10217 22983 10251
rect 23106 10248 23112 10260
rect 23067 10220 23112 10248
rect 22925 10211 22983 10217
rect 23106 10208 23112 10220
rect 23164 10208 23170 10260
rect 31665 10251 31723 10257
rect 31665 10217 31677 10251
rect 31711 10248 31723 10251
rect 32306 10248 32312 10260
rect 31711 10220 32312 10248
rect 31711 10217 31723 10220
rect 31665 10211 31723 10217
rect 32306 10208 32312 10220
rect 32364 10208 32370 10260
rect 21968 10152 22416 10180
rect 22465 10183 22523 10189
rect 21968 10140 21974 10152
rect 22465 10149 22477 10183
rect 22511 10180 22523 10183
rect 23658 10180 23664 10192
rect 22511 10152 23664 10180
rect 22511 10149 22523 10152
rect 22465 10143 22523 10149
rect 23658 10140 23664 10152
rect 23716 10140 23722 10192
rect 17313 10115 17371 10121
rect 17313 10081 17325 10115
rect 17359 10081 17371 10115
rect 17313 10075 17371 10081
rect 19426 10072 19432 10124
rect 19484 10112 19490 10124
rect 19613 10115 19671 10121
rect 19613 10112 19625 10115
rect 19484 10084 19625 10112
rect 19484 10072 19490 10084
rect 19613 10081 19625 10084
rect 19659 10081 19671 10115
rect 19613 10075 19671 10081
rect 24210 10072 24216 10124
rect 24268 10112 24274 10124
rect 24397 10115 24455 10121
rect 24397 10112 24409 10115
rect 24268 10084 24409 10112
rect 24268 10072 24274 10084
rect 24397 10081 24409 10084
rect 24443 10081 24455 10115
rect 24397 10075 24455 10081
rect 28442 10072 28448 10124
rect 28500 10112 28506 10124
rect 30285 10115 30343 10121
rect 30285 10112 30297 10115
rect 28500 10084 30297 10112
rect 28500 10072 28506 10084
rect 30285 10081 30297 10084
rect 30331 10081 30343 10115
rect 30285 10075 30343 10081
rect 3970 10044 3976 10056
rect 3931 10016 3976 10044
rect 3970 10004 3976 10016
rect 4028 10004 4034 10056
rect 19797 10047 19855 10053
rect 19797 10013 19809 10047
rect 19843 10013 19855 10047
rect 19797 10007 19855 10013
rect 19889 10047 19947 10053
rect 19889 10013 19901 10047
rect 19935 10044 19947 10047
rect 20346 10044 20352 10056
rect 19935 10016 20352 10044
rect 19935 10013 19947 10016
rect 19889 10007 19947 10013
rect 3053 9979 3111 9985
rect 3053 9945 3065 9979
rect 3099 9976 3111 9979
rect 3881 9979 3939 9985
rect 3881 9976 3893 9979
rect 3099 9948 3893 9976
rect 3099 9945 3111 9948
rect 3053 9939 3111 9945
rect 3881 9945 3893 9948
rect 3927 9945 3939 9979
rect 3881 9939 3939 9945
rect 17580 9979 17638 9985
rect 17580 9945 17592 9979
rect 17626 9976 17638 9979
rect 17678 9976 17684 9988
rect 17626 9948 17684 9976
rect 17626 9945 17638 9948
rect 17580 9939 17638 9945
rect 17678 9936 17684 9948
rect 17736 9936 17742 9988
rect 19812 9976 19840 10007
rect 20346 10004 20352 10016
rect 20404 10004 20410 10056
rect 22922 10004 22928 10056
rect 22980 10044 22986 10056
rect 24581 10047 24639 10053
rect 24581 10044 24593 10047
rect 22980 10016 24593 10044
rect 22980 10004 22986 10016
rect 20530 9976 20536 9988
rect 19812 9948 20536 9976
rect 20530 9936 20536 9948
rect 20588 9936 20594 9988
rect 23308 9985 23336 10016
rect 24581 10013 24593 10016
rect 24627 10013 24639 10047
rect 24581 10007 24639 10013
rect 24854 10004 24860 10056
rect 24912 10044 24918 10056
rect 25225 10047 25283 10053
rect 25225 10044 25237 10047
rect 24912 10016 25237 10044
rect 24912 10004 24918 10016
rect 25225 10013 25237 10016
rect 25271 10044 25283 10047
rect 27433 10047 27491 10053
rect 27433 10044 27445 10047
rect 25271 10016 27445 10044
rect 25271 10013 25283 10016
rect 25225 10007 25283 10013
rect 27433 10013 27445 10016
rect 27479 10013 27491 10047
rect 27433 10007 27491 10013
rect 30552 10047 30610 10053
rect 30552 10013 30564 10047
rect 30598 10044 30610 10047
rect 30834 10044 30840 10056
rect 30598 10016 30840 10044
rect 30598 10013 30610 10016
rect 30552 10007 30610 10013
rect 30834 10004 30840 10016
rect 30892 10004 30898 10056
rect 23293 9979 23351 9985
rect 23293 9945 23305 9979
rect 23339 9945 23351 9979
rect 23293 9939 23351 9945
rect 25492 9979 25550 9985
rect 25492 9945 25504 9979
rect 25538 9976 25550 9979
rect 25590 9976 25596 9988
rect 25538 9948 25596 9976
rect 25538 9945 25550 9948
rect 25492 9939 25550 9945
rect 25590 9936 25596 9948
rect 25648 9936 25654 9988
rect 27614 9976 27620 9988
rect 26620 9948 27620 9976
rect 19426 9868 19432 9920
rect 19484 9908 19490 9920
rect 19613 9911 19671 9917
rect 19613 9908 19625 9911
rect 19484 9880 19625 9908
rect 19484 9868 19490 9880
rect 19613 9877 19625 9880
rect 19659 9877 19671 9911
rect 20990 9908 20996 9920
rect 20951 9880 20996 9908
rect 19613 9871 19671 9877
rect 20990 9868 20996 9880
rect 21048 9868 21054 9920
rect 22278 9908 22284 9920
rect 22239 9880 22284 9908
rect 22278 9868 22284 9880
rect 22336 9868 22342 9920
rect 23106 9917 23112 9920
rect 23093 9911 23112 9917
rect 23093 9877 23105 9911
rect 23093 9871 23112 9877
rect 23106 9868 23112 9871
rect 23164 9868 23170 9920
rect 24670 9868 24676 9920
rect 24728 9908 24734 9920
rect 26620 9917 26648 9948
rect 27614 9936 27620 9948
rect 27672 9985 27678 9988
rect 27672 9979 27736 9985
rect 27672 9945 27690 9979
rect 27724 9945 27736 9979
rect 27672 9939 27736 9945
rect 27672 9936 27678 9939
rect 24765 9911 24823 9917
rect 24765 9908 24777 9911
rect 24728 9880 24777 9908
rect 24728 9868 24734 9880
rect 24765 9877 24777 9880
rect 24811 9877 24823 9911
rect 24765 9871 24823 9877
rect 26605 9911 26663 9917
rect 26605 9877 26617 9911
rect 26651 9877 26663 9911
rect 26605 9871 26663 9877
rect 1104 9818 44896 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 44896 9818
rect 1104 9744 44896 9766
rect 17678 9704 17684 9716
rect 17639 9676 17684 9704
rect 17678 9664 17684 9676
rect 17736 9664 17742 9716
rect 24946 9704 24952 9716
rect 24907 9676 24952 9704
rect 24946 9664 24952 9676
rect 25004 9664 25010 9716
rect 25590 9704 25596 9716
rect 25551 9676 25596 9704
rect 25590 9664 25596 9676
rect 25648 9664 25654 9716
rect 3970 9596 3976 9648
rect 4028 9636 4034 9648
rect 4028 9608 26234 9636
rect 4028 9596 4034 9608
rect 17589 9571 17647 9577
rect 17589 9537 17601 9571
rect 17635 9537 17647 9571
rect 17770 9568 17776 9580
rect 17731 9540 17776 9568
rect 17589 9531 17647 9537
rect 1946 9500 1952 9512
rect 1907 9472 1952 9500
rect 1946 9460 1952 9472
rect 2004 9460 2010 9512
rect 2133 9503 2191 9509
rect 2133 9469 2145 9503
rect 2179 9500 2191 9503
rect 2498 9500 2504 9512
rect 2179 9472 2504 9500
rect 2179 9469 2191 9472
rect 2133 9463 2191 9469
rect 2498 9460 2504 9472
rect 2556 9460 2562 9512
rect 2774 9460 2780 9512
rect 2832 9500 2838 9512
rect 2832 9472 2877 9500
rect 2832 9460 2838 9472
rect 17604 9432 17632 9531
rect 17770 9528 17776 9540
rect 17828 9528 17834 9580
rect 18414 9568 18420 9580
rect 18375 9540 18420 9568
rect 18414 9528 18420 9540
rect 18472 9528 18478 9580
rect 18509 9571 18567 9577
rect 18509 9537 18521 9571
rect 18555 9568 18567 9571
rect 18690 9568 18696 9580
rect 18555 9540 18696 9568
rect 18555 9537 18567 9540
rect 18509 9531 18567 9537
rect 18690 9528 18696 9540
rect 18748 9528 18754 9580
rect 19334 9568 19340 9580
rect 19295 9540 19340 9568
rect 19334 9528 19340 9540
rect 19392 9528 19398 9580
rect 19610 9577 19616 9580
rect 19604 9568 19616 9577
rect 19571 9540 19616 9568
rect 19604 9531 19616 9540
rect 19610 9528 19616 9531
rect 19668 9528 19674 9580
rect 22370 9568 22376 9580
rect 22283 9540 22376 9568
rect 22370 9528 22376 9540
rect 22428 9568 22434 9580
rect 23106 9568 23112 9580
rect 22428 9540 23112 9568
rect 22428 9528 22434 9540
rect 23106 9528 23112 9540
rect 23164 9528 23170 9580
rect 23658 9568 23664 9580
rect 23619 9540 23664 9568
rect 23658 9528 23664 9540
rect 23716 9528 23722 9580
rect 24670 9528 24676 9580
rect 24728 9568 24734 9580
rect 24765 9571 24823 9577
rect 24765 9568 24777 9571
rect 24728 9540 24777 9568
rect 24728 9528 24734 9540
rect 24765 9537 24777 9540
rect 24811 9537 24823 9571
rect 25406 9568 25412 9580
rect 25367 9540 25412 9568
rect 24765 9531 24823 9537
rect 25406 9528 25412 9540
rect 25464 9528 25470 9580
rect 26206 9568 26234 9608
rect 42797 9571 42855 9577
rect 42797 9568 42809 9571
rect 26206 9540 42809 9568
rect 42797 9537 42809 9540
rect 42843 9537 42855 9571
rect 42797 9531 42855 9537
rect 18230 9500 18236 9512
rect 18191 9472 18236 9500
rect 18230 9460 18236 9472
rect 18288 9460 18294 9512
rect 20530 9460 20536 9512
rect 20588 9500 20594 9512
rect 22649 9503 22707 9509
rect 22649 9500 22661 9503
rect 20588 9472 22661 9500
rect 20588 9460 20594 9472
rect 22649 9469 22661 9472
rect 22695 9500 22707 9503
rect 23474 9500 23480 9512
rect 22695 9472 23480 9500
rect 22695 9469 22707 9472
rect 22649 9463 22707 9469
rect 23474 9460 23480 9472
rect 23532 9460 23538 9512
rect 18325 9435 18383 9441
rect 18325 9432 18337 9435
rect 17604 9404 18337 9432
rect 18325 9401 18337 9404
rect 18371 9401 18383 9435
rect 18325 9395 18383 9401
rect 20346 9392 20352 9444
rect 20404 9432 20410 9444
rect 20717 9435 20775 9441
rect 20717 9432 20729 9435
rect 20404 9404 20729 9432
rect 20404 9392 20410 9404
rect 20717 9401 20729 9404
rect 20763 9432 20775 9435
rect 23014 9432 23020 9444
rect 20763 9404 23020 9432
rect 20763 9401 20775 9404
rect 20717 9395 20775 9401
rect 23014 9392 23020 9404
rect 23072 9392 23078 9444
rect 23842 9364 23848 9376
rect 23803 9336 23848 9364
rect 23842 9324 23848 9336
rect 23900 9324 23906 9376
rect 42518 9324 42524 9376
rect 42576 9364 42582 9376
rect 42889 9367 42947 9373
rect 42889 9364 42901 9367
rect 42576 9336 42901 9364
rect 42576 9324 42582 9336
rect 42889 9333 42901 9336
rect 42935 9333 42947 9367
rect 42889 9327 42947 9333
rect 1104 9274 44896 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 44896 9274
rect 1104 9200 44896 9222
rect 1946 9160 1952 9172
rect 1907 9132 1952 9160
rect 1946 9120 1952 9132
rect 2004 9120 2010 9172
rect 2498 9160 2504 9172
rect 2459 9132 2504 9160
rect 2498 9120 2504 9132
rect 2556 9120 2562 9172
rect 19610 9160 19616 9172
rect 19571 9132 19616 9160
rect 19610 9120 19616 9132
rect 19668 9120 19674 9172
rect 22278 9120 22284 9172
rect 22336 9160 22342 9172
rect 22741 9163 22799 9169
rect 22741 9160 22753 9163
rect 22336 9132 22753 9160
rect 22336 9120 22342 9132
rect 22741 9129 22753 9132
rect 22787 9129 22799 9163
rect 22741 9123 22799 9129
rect 42518 9024 42524 9036
rect 42479 8996 42524 9024
rect 42518 8984 42524 8996
rect 42576 8984 42582 9036
rect 2590 8956 2596 8968
rect 2551 8928 2596 8956
rect 2590 8916 2596 8928
rect 2648 8916 2654 8968
rect 19426 8916 19432 8968
rect 19484 8956 19490 8968
rect 19613 8959 19671 8965
rect 19613 8956 19625 8959
rect 19484 8928 19625 8956
rect 19484 8916 19490 8928
rect 19613 8925 19625 8928
rect 19659 8925 19671 8959
rect 19613 8919 19671 8925
rect 19889 8959 19947 8965
rect 19889 8925 19901 8959
rect 19935 8956 19947 8959
rect 20530 8956 20536 8968
rect 19935 8928 20536 8956
rect 19935 8925 19947 8928
rect 19889 8919 19947 8925
rect 20530 8916 20536 8928
rect 20588 8916 20594 8968
rect 20901 8959 20959 8965
rect 20901 8925 20913 8959
rect 20947 8956 20959 8959
rect 22830 8956 22836 8968
rect 20947 8928 22836 8956
rect 20947 8925 20959 8928
rect 20901 8919 20959 8925
rect 22830 8916 22836 8928
rect 22888 8916 22894 8968
rect 22922 8916 22928 8968
rect 22980 8956 22986 8968
rect 23201 8959 23259 8965
rect 22980 8928 23025 8956
rect 22980 8916 22986 8928
rect 23201 8925 23213 8959
rect 23247 8956 23259 8959
rect 23474 8956 23480 8968
rect 23247 8928 23480 8956
rect 23247 8925 23259 8928
rect 23201 8919 23259 8925
rect 23474 8916 23480 8928
rect 23532 8916 23538 8968
rect 42334 8956 42340 8968
rect 42295 8928 42340 8956
rect 42334 8916 42340 8928
rect 42392 8916 42398 8968
rect 19797 8891 19855 8897
rect 19797 8857 19809 8891
rect 19843 8888 19855 8891
rect 20346 8888 20352 8900
rect 19843 8860 20352 8888
rect 19843 8857 19855 8860
rect 19797 8851 19855 8857
rect 20346 8848 20352 8860
rect 20404 8848 20410 8900
rect 21174 8897 21180 8900
rect 21168 8851 21180 8897
rect 21232 8888 21238 8900
rect 21232 8860 21268 8888
rect 21174 8848 21180 8851
rect 21232 8848 21238 8860
rect 23014 8848 23020 8900
rect 23072 8888 23078 8900
rect 23109 8891 23167 8897
rect 23109 8888 23121 8891
rect 23072 8860 23121 8888
rect 23072 8848 23078 8860
rect 23109 8857 23121 8860
rect 23155 8857 23167 8891
rect 23109 8851 23167 8857
rect 44177 8891 44235 8897
rect 44177 8857 44189 8891
rect 44223 8888 44235 8891
rect 45094 8888 45100 8900
rect 44223 8860 45100 8888
rect 44223 8857 44235 8860
rect 44177 8851 44235 8857
rect 45094 8848 45100 8860
rect 45152 8848 45158 8900
rect 22281 8823 22339 8829
rect 22281 8789 22293 8823
rect 22327 8820 22339 8823
rect 22370 8820 22376 8832
rect 22327 8792 22376 8820
rect 22327 8789 22339 8792
rect 22281 8783 22339 8789
rect 22370 8780 22376 8792
rect 22428 8780 22434 8832
rect 1104 8730 44896 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 44896 8730
rect 1104 8656 44896 8678
rect 21174 8616 21180 8628
rect 21135 8588 21180 8616
rect 21174 8576 21180 8588
rect 21232 8576 21238 8628
rect 22741 8619 22799 8625
rect 22741 8585 22753 8619
rect 22787 8616 22799 8619
rect 22922 8616 22928 8628
rect 22787 8588 22928 8616
rect 22787 8585 22799 8588
rect 22741 8579 22799 8585
rect 22922 8576 22928 8588
rect 22980 8576 22986 8628
rect 2130 8548 2136 8560
rect 2091 8520 2136 8548
rect 2130 8508 2136 8520
rect 2188 8508 2194 8560
rect 23842 8508 23848 8560
rect 23900 8557 23906 8560
rect 23900 8548 23912 8557
rect 23900 8520 23945 8548
rect 23900 8511 23912 8520
rect 23900 8508 23906 8511
rect 1854 8440 1860 8492
rect 1912 8480 1918 8492
rect 1949 8483 2007 8489
rect 1949 8480 1961 8483
rect 1912 8452 1961 8480
rect 1912 8440 1918 8452
rect 1949 8449 1961 8452
rect 1995 8449 2007 8483
rect 20990 8480 20996 8492
rect 20951 8452 20996 8480
rect 1949 8443 2007 8449
rect 20990 8440 20996 8452
rect 21048 8440 21054 8492
rect 24121 8483 24179 8489
rect 24121 8449 24133 8483
rect 24167 8480 24179 8483
rect 24762 8480 24768 8492
rect 24167 8452 24768 8480
rect 24167 8449 24179 8452
rect 24121 8443 24179 8449
rect 24762 8440 24768 8452
rect 24820 8440 24826 8492
rect 42334 8440 42340 8492
rect 42392 8480 42398 8492
rect 43625 8483 43683 8489
rect 43625 8480 43637 8483
rect 42392 8452 43637 8480
rect 42392 8440 42398 8452
rect 43625 8449 43637 8452
rect 43671 8449 43683 8483
rect 43625 8443 43683 8449
rect 2866 8412 2872 8424
rect 2827 8384 2872 8412
rect 2866 8372 2872 8384
rect 2924 8372 2930 8424
rect 1104 8186 44896 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 44896 8186
rect 1104 8112 44896 8134
rect 44174 7868 44180 7880
rect 44135 7840 44180 7868
rect 44174 7828 44180 7840
rect 44232 7828 44238 7880
rect 26326 7692 26332 7744
rect 26384 7732 26390 7744
rect 43993 7735 44051 7741
rect 43993 7732 44005 7735
rect 26384 7704 44005 7732
rect 26384 7692 26390 7704
rect 43993 7701 44005 7704
rect 44039 7701 44051 7735
rect 43993 7695 44051 7701
rect 1104 7642 44896 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 44896 7642
rect 1104 7568 44896 7590
rect 3418 7392 3424 7404
rect 3379 7364 3424 7392
rect 3418 7352 3424 7364
rect 3476 7352 3482 7404
rect 43533 7395 43591 7401
rect 43533 7361 43545 7395
rect 43579 7392 43591 7395
rect 43622 7392 43628 7404
rect 43579 7364 43628 7392
rect 43579 7361 43591 7364
rect 43533 7355 43591 7361
rect 43622 7352 43628 7364
rect 43680 7352 43686 7404
rect 3510 7188 3516 7200
rect 3471 7160 3516 7188
rect 3510 7148 3516 7160
rect 3568 7148 3574 7200
rect 4062 7188 4068 7200
rect 4023 7160 4068 7188
rect 4062 7148 4068 7160
rect 4120 7148 4126 7200
rect 43625 7191 43683 7197
rect 43625 7157 43637 7191
rect 43671 7188 43683 7191
rect 43990 7188 43996 7200
rect 43671 7160 43996 7188
rect 43671 7157 43683 7160
rect 43625 7151 43683 7157
rect 43990 7148 43996 7160
rect 44048 7148 44054 7200
rect 1104 7098 44896 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 44896 7098
rect 1104 7024 44896 7046
rect 3789 6851 3847 6857
rect 3789 6817 3801 6851
rect 3835 6848 3847 6851
rect 4062 6848 4068 6860
rect 3835 6820 4068 6848
rect 3835 6817 3847 6820
rect 3789 6811 3847 6817
rect 4062 6808 4068 6820
rect 4120 6808 4126 6860
rect 4706 6848 4712 6860
rect 4667 6820 4712 6848
rect 4706 6808 4712 6820
rect 4764 6808 4770 6860
rect 14734 6848 14740 6860
rect 5184 6820 14740 6848
rect 1670 6740 1676 6792
rect 1728 6780 1734 6792
rect 1765 6783 1823 6789
rect 1765 6780 1777 6783
rect 1728 6752 1777 6780
rect 1728 6740 1734 6752
rect 1765 6749 1777 6752
rect 1811 6749 1823 6783
rect 1765 6743 1823 6749
rect 3510 6672 3516 6724
rect 3568 6712 3574 6724
rect 3973 6715 4031 6721
rect 3973 6712 3985 6715
rect 3568 6684 3985 6712
rect 3568 6672 3574 6684
rect 3973 6681 3985 6684
rect 4019 6681 4031 6715
rect 3973 6675 4031 6681
rect 4062 6672 4068 6724
rect 4120 6712 4126 6724
rect 5184 6712 5212 6820
rect 14734 6808 14740 6820
rect 14792 6808 14798 6860
rect 42702 6848 42708 6860
rect 42663 6820 42708 6848
rect 42702 6808 42708 6820
rect 42760 6808 42766 6860
rect 43990 6848 43996 6860
rect 43951 6820 43996 6848
rect 43990 6808 43996 6820
rect 44048 6808 44054 6860
rect 44174 6740 44180 6792
rect 44232 6780 44238 6792
rect 44232 6752 44277 6780
rect 44232 6740 44238 6752
rect 4120 6684 5212 6712
rect 4120 6672 4126 6684
rect 1104 6554 44896 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 44896 6554
rect 1104 6480 44896 6502
rect 1670 6304 1676 6316
rect 1631 6276 1676 6304
rect 1670 6264 1676 6276
rect 1728 6264 1734 6316
rect 43809 6307 43867 6313
rect 43809 6273 43821 6307
rect 43855 6304 43867 6307
rect 44174 6304 44180 6316
rect 43855 6276 44180 6304
rect 43855 6273 43867 6276
rect 43809 6267 43867 6273
rect 44174 6264 44180 6276
rect 44232 6264 44238 6316
rect 1857 6239 1915 6245
rect 1857 6205 1869 6239
rect 1903 6236 1915 6239
rect 2130 6236 2136 6248
rect 1903 6208 2136 6236
rect 1903 6205 1915 6208
rect 1857 6199 1915 6205
rect 2130 6196 2136 6208
rect 2188 6196 2194 6248
rect 2774 6196 2780 6248
rect 2832 6236 2838 6248
rect 2832 6208 2877 6236
rect 2832 6196 2838 6208
rect 1104 6010 44896 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 44896 6010
rect 1104 5936 44896 5958
rect 2130 5896 2136 5908
rect 2091 5868 2136 5896
rect 2130 5856 2136 5868
rect 2188 5856 2194 5908
rect 5902 5828 5908 5840
rect 2240 5800 5908 5828
rect 1578 5692 1584 5704
rect 1539 5664 1584 5692
rect 1578 5652 1584 5664
rect 1636 5652 1642 5704
rect 2038 5652 2044 5704
rect 2096 5692 2102 5704
rect 2240 5701 2268 5800
rect 5902 5788 5908 5800
rect 5960 5788 5966 5840
rect 6270 5760 6276 5772
rect 2976 5732 6276 5760
rect 2976 5701 3004 5732
rect 6270 5720 6276 5732
rect 6328 5720 6334 5772
rect 42702 5760 42708 5772
rect 42663 5732 42708 5760
rect 42702 5720 42708 5732
rect 42760 5720 42766 5772
rect 2225 5695 2283 5701
rect 2225 5692 2237 5695
rect 2096 5664 2237 5692
rect 2096 5652 2102 5664
rect 2225 5661 2237 5664
rect 2271 5661 2283 5695
rect 2225 5655 2283 5661
rect 2961 5695 3019 5701
rect 2961 5661 2973 5695
rect 3007 5661 3019 5695
rect 3786 5692 3792 5704
rect 3747 5664 3792 5692
rect 2961 5655 3019 5661
rect 3786 5652 3792 5664
rect 3844 5652 3850 5704
rect 4154 5652 4160 5704
rect 4212 5692 4218 5704
rect 4433 5695 4491 5701
rect 4433 5692 4445 5695
rect 4212 5664 4445 5692
rect 4212 5652 4218 5664
rect 4433 5661 4445 5664
rect 4479 5661 4491 5695
rect 4433 5655 4491 5661
rect 44174 5652 44180 5704
rect 44232 5692 44238 5704
rect 44232 5664 44277 5692
rect 44232 5652 44238 5664
rect 43990 5624 43996 5636
rect 43951 5596 43996 5624
rect 43990 5584 43996 5596
rect 44048 5584 44054 5636
rect 2866 5556 2872 5568
rect 2827 5528 2872 5556
rect 2866 5516 2872 5528
rect 2924 5516 2930 5568
rect 1104 5466 44896 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 44896 5466
rect 1104 5392 44896 5414
rect 2133 5287 2191 5293
rect 2133 5253 2145 5287
rect 2179 5284 2191 5287
rect 2866 5284 2872 5296
rect 2179 5256 2872 5284
rect 2179 5253 2191 5256
rect 2133 5247 2191 5253
rect 2866 5244 2872 5256
rect 2924 5244 2930 5296
rect 1578 5176 1584 5228
rect 1636 5216 1642 5228
rect 1949 5219 2007 5225
rect 1949 5216 1961 5219
rect 1636 5188 1961 5216
rect 1636 5176 1642 5188
rect 1949 5185 1961 5188
rect 1995 5185 2007 5219
rect 1949 5179 2007 5185
rect 4433 5219 4491 5225
rect 4433 5185 4445 5219
rect 4479 5216 4491 5219
rect 4614 5216 4620 5228
rect 4479 5188 4620 5216
rect 4479 5185 4491 5188
rect 4433 5179 4491 5185
rect 4614 5176 4620 5188
rect 4672 5176 4678 5228
rect 42794 5216 42800 5228
rect 42755 5188 42800 5216
rect 42794 5176 42800 5188
rect 42852 5176 42858 5228
rect 2774 5108 2780 5160
rect 2832 5148 2838 5160
rect 2832 5120 2877 5148
rect 2832 5108 2838 5120
rect 4341 5015 4399 5021
rect 4341 4981 4353 5015
rect 4387 5012 4399 5015
rect 4614 5012 4620 5024
rect 4387 4984 4620 5012
rect 4387 4981 4399 4984
rect 4341 4975 4399 4981
rect 4614 4972 4620 4984
rect 4672 4972 4678 5024
rect 4890 5012 4896 5024
rect 4851 4984 4896 5012
rect 4890 4972 4896 4984
rect 4948 4972 4954 5024
rect 42518 4972 42524 5024
rect 42576 5012 42582 5024
rect 42889 5015 42947 5021
rect 42889 5012 42901 5015
rect 42576 4984 42901 5012
rect 42576 4972 42582 4984
rect 42889 4981 42901 4984
rect 42935 4981 42947 5015
rect 43622 5012 43628 5024
rect 43583 4984 43628 5012
rect 42889 4975 42947 4981
rect 43622 4972 43628 4984
rect 43680 4972 43686 5024
rect 1104 4922 44896 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 44896 4922
rect 1104 4848 44896 4870
rect 4798 4768 4804 4820
rect 4856 4768 4862 4820
rect 4816 4740 4844 4768
rect 11790 4740 11796 4752
rect 3252 4712 11796 4740
rect 1949 4675 2007 4681
rect 1949 4641 1961 4675
rect 1995 4672 2007 4675
rect 2958 4672 2964 4684
rect 1995 4644 2964 4672
rect 1995 4641 2007 4644
rect 1949 4635 2007 4641
rect 2958 4632 2964 4644
rect 3016 4632 3022 4684
rect 2593 4607 2651 4613
rect 2593 4573 2605 4607
rect 2639 4604 2651 4607
rect 3142 4604 3148 4616
rect 2639 4576 3148 4604
rect 2639 4573 2651 4576
rect 2593 4567 2651 4573
rect 3142 4564 3148 4576
rect 3200 4564 3206 4616
rect 3252 4613 3280 4712
rect 11790 4700 11796 4712
rect 11848 4700 11854 4752
rect 43622 4740 43628 4752
rect 42352 4712 43628 4740
rect 4062 4672 4068 4684
rect 4023 4644 4068 4672
rect 4062 4632 4068 4644
rect 4120 4632 4126 4684
rect 4249 4675 4307 4681
rect 4249 4641 4261 4675
rect 4295 4672 4307 4675
rect 4614 4672 4620 4684
rect 4295 4644 4620 4672
rect 4295 4641 4307 4644
rect 4249 4635 4307 4641
rect 4614 4632 4620 4644
rect 4672 4632 4678 4684
rect 4798 4672 4804 4684
rect 4759 4644 4804 4672
rect 4798 4632 4804 4644
rect 4856 4632 4862 4684
rect 38010 4672 38016 4684
rect 37971 4644 38016 4672
rect 38010 4632 38016 4644
rect 38068 4632 38074 4684
rect 42352 4681 42380 4712
rect 43622 4700 43628 4712
rect 43680 4700 43686 4752
rect 42337 4675 42395 4681
rect 42337 4641 42349 4675
rect 42383 4641 42395 4675
rect 42518 4672 42524 4684
rect 42479 4644 42524 4672
rect 42337 4635 42395 4641
rect 42518 4632 42524 4644
rect 42576 4632 42582 4684
rect 44082 4672 44088 4684
rect 44043 4644 44088 4672
rect 44082 4632 44088 4644
rect 44140 4632 44146 4684
rect 3237 4607 3295 4613
rect 3237 4573 3249 4607
rect 3283 4573 3295 4607
rect 3237 4567 3295 4573
rect 6270 4564 6276 4616
rect 6328 4604 6334 4616
rect 6365 4607 6423 4613
rect 6365 4604 6377 4607
rect 6328 4576 6377 4604
rect 6328 4564 6334 4576
rect 6365 4573 6377 4576
rect 6411 4573 6423 4607
rect 37366 4604 37372 4616
rect 37327 4576 37372 4604
rect 6365 4567 6423 4573
rect 37366 4564 37372 4576
rect 37424 4564 37430 4616
rect 37550 4536 37556 4548
rect 37511 4508 37556 4536
rect 37550 4496 37556 4508
rect 37608 4496 37614 4548
rect 3145 4471 3203 4477
rect 3145 4437 3157 4471
rect 3191 4468 3203 4471
rect 4154 4468 4160 4480
rect 3191 4440 4160 4468
rect 3191 4437 3203 4440
rect 3145 4431 3203 4437
rect 4154 4428 4160 4440
rect 4212 4428 4218 4480
rect 1104 4378 44896 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 44896 4378
rect 1104 4304 44896 4326
rect 2038 4128 2044 4140
rect 1999 4100 2044 4128
rect 2038 4088 2044 4100
rect 2096 4088 2102 4140
rect 4341 4131 4399 4137
rect 4341 4097 4353 4131
rect 4387 4128 4399 4131
rect 4890 4128 4896 4140
rect 4387 4100 4896 4128
rect 4387 4097 4399 4100
rect 4341 4091 4399 4097
rect 4890 4088 4896 4100
rect 4948 4088 4954 4140
rect 5353 4131 5411 4137
rect 5353 4097 5365 4131
rect 5399 4097 5411 4131
rect 11790 4128 11796 4140
rect 11751 4100 11796 4128
rect 5353 4091 5411 4097
rect 2774 4020 2780 4072
rect 2832 4060 2838 4072
rect 4154 4060 4160 4072
rect 2832 4032 2877 4060
rect 4115 4032 4160 4060
rect 2832 4020 2838 4032
rect 4154 4020 4160 4032
rect 4212 4020 4218 4072
rect 5368 4060 5396 4091
rect 11790 4088 11796 4100
rect 11848 4128 11854 4140
rect 11848 4100 16574 4128
rect 11848 4088 11854 4100
rect 16546 4060 16574 4100
rect 18690 4088 18696 4140
rect 18748 4128 18754 4140
rect 20993 4131 21051 4137
rect 20993 4128 21005 4131
rect 18748 4100 21005 4128
rect 18748 4088 18754 4100
rect 20993 4097 21005 4100
rect 21039 4097 21051 4131
rect 36538 4128 36544 4140
rect 36499 4100 36544 4128
rect 20993 4091 21051 4097
rect 36538 4088 36544 4100
rect 36596 4088 36602 4140
rect 37366 4088 37372 4140
rect 37424 4128 37430 4140
rect 37921 4131 37979 4137
rect 37921 4128 37933 4131
rect 37424 4100 37933 4128
rect 37424 4088 37430 4100
rect 37921 4097 37933 4100
rect 37967 4097 37979 4131
rect 37921 4091 37979 4097
rect 41693 4131 41751 4137
rect 41693 4097 41705 4131
rect 41739 4128 41751 4131
rect 42978 4128 42984 4140
rect 41739 4100 42984 4128
rect 41739 4097 41751 4100
rect 41693 4091 41751 4097
rect 42978 4088 42984 4100
rect 43036 4088 43042 4140
rect 43346 4128 43352 4140
rect 43307 4100 43352 4128
rect 43346 4088 43352 4100
rect 43404 4088 43410 4140
rect 38194 4060 38200 4072
rect 5368 4032 12434 4060
rect 16546 4032 38200 4060
rect 2314 3952 2320 4004
rect 2372 3992 2378 4004
rect 5368 3992 5396 4032
rect 2372 3964 5396 3992
rect 2372 3952 2378 3964
rect 6178 3952 6184 4004
rect 6236 3992 6242 4004
rect 9490 3992 9496 4004
rect 6236 3964 9496 3992
rect 6236 3952 6242 3964
rect 9490 3952 9496 3964
rect 9548 3952 9554 4004
rect 12406 3992 12434 4032
rect 38194 4020 38200 4032
rect 38252 4020 38258 4072
rect 38838 4060 38844 4072
rect 38799 4032 38844 4060
rect 38838 4020 38844 4032
rect 38896 4020 38902 4072
rect 39025 4063 39083 4069
rect 39025 4029 39037 4063
rect 39071 4029 39083 4063
rect 39025 4023 39083 4029
rect 40681 4063 40739 4069
rect 40681 4029 40693 4063
rect 40727 4060 40739 4063
rect 41322 4060 41328 4072
rect 40727 4032 41328 4060
rect 40727 4029 40739 4032
rect 40681 4023 40739 4029
rect 36446 3992 36452 4004
rect 12406 3964 36452 3992
rect 36446 3952 36452 3964
rect 36504 3952 36510 4004
rect 36633 3995 36691 4001
rect 36633 3961 36645 3995
rect 36679 3992 36691 3995
rect 37458 3992 37464 4004
rect 36679 3964 37464 3992
rect 36679 3961 36691 3964
rect 36633 3955 36691 3961
rect 37458 3952 37464 3964
rect 37516 3952 37522 4004
rect 38286 3952 38292 4004
rect 38344 3992 38350 4004
rect 39040 3992 39068 4023
rect 41322 4020 41328 4032
rect 41380 4020 41386 4072
rect 38344 3964 39068 3992
rect 38344 3952 38350 3964
rect 1578 3884 1584 3936
rect 1636 3924 1642 3936
rect 1949 3927 2007 3933
rect 1949 3924 1961 3927
rect 1636 3896 1961 3924
rect 1636 3884 1642 3896
rect 1949 3893 1961 3896
rect 1995 3893 2007 3927
rect 1949 3887 2007 3893
rect 3878 3884 3884 3936
rect 3936 3924 3942 3936
rect 4706 3924 4712 3936
rect 3936 3896 4712 3924
rect 3936 3884 3942 3896
rect 4706 3884 4712 3896
rect 4764 3884 4770 3936
rect 5445 3927 5503 3933
rect 5445 3893 5457 3927
rect 5491 3924 5503 3927
rect 5534 3924 5540 3936
rect 5491 3896 5540 3924
rect 5491 3893 5503 3896
rect 5445 3887 5503 3893
rect 5534 3884 5540 3896
rect 5592 3884 5598 3936
rect 6362 3924 6368 3936
rect 6323 3896 6368 3924
rect 6362 3884 6368 3896
rect 6420 3884 6426 3936
rect 7282 3884 7288 3936
rect 7340 3924 7346 3936
rect 7377 3927 7435 3933
rect 7377 3924 7389 3927
rect 7340 3896 7389 3924
rect 7340 3884 7346 3896
rect 7377 3893 7389 3896
rect 7423 3893 7435 3927
rect 7377 3887 7435 3893
rect 9214 3884 9220 3936
rect 9272 3924 9278 3936
rect 9309 3927 9367 3933
rect 9309 3924 9321 3927
rect 9272 3896 9321 3924
rect 9272 3884 9278 3896
rect 9309 3893 9321 3896
rect 9355 3893 9367 3927
rect 11882 3924 11888 3936
rect 11843 3896 11888 3924
rect 9309 3887 9367 3893
rect 11882 3884 11888 3896
rect 11940 3884 11946 3936
rect 12434 3924 12440 3936
rect 12395 3896 12440 3924
rect 12434 3884 12440 3896
rect 12492 3884 12498 3936
rect 15470 3884 15476 3936
rect 15528 3924 15534 3936
rect 15565 3927 15623 3933
rect 15565 3924 15577 3927
rect 15528 3896 15577 3924
rect 15528 3884 15534 3896
rect 15565 3893 15577 3896
rect 15611 3893 15623 3927
rect 15565 3887 15623 3893
rect 20806 3884 20812 3936
rect 20864 3924 20870 3936
rect 20901 3927 20959 3933
rect 20901 3924 20913 3927
rect 20864 3896 20913 3924
rect 20864 3884 20870 3896
rect 20901 3893 20913 3896
rect 20947 3893 20959 3927
rect 24210 3924 24216 3936
rect 24171 3896 24216 3924
rect 20901 3887 20959 3893
rect 24210 3884 24216 3896
rect 24268 3884 24274 3936
rect 37274 3924 37280 3936
rect 37235 3896 37280 3924
rect 37274 3884 37280 3896
rect 37332 3884 37338 3936
rect 41785 3927 41843 3933
rect 41785 3893 41797 3927
rect 41831 3924 41843 3927
rect 41874 3924 41880 3936
rect 41831 3896 41880 3924
rect 41831 3893 41843 3896
rect 41785 3887 41843 3893
rect 41874 3884 41880 3896
rect 41932 3884 41938 3936
rect 42426 3924 42432 3936
rect 42387 3896 42432 3924
rect 42426 3884 42432 3896
rect 42484 3884 42490 3936
rect 43438 3924 43444 3936
rect 43399 3896 43444 3924
rect 43438 3884 43444 3896
rect 43496 3884 43502 3936
rect 43530 3884 43536 3936
rect 43588 3924 43594 3936
rect 43993 3927 44051 3933
rect 43993 3924 44005 3927
rect 43588 3896 44005 3924
rect 43588 3884 43594 3896
rect 43993 3893 44005 3896
rect 44039 3893 44051 3927
rect 43993 3887 44051 3893
rect 1104 3834 44896 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 44896 3834
rect 1104 3760 44896 3782
rect 12802 3720 12808 3732
rect 8312 3692 12808 3720
rect 6362 3652 6368 3664
rect 5368 3624 6368 3652
rect 2958 3544 2964 3596
rect 3016 3584 3022 3596
rect 5368 3593 5396 3624
rect 6362 3612 6368 3624
rect 6420 3612 6426 3664
rect 3237 3587 3295 3593
rect 3237 3584 3249 3587
rect 3016 3556 3249 3584
rect 3016 3544 3022 3556
rect 3237 3553 3249 3556
rect 3283 3553 3295 3587
rect 3237 3547 3295 3553
rect 5353 3587 5411 3593
rect 5353 3553 5365 3587
rect 5399 3553 5411 3587
rect 5534 3584 5540 3596
rect 5495 3556 5540 3584
rect 5353 3547 5411 3553
rect 5534 3544 5540 3556
rect 5592 3544 5598 3596
rect 5810 3584 5816 3596
rect 5771 3556 5816 3584
rect 5810 3544 5816 3556
rect 5868 3544 5874 3596
rect 1394 3516 1400 3528
rect 1355 3488 1400 3516
rect 1394 3476 1400 3488
rect 1452 3476 1458 3528
rect 4522 3516 4528 3528
rect 4483 3488 4528 3516
rect 4522 3476 4528 3488
rect 4580 3476 4586 3528
rect 8312 3525 8340 3692
rect 12802 3680 12808 3692
rect 12860 3720 12866 3732
rect 13262 3720 13268 3732
rect 12860 3692 13268 3720
rect 12860 3680 12866 3692
rect 13262 3680 13268 3692
rect 13320 3680 13326 3732
rect 38286 3720 38292 3732
rect 38247 3692 38292 3720
rect 38286 3680 38292 3692
rect 38344 3680 38350 3732
rect 38838 3720 38844 3732
rect 38799 3692 38844 3720
rect 38838 3680 38844 3692
rect 38896 3680 38902 3732
rect 42794 3720 42800 3732
rect 40880 3692 42800 3720
rect 9490 3612 9496 3664
rect 9548 3652 9554 3664
rect 36538 3652 36544 3664
rect 9548 3624 36544 3652
rect 9548 3612 9554 3624
rect 9214 3544 9220 3596
rect 9272 3584 9278 3596
rect 9398 3584 9404 3596
rect 9272 3556 9317 3584
rect 9359 3556 9404 3584
rect 9272 3544 9278 3556
rect 9398 3544 9404 3556
rect 9456 3544 9462 3596
rect 9674 3584 9680 3596
rect 9635 3556 9680 3584
rect 9674 3544 9680 3556
rect 9732 3544 9738 3596
rect 12986 3584 12992 3596
rect 12406 3556 12992 3584
rect 8297 3519 8355 3525
rect 8297 3485 8309 3519
rect 8343 3485 8355 3519
rect 8297 3479 8355 3485
rect 12253 3519 12311 3525
rect 12253 3485 12265 3519
rect 12299 3516 12311 3519
rect 12406 3516 12434 3556
rect 12986 3544 12992 3556
rect 13044 3544 13050 3596
rect 15470 3584 15476 3596
rect 15431 3556 15476 3584
rect 15470 3544 15476 3556
rect 15528 3544 15534 3596
rect 16114 3584 16120 3596
rect 16075 3556 16120 3584
rect 16114 3544 16120 3556
rect 16172 3544 16178 3596
rect 12299 3488 12434 3516
rect 12897 3519 12955 3525
rect 12299 3485 12311 3488
rect 12253 3479 12311 3485
rect 12897 3485 12909 3519
rect 12943 3516 12955 3519
rect 13354 3516 13360 3528
rect 12943 3488 13360 3516
rect 12943 3485 12955 3488
rect 12897 3479 12955 3485
rect 13354 3476 13360 3488
rect 13412 3476 13418 3528
rect 16850 3476 16856 3528
rect 16908 3516 16914 3528
rect 17773 3519 17831 3525
rect 17773 3516 17785 3519
rect 16908 3488 17785 3516
rect 16908 3476 16914 3488
rect 17773 3485 17785 3488
rect 17819 3485 17831 3519
rect 17773 3479 17831 3485
rect 18693 3519 18751 3525
rect 18693 3485 18705 3519
rect 18739 3516 18751 3519
rect 18782 3516 18788 3528
rect 18739 3488 18788 3516
rect 18739 3485 18751 3488
rect 18693 3479 18751 3485
rect 18782 3476 18788 3488
rect 18840 3476 18846 3528
rect 19444 3525 19472 3624
rect 36538 3612 36544 3624
rect 36596 3612 36602 3664
rect 20806 3584 20812 3596
rect 20767 3556 20812 3584
rect 20806 3544 20812 3556
rect 20864 3544 20870 3596
rect 21266 3584 21272 3596
rect 21227 3556 21272 3584
rect 21266 3544 21272 3556
rect 21324 3544 21330 3596
rect 24780 3556 29776 3584
rect 24780 3528 24808 3556
rect 19429 3519 19487 3525
rect 19429 3485 19441 3519
rect 19475 3485 19487 3519
rect 19429 3479 19487 3485
rect 20165 3519 20223 3525
rect 20165 3485 20177 3519
rect 20211 3516 20223 3519
rect 20625 3519 20683 3525
rect 20625 3516 20637 3519
rect 20211 3488 20637 3516
rect 20211 3485 20223 3488
rect 20165 3479 20223 3485
rect 20625 3485 20637 3488
rect 20671 3485 20683 3519
rect 20625 3479 20683 3485
rect 22094 3476 22100 3528
rect 22152 3516 22158 3528
rect 22925 3519 22983 3525
rect 22925 3516 22937 3519
rect 22152 3488 22937 3516
rect 22152 3476 22158 3488
rect 22925 3485 22937 3488
rect 22971 3485 22983 3519
rect 22925 3479 22983 3485
rect 23661 3519 23719 3525
rect 23661 3485 23673 3519
rect 23707 3485 23719 3519
rect 24762 3516 24768 3528
rect 24723 3488 24768 3516
rect 23661 3479 23719 3485
rect 2222 3408 2228 3460
rect 2280 3448 2286 3460
rect 3053 3451 3111 3457
rect 3053 3448 3065 3451
rect 2280 3420 3065 3448
rect 2280 3408 2286 3420
rect 3053 3417 3065 3420
rect 3099 3417 3111 3451
rect 3053 3411 3111 3417
rect 3694 3408 3700 3460
rect 3752 3448 3758 3460
rect 13078 3448 13084 3460
rect 3752 3420 13084 3448
rect 3752 3408 3758 3420
rect 13078 3408 13084 3420
rect 13136 3408 13142 3460
rect 15657 3451 15715 3457
rect 15657 3417 15669 3451
rect 15703 3448 15715 3451
rect 15746 3448 15752 3460
rect 15703 3420 15752 3448
rect 15703 3417 15715 3420
rect 15657 3411 15715 3417
rect 15746 3408 15752 3420
rect 15804 3408 15810 3460
rect 23676 3448 23704 3479
rect 24762 3476 24768 3488
rect 24820 3476 24826 3528
rect 25225 3519 25283 3525
rect 25225 3485 25237 3519
rect 25271 3485 25283 3519
rect 25225 3479 25283 3485
rect 28997 3519 29055 3525
rect 28997 3485 29009 3519
rect 29043 3516 29055 3519
rect 29178 3516 29184 3528
rect 29043 3488 29184 3516
rect 29043 3485 29055 3488
rect 28997 3479 29055 3485
rect 16546 3420 23704 3448
rect 4433 3383 4491 3389
rect 4433 3349 4445 3383
rect 4479 3380 4491 3383
rect 4614 3380 4620 3392
rect 4479 3352 4620 3380
rect 4479 3349 4491 3352
rect 4433 3343 4491 3349
rect 4614 3340 4620 3352
rect 4672 3340 4678 3392
rect 7466 3340 7472 3392
rect 7524 3380 7530 3392
rect 8205 3383 8263 3389
rect 8205 3380 8217 3383
rect 7524 3352 8217 3380
rect 7524 3340 7530 3352
rect 8205 3349 8217 3352
rect 8251 3349 8263 3383
rect 8205 3343 8263 3349
rect 12161 3383 12219 3389
rect 12161 3349 12173 3383
rect 12207 3380 12219 3383
rect 13170 3380 13176 3392
rect 12207 3352 13176 3380
rect 12207 3349 12219 3352
rect 12161 3343 12219 3349
rect 13170 3340 13176 3352
rect 13228 3340 13234 3392
rect 13262 3340 13268 3392
rect 13320 3380 13326 3392
rect 16546 3380 16574 3420
rect 24394 3408 24400 3460
rect 24452 3448 24458 3460
rect 25240 3448 25268 3479
rect 29178 3476 29184 3488
rect 29236 3476 29242 3528
rect 29748 3525 29776 3556
rect 35526 3544 35532 3596
rect 35584 3584 35590 3596
rect 35805 3587 35863 3593
rect 35805 3584 35817 3587
rect 35584 3556 35817 3584
rect 35584 3544 35590 3556
rect 35805 3553 35817 3556
rect 35851 3553 35863 3587
rect 36078 3584 36084 3596
rect 36039 3556 36084 3584
rect 35805 3547 35863 3553
rect 36078 3544 36084 3556
rect 36136 3544 36142 3596
rect 36446 3544 36452 3596
rect 36504 3584 36510 3596
rect 40880 3584 40908 3692
rect 42794 3680 42800 3692
rect 42852 3680 42858 3732
rect 43990 3680 43996 3732
rect 44048 3720 44054 3732
rect 44085 3723 44143 3729
rect 44085 3720 44097 3723
rect 44048 3692 44097 3720
rect 44048 3680 44054 3692
rect 44085 3689 44097 3692
rect 44131 3689 44143 3723
rect 44085 3683 44143 3689
rect 42426 3652 42432 3664
rect 41708 3624 42432 3652
rect 41708 3593 41736 3624
rect 42426 3612 42432 3624
rect 42484 3612 42490 3664
rect 36504 3556 40908 3584
rect 36504 3544 36510 3556
rect 29733 3519 29791 3525
rect 29733 3485 29745 3519
rect 29779 3485 29791 3519
rect 35618 3516 35624 3528
rect 35579 3488 35624 3516
rect 29733 3479 29791 3485
rect 35618 3476 35624 3488
rect 35676 3476 35682 3528
rect 38194 3516 38200 3528
rect 38155 3488 38200 3516
rect 38194 3476 38200 3488
rect 38252 3476 38258 3528
rect 40034 3516 40040 3528
rect 39995 3488 40040 3516
rect 40034 3476 40040 3488
rect 40092 3476 40098 3528
rect 40880 3525 40908 3556
rect 41693 3587 41751 3593
rect 41693 3553 41705 3587
rect 41739 3553 41751 3587
rect 41874 3584 41880 3596
rect 41835 3556 41880 3584
rect 41693 3547 41751 3553
rect 41874 3544 41880 3556
rect 41932 3544 41938 3596
rect 42518 3584 42524 3596
rect 42479 3556 42524 3584
rect 42518 3544 42524 3556
rect 42576 3544 42582 3596
rect 40865 3519 40923 3525
rect 40865 3485 40877 3519
rect 40911 3485 40923 3519
rect 40865 3479 40923 3485
rect 43898 3476 43904 3528
rect 43956 3516 43962 3528
rect 43993 3519 44051 3525
rect 43993 3516 44005 3519
rect 43956 3488 44005 3516
rect 43956 3476 43962 3488
rect 43993 3485 44005 3488
rect 44039 3485 44051 3519
rect 43993 3479 44051 3485
rect 24452 3420 25268 3448
rect 24452 3408 24458 3420
rect 37366 3408 37372 3460
rect 37424 3448 37430 3460
rect 39942 3448 39948 3460
rect 37424 3420 39948 3448
rect 37424 3408 37430 3420
rect 39942 3408 39948 3420
rect 40000 3408 40006 3460
rect 42886 3448 42892 3460
rect 40144 3420 42892 3448
rect 13320 3352 16574 3380
rect 13320 3340 13326 3352
rect 18966 3340 18972 3392
rect 19024 3380 19030 3392
rect 19337 3383 19395 3389
rect 19337 3380 19349 3383
rect 19024 3352 19349 3380
rect 19024 3340 19030 3352
rect 19337 3349 19349 3352
rect 19383 3349 19395 3383
rect 23750 3380 23756 3392
rect 23711 3352 23756 3380
rect 19337 3343 19395 3349
rect 23750 3340 23756 3352
rect 23808 3340 23814 3392
rect 24578 3340 24584 3392
rect 24636 3380 24642 3392
rect 24673 3383 24731 3389
rect 24673 3380 24685 3383
rect 24636 3352 24685 3380
rect 24636 3340 24642 3352
rect 24673 3349 24685 3352
rect 24719 3349 24731 3383
rect 24673 3343 24731 3349
rect 29362 3340 29368 3392
rect 29420 3380 29426 3392
rect 29641 3383 29699 3389
rect 29641 3380 29653 3383
rect 29420 3352 29653 3380
rect 29420 3340 29426 3352
rect 29641 3349 29653 3352
rect 29687 3349 29699 3383
rect 29641 3343 29699 3349
rect 36538 3340 36544 3392
rect 36596 3380 36602 3392
rect 40144 3380 40172 3420
rect 42886 3408 42892 3420
rect 42944 3408 42950 3460
rect 36596 3352 40172 3380
rect 36596 3340 36602 3352
rect 40218 3340 40224 3392
rect 40276 3380 40282 3392
rect 40773 3383 40831 3389
rect 40773 3380 40785 3383
rect 40276 3352 40785 3380
rect 40276 3340 40282 3352
rect 40773 3349 40785 3352
rect 40819 3349 40831 3383
rect 40773 3343 40831 3349
rect 1104 3290 44896 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 44896 3290
rect 1104 3216 44896 3238
rect 2222 3176 2228 3188
rect 2183 3148 2228 3176
rect 2222 3136 2228 3148
rect 2280 3136 2286 3188
rect 4522 3136 4528 3188
rect 4580 3176 4586 3188
rect 9582 3176 9588 3188
rect 4580 3148 9588 3176
rect 4580 3136 4586 3148
rect 2961 3111 3019 3117
rect 2961 3077 2973 3111
rect 3007 3108 3019 3111
rect 3697 3111 3755 3117
rect 3697 3108 3709 3111
rect 3007 3080 3709 3108
rect 3007 3077 3019 3080
rect 2961 3071 3019 3077
rect 3697 3077 3709 3080
rect 3743 3077 3755 3111
rect 3697 3071 3755 3077
rect 2314 3040 2320 3052
rect 2275 3012 2320 3040
rect 2314 3000 2320 3012
rect 2372 3000 2378 3052
rect 3053 3043 3111 3049
rect 3053 3009 3065 3043
rect 3099 3009 3111 3043
rect 3053 3003 3111 3009
rect 3068 2972 3096 3003
rect 3142 3000 3148 3052
rect 3200 3040 3206 3052
rect 6380 3049 6408 3148
rect 9582 3136 9588 3148
rect 9640 3136 9646 3188
rect 15746 3176 15752 3188
rect 12406 3148 13584 3176
rect 15707 3148 15752 3176
rect 7466 3108 7472 3120
rect 7427 3080 7472 3108
rect 7466 3068 7472 3080
rect 7524 3068 7530 3120
rect 12406 3108 12434 3148
rect 13170 3108 13176 3120
rect 8680 3080 12434 3108
rect 13131 3080 13176 3108
rect 3513 3043 3571 3049
rect 3513 3040 3525 3043
rect 3200 3012 3525 3040
rect 3200 3000 3206 3012
rect 3513 3009 3525 3012
rect 3559 3009 3571 3043
rect 3513 3003 3571 3009
rect 6365 3043 6423 3049
rect 6365 3009 6377 3043
rect 6411 3009 6423 3043
rect 7282 3040 7288 3052
rect 7243 3012 7288 3040
rect 6365 3003 6423 3009
rect 7282 3000 7288 3012
rect 7340 3000 7346 3052
rect 3694 2972 3700 2984
rect 3068 2944 3700 2972
rect 3694 2932 3700 2944
rect 3752 2932 3758 2984
rect 3970 2972 3976 2984
rect 3931 2944 3976 2972
rect 3970 2932 3976 2944
rect 4028 2932 4034 2984
rect 7098 2932 7104 2984
rect 7156 2972 7162 2984
rect 7745 2975 7803 2981
rect 7745 2972 7757 2975
rect 7156 2944 7757 2972
rect 7156 2932 7162 2944
rect 7745 2941 7757 2944
rect 7791 2941 7803 2975
rect 7745 2935 7803 2941
rect 658 2864 664 2916
rect 716 2904 722 2916
rect 4706 2904 4712 2916
rect 716 2876 4712 2904
rect 716 2864 722 2876
rect 4706 2864 4712 2876
rect 4764 2864 4770 2916
rect 5166 2864 5172 2916
rect 5224 2904 5230 2916
rect 8680 2904 8708 3080
rect 13170 3068 13176 3080
rect 13228 3068 13234 3120
rect 13354 3000 13360 3052
rect 13412 3040 13418 3052
rect 13556 3040 13584 3148
rect 15746 3136 15752 3148
rect 15804 3136 15810 3188
rect 36633 3179 36691 3185
rect 36633 3145 36645 3179
rect 36679 3176 36691 3179
rect 37550 3176 37556 3188
rect 36679 3148 37556 3176
rect 36679 3145 36691 3148
rect 36633 3139 36691 3145
rect 37550 3136 37556 3148
rect 37608 3136 37614 3188
rect 42978 3176 42984 3188
rect 39776 3148 42984 3176
rect 18690 3108 18696 3120
rect 16546 3080 18696 3108
rect 15841 3043 15899 3049
rect 15841 3040 15853 3043
rect 13412 3012 13457 3040
rect 13556 3012 15853 3040
rect 13412 3000 13418 3012
rect 15841 3009 15853 3012
rect 15887 3040 15899 3043
rect 16546 3040 16574 3080
rect 18690 3068 18696 3080
rect 18748 3068 18754 3120
rect 18966 3108 18972 3120
rect 18927 3080 18972 3108
rect 18966 3068 18972 3080
rect 19024 3068 19030 3120
rect 24578 3108 24584 3120
rect 24539 3080 24584 3108
rect 24578 3068 24584 3080
rect 24636 3068 24642 3120
rect 29362 3108 29368 3120
rect 29323 3080 29368 3108
rect 29362 3068 29368 3080
rect 29420 3068 29426 3120
rect 15887 3012 16574 3040
rect 16945 3043 17003 3049
rect 15887 3009 15899 3012
rect 15841 3003 15899 3009
rect 16945 3009 16957 3043
rect 16991 3009 17003 3043
rect 18782 3040 18788 3052
rect 18743 3012 18788 3040
rect 16945 3003 17003 3009
rect 11606 2972 11612 2984
rect 11567 2944 11612 2972
rect 11606 2932 11612 2944
rect 11664 2932 11670 2984
rect 11698 2932 11704 2984
rect 11756 2972 11762 2984
rect 16960 2972 16988 3003
rect 18782 3000 18788 3012
rect 18840 3000 18846 3052
rect 22094 3040 22100 3052
rect 22055 3012 22100 3040
rect 22094 3000 22100 3012
rect 22152 3000 22158 3052
rect 24394 3040 24400 3052
rect 24355 3012 24400 3040
rect 24394 3000 24400 3012
rect 24452 3000 24458 3052
rect 29178 3040 29184 3052
rect 29139 3012 29184 3040
rect 29178 3000 29184 3012
rect 29236 3000 29242 3052
rect 35618 3000 35624 3052
rect 35676 3040 35682 3052
rect 35713 3043 35771 3049
rect 35713 3040 35725 3043
rect 35676 3012 35725 3040
rect 35676 3000 35682 3012
rect 35713 3009 35725 3012
rect 35759 3009 35771 3043
rect 36538 3040 36544 3052
rect 36499 3012 36544 3040
rect 35713 3003 35771 3009
rect 36538 3000 36544 3012
rect 36596 3000 36602 3052
rect 39577 3043 39635 3049
rect 39577 3009 39589 3043
rect 39623 3040 39635 3043
rect 39776 3040 39804 3148
rect 42978 3136 42984 3148
rect 43036 3136 43042 3188
rect 40034 3040 40040 3052
rect 39623 3012 39804 3040
rect 39995 3012 40040 3040
rect 39623 3009 39635 3012
rect 39577 3003 39635 3009
rect 40034 3000 40040 3012
rect 40092 3000 40098 3052
rect 42886 3000 42892 3052
rect 42944 3040 42950 3052
rect 42981 3043 43039 3049
rect 42981 3040 42993 3043
rect 42944 3012 42993 3040
rect 42944 3000 42950 3012
rect 42981 3009 42993 3012
rect 43027 3009 43039 3043
rect 42981 3003 43039 3009
rect 43809 3043 43867 3049
rect 43809 3009 43821 3043
rect 43855 3040 43867 3043
rect 44174 3040 44180 3052
rect 43855 3012 44180 3040
rect 43855 3009 43867 3012
rect 43809 3003 43867 3009
rect 44174 3000 44180 3012
rect 44232 3000 44238 3052
rect 19334 2972 19340 2984
rect 11756 2944 16988 2972
rect 19295 2944 19340 2972
rect 11756 2932 11762 2944
rect 5224 2876 8708 2904
rect 16960 2904 16988 2944
rect 19334 2932 19340 2944
rect 19392 2932 19398 2984
rect 22278 2972 22284 2984
rect 22239 2944 22284 2972
rect 22278 2932 22284 2944
rect 22336 2932 22342 2984
rect 23198 2972 23204 2984
rect 23159 2944 23204 2972
rect 23198 2932 23204 2944
rect 23256 2932 23262 2984
rect 25130 2972 25136 2984
rect 25091 2944 25136 2972
rect 25130 2932 25136 2944
rect 25188 2932 25194 2984
rect 29638 2972 29644 2984
rect 29599 2944 29644 2972
rect 29638 2932 29644 2944
rect 29696 2932 29702 2984
rect 39117 2975 39175 2981
rect 39117 2941 39129 2975
rect 39163 2941 39175 2975
rect 39117 2935 39175 2941
rect 39393 2975 39451 2981
rect 39393 2941 39405 2975
rect 39439 2941 39451 2975
rect 40218 2972 40224 2984
rect 40179 2944 40224 2972
rect 39393 2935 39451 2941
rect 23014 2904 23020 2916
rect 16960 2876 23020 2904
rect 5224 2864 5230 2876
rect 23014 2864 23020 2876
rect 23072 2864 23078 2916
rect 1394 2796 1400 2848
rect 1452 2836 1458 2848
rect 1489 2839 1547 2845
rect 1489 2836 1501 2839
rect 1452 2808 1501 2836
rect 1452 2796 1458 2808
rect 1489 2805 1501 2808
rect 1535 2805 1547 2839
rect 1489 2799 1547 2805
rect 3234 2796 3240 2848
rect 3292 2836 3298 2848
rect 3970 2836 3976 2848
rect 3292 2808 3976 2836
rect 3292 2796 3298 2808
rect 3970 2796 3976 2808
rect 4028 2796 4034 2848
rect 6457 2839 6515 2845
rect 6457 2805 6469 2839
rect 6503 2836 6515 2839
rect 6546 2836 6552 2848
rect 6503 2808 6552 2836
rect 6503 2805 6515 2808
rect 6457 2799 6515 2805
rect 6546 2796 6552 2808
rect 6604 2796 6610 2848
rect 17034 2836 17040 2848
rect 16995 2808 17040 2836
rect 17034 2796 17040 2808
rect 17092 2796 17098 2848
rect 39132 2836 39160 2935
rect 39408 2904 39436 2935
rect 40218 2932 40224 2944
rect 40276 2932 40282 2984
rect 41230 2972 41236 2984
rect 41191 2944 41236 2972
rect 41230 2932 41236 2944
rect 41288 2932 41294 2984
rect 42889 2907 42947 2913
rect 42889 2904 42901 2907
rect 39408 2876 42901 2904
rect 42889 2873 42901 2876
rect 42935 2873 42947 2907
rect 42889 2867 42947 2873
rect 43806 2836 43812 2848
rect 39132 2808 43812 2836
rect 43806 2796 43812 2808
rect 43864 2796 43870 2848
rect 1104 2746 44896 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 44896 2746
rect 1104 2672 44896 2694
rect 3418 2592 3424 2644
rect 3476 2632 3482 2644
rect 15930 2632 15936 2644
rect 3476 2604 15936 2632
rect 3476 2592 3482 2604
rect 15930 2592 15936 2604
rect 15988 2592 15994 2644
rect 22278 2592 22284 2644
rect 22336 2632 22342 2644
rect 22925 2635 22983 2641
rect 22925 2632 22937 2635
rect 22336 2604 22937 2632
rect 22336 2592 22342 2604
rect 22925 2601 22937 2604
rect 22971 2601 22983 2635
rect 42978 2632 42984 2644
rect 42939 2604 42984 2632
rect 22925 2595 22983 2601
rect 42978 2592 42984 2604
rect 43036 2592 43042 2644
rect 12434 2564 12440 2576
rect 11716 2536 12440 2564
rect 1394 2496 1400 2508
rect 1355 2468 1400 2496
rect 1394 2456 1400 2468
rect 1452 2456 1458 2508
rect 1578 2496 1584 2508
rect 1539 2468 1584 2496
rect 1578 2456 1584 2468
rect 1636 2456 1642 2508
rect 2774 2496 2780 2508
rect 2735 2468 2780 2496
rect 2774 2456 2780 2468
rect 2832 2456 2838 2508
rect 3786 2496 3792 2508
rect 3747 2468 3792 2496
rect 3786 2456 3792 2468
rect 3844 2456 3850 2508
rect 3973 2499 4031 2505
rect 3973 2465 3985 2499
rect 4019 2496 4031 2499
rect 4614 2496 4620 2508
rect 4019 2468 4620 2496
rect 4019 2465 4031 2468
rect 3973 2459 4031 2465
rect 4614 2456 4620 2468
rect 4672 2456 4678 2508
rect 4706 2456 4712 2508
rect 4764 2496 4770 2508
rect 6362 2496 6368 2508
rect 4764 2468 4809 2496
rect 6323 2468 6368 2496
rect 4764 2456 4770 2468
rect 6362 2456 6368 2468
rect 6420 2456 6426 2508
rect 6546 2496 6552 2508
rect 6507 2468 6552 2496
rect 6546 2456 6552 2468
rect 6604 2456 6610 2508
rect 6638 2456 6644 2508
rect 6696 2496 6702 2508
rect 11716 2505 11744 2536
rect 12434 2524 12440 2536
rect 12492 2524 12498 2576
rect 23014 2564 23020 2576
rect 22927 2536 23020 2564
rect 23014 2524 23020 2536
rect 23072 2564 23078 2576
rect 43346 2564 43352 2576
rect 23072 2536 43352 2564
rect 23072 2524 23078 2536
rect 43346 2524 43352 2536
rect 43404 2524 43410 2576
rect 6917 2499 6975 2505
rect 6917 2496 6929 2499
rect 6696 2468 6929 2496
rect 6696 2456 6702 2468
rect 6917 2465 6929 2468
rect 6963 2465 6975 2499
rect 6917 2459 6975 2465
rect 11701 2499 11759 2505
rect 11701 2465 11713 2499
rect 11747 2465 11759 2499
rect 11882 2496 11888 2508
rect 11843 2468 11888 2496
rect 11701 2459 11759 2465
rect 11882 2456 11888 2468
rect 11940 2456 11946 2508
rect 12250 2496 12256 2508
rect 12211 2468 12256 2496
rect 12250 2456 12256 2468
rect 12308 2456 12314 2508
rect 16850 2496 16856 2508
rect 16811 2468 16856 2496
rect 16850 2456 16856 2468
rect 16908 2456 16914 2508
rect 17034 2496 17040 2508
rect 16995 2468 17040 2496
rect 17034 2456 17040 2468
rect 17092 2456 17098 2508
rect 17402 2496 17408 2508
rect 17363 2468 17408 2496
rect 17402 2456 17408 2468
rect 17460 2456 17466 2508
rect 23032 2437 23060 2524
rect 24210 2456 24216 2508
rect 24268 2496 24274 2508
rect 24397 2499 24455 2505
rect 24397 2496 24409 2499
rect 24268 2468 24409 2496
rect 24268 2456 24274 2468
rect 24397 2465 24409 2468
rect 24443 2465 24455 2499
rect 24397 2459 24455 2465
rect 24578 2456 24584 2508
rect 24636 2496 24642 2508
rect 24857 2499 24915 2505
rect 24857 2496 24869 2499
rect 24636 2468 24869 2496
rect 24636 2456 24642 2468
rect 24857 2465 24869 2468
rect 24903 2465 24915 2499
rect 37274 2496 37280 2508
rect 37235 2468 37280 2496
rect 24857 2459 24915 2465
rect 37274 2456 37280 2468
rect 37332 2456 37338 2508
rect 37458 2496 37464 2508
rect 37419 2468 37464 2496
rect 37458 2456 37464 2468
rect 37516 2456 37522 2508
rect 38654 2496 38660 2508
rect 38615 2468 38660 2496
rect 38654 2456 38660 2468
rect 38712 2456 38718 2508
rect 41322 2496 41328 2508
rect 41283 2468 41328 2496
rect 41322 2456 41328 2468
rect 41380 2456 41386 2508
rect 41693 2499 41751 2505
rect 41693 2465 41705 2499
rect 41739 2496 41751 2499
rect 43438 2496 43444 2508
rect 41739 2468 43444 2496
rect 41739 2465 41751 2468
rect 41693 2459 41751 2465
rect 43438 2456 43444 2468
rect 43496 2456 43502 2508
rect 23017 2431 23075 2437
rect 23017 2397 23029 2431
rect 23063 2397 23075 2431
rect 23017 2391 23075 2397
rect 41877 2431 41935 2437
rect 41877 2397 41889 2431
rect 41923 2428 41935 2431
rect 43530 2428 43536 2440
rect 41923 2400 43536 2428
rect 41923 2397 41935 2400
rect 41877 2391 41935 2397
rect 43530 2388 43536 2400
rect 43588 2388 43594 2440
rect 23750 2320 23756 2372
rect 23808 2360 23814 2372
rect 24581 2363 24639 2369
rect 24581 2360 24593 2363
rect 23808 2332 24593 2360
rect 23808 2320 23814 2332
rect 24581 2329 24593 2332
rect 24627 2329 24639 2363
rect 24581 2323 24639 2329
rect 1104 2202 44896 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 44896 2202
rect 1104 2128 44896 2150
<< via1 >>
rect 23848 44072 23900 44124
rect 24860 44072 24912 44124
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 1860 43299 1912 43308
rect 1860 43265 1869 43299
rect 1869 43265 1903 43299
rect 1903 43265 1912 43299
rect 1860 43256 1912 43265
rect 3332 43256 3384 43308
rect 7748 43256 7800 43308
rect 12532 43299 12584 43308
rect 12532 43265 12541 43299
rect 12541 43265 12575 43299
rect 12575 43265 12584 43299
rect 12532 43256 12584 43265
rect 13084 43299 13136 43308
rect 13084 43265 13093 43299
rect 13093 43265 13127 43299
rect 13127 43265 13136 43299
rect 13084 43256 13136 43265
rect 3608 43188 3660 43240
rect 3792 43231 3844 43240
rect 3792 43197 3801 43231
rect 3801 43197 3835 43231
rect 3835 43197 3844 43231
rect 3792 43188 3844 43197
rect 3976 43231 4028 43240
rect 3976 43197 3985 43231
rect 3985 43197 4019 43231
rect 4019 43197 4028 43231
rect 3976 43188 4028 43197
rect 14096 43231 14148 43240
rect 2044 43120 2096 43172
rect 14096 43197 14105 43231
rect 14105 43197 14139 43231
rect 14139 43197 14148 43231
rect 14096 43188 14148 43197
rect 13544 43120 13596 43172
rect 23480 43324 23532 43376
rect 25780 43324 25832 43376
rect 24860 43231 24912 43240
rect 24860 43197 24869 43231
rect 24869 43197 24903 43231
rect 24903 43197 24912 43231
rect 24860 43188 24912 43197
rect 33324 43188 33376 43240
rect 33508 43231 33560 43240
rect 33508 43197 33517 43231
rect 33517 43197 33551 43231
rect 33551 43197 33560 43231
rect 33508 43188 33560 43197
rect 2780 43095 2832 43104
rect 2780 43061 2789 43095
rect 2789 43061 2823 43095
rect 2823 43061 2832 43095
rect 2780 43052 2832 43061
rect 6552 43095 6604 43104
rect 6552 43061 6561 43095
rect 6561 43061 6595 43095
rect 6595 43061 6604 43095
rect 6552 43052 6604 43061
rect 8024 43095 8076 43104
rect 8024 43061 8033 43095
rect 8033 43061 8067 43095
rect 8067 43061 8076 43095
rect 8024 43052 8076 43061
rect 11520 43052 11572 43104
rect 11612 43052 11664 43104
rect 12440 43095 12492 43104
rect 12440 43061 12449 43095
rect 12449 43061 12483 43095
rect 12483 43061 12492 43095
rect 12440 43052 12492 43061
rect 20812 43095 20864 43104
rect 20812 43061 20821 43095
rect 20821 43061 20855 43095
rect 20855 43061 20864 43095
rect 20812 43052 20864 43061
rect 22652 43095 22704 43104
rect 22652 43061 22661 43095
rect 22661 43061 22695 43095
rect 22695 43061 22704 43095
rect 22652 43052 22704 43061
rect 27160 43052 27212 43104
rect 27804 43052 27856 43104
rect 30472 43095 30524 43104
rect 30472 43061 30481 43095
rect 30481 43061 30515 43095
rect 30515 43061 30524 43095
rect 30472 43052 30524 43061
rect 33140 43120 33192 43172
rect 34520 43052 34572 43104
rect 40040 43095 40092 43104
rect 40040 43061 40049 43095
rect 40049 43061 40083 43095
rect 40083 43061 40092 43095
rect 40040 43052 40092 43061
rect 42892 43095 42944 43104
rect 42892 43061 42901 43095
rect 42901 43061 42935 43095
rect 42935 43061 42944 43095
rect 42892 43052 42944 43061
rect 44180 43052 44232 43104
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 13084 42848 13136 42900
rect 22560 42848 22612 42900
rect 24492 42780 24544 42832
rect 40040 42780 40092 42832
rect 2872 42712 2924 42764
rect 10324 42755 10376 42764
rect 10324 42721 10333 42755
rect 10333 42721 10367 42755
rect 10367 42721 10376 42755
rect 10324 42712 10376 42721
rect 11612 42755 11664 42764
rect 11612 42721 11621 42755
rect 11621 42721 11655 42755
rect 11655 42721 11664 42755
rect 11612 42712 11664 42721
rect 12256 42712 12308 42764
rect 14832 42755 14884 42764
rect 14832 42721 14841 42755
rect 14841 42721 14875 42755
rect 14875 42721 14884 42755
rect 14832 42712 14884 42721
rect 20812 42755 20864 42764
rect 20812 42721 20821 42755
rect 20821 42721 20855 42755
rect 20855 42721 20864 42755
rect 20812 42712 20864 42721
rect 21272 42755 21324 42764
rect 21272 42721 21281 42755
rect 21281 42721 21315 42755
rect 21315 42721 21324 42755
rect 21272 42712 21324 42721
rect 27068 42712 27120 42764
rect 30472 42755 30524 42764
rect 30472 42721 30481 42755
rect 30481 42721 30515 42755
rect 30515 42721 30524 42755
rect 30472 42712 30524 42721
rect 30932 42755 30984 42764
rect 30932 42721 30941 42755
rect 30941 42721 30975 42755
rect 30975 42721 30984 42755
rect 30932 42712 30984 42721
rect 33140 42755 33192 42764
rect 33140 42721 33149 42755
rect 33149 42721 33183 42755
rect 33183 42721 33192 42755
rect 33140 42712 33192 42721
rect 37372 42755 37424 42764
rect 37372 42721 37381 42755
rect 37381 42721 37415 42755
rect 37415 42721 37424 42755
rect 37372 42712 37424 42721
rect 41788 42755 41840 42764
rect 41788 42721 41797 42755
rect 41797 42721 41831 42755
rect 41831 42721 41840 42755
rect 41788 42712 41840 42721
rect 42892 42712 42944 42764
rect 43812 42755 43864 42764
rect 43812 42721 43821 42755
rect 43821 42721 43855 42755
rect 43855 42721 43864 42755
rect 43812 42712 43864 42721
rect 3240 42687 3292 42696
rect 3240 42653 3249 42687
rect 3249 42653 3283 42687
rect 3283 42653 3292 42687
rect 3240 42644 3292 42653
rect 4620 42644 4672 42696
rect 7104 42687 7156 42696
rect 7104 42653 7113 42687
rect 7113 42653 7147 42687
rect 7147 42653 7156 42687
rect 7104 42644 7156 42653
rect 9312 42687 9364 42696
rect 9312 42653 9321 42687
rect 9321 42653 9355 42687
rect 9355 42653 9364 42687
rect 9312 42644 9364 42653
rect 14372 42687 14424 42696
rect 14372 42653 14381 42687
rect 14381 42653 14415 42687
rect 14415 42653 14424 42687
rect 14372 42644 14424 42653
rect 15752 42644 15804 42696
rect 26424 42644 26476 42696
rect 33968 42687 34020 42696
rect 33968 42653 33977 42687
rect 33977 42653 34011 42687
rect 34011 42653 34020 42687
rect 33968 42644 34020 42653
rect 35440 42687 35492 42696
rect 35440 42653 35449 42687
rect 35449 42653 35483 42687
rect 35483 42653 35492 42687
rect 35440 42644 35492 42653
rect 6460 42619 6512 42628
rect 6460 42585 6469 42619
rect 6469 42585 6503 42619
rect 6503 42585 6512 42619
rect 6460 42576 6512 42585
rect 10048 42576 10100 42628
rect 11796 42619 11848 42628
rect 11796 42585 11805 42619
rect 11805 42585 11839 42619
rect 11839 42585 11848 42619
rect 11796 42576 11848 42585
rect 14556 42619 14608 42628
rect 14556 42585 14565 42619
rect 14565 42585 14599 42619
rect 14599 42585 14608 42619
rect 14556 42576 14608 42585
rect 20996 42619 21048 42628
rect 20996 42585 21005 42619
rect 21005 42585 21039 42619
rect 21039 42585 21048 42619
rect 20996 42576 21048 42585
rect 24584 42619 24636 42628
rect 24584 42585 24593 42619
rect 24593 42585 24627 42619
rect 24627 42585 24636 42619
rect 24584 42576 24636 42585
rect 27068 42576 27120 42628
rect 30656 42619 30708 42628
rect 30656 42585 30665 42619
rect 30665 42585 30699 42619
rect 30699 42585 30708 42619
rect 30656 42576 30708 42585
rect 37832 42576 37884 42628
rect 39948 42576 40000 42628
rect 42708 42576 42760 42628
rect 3148 42508 3200 42560
rect 12532 42508 12584 42560
rect 33416 42508 33468 42560
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 2596 42304 2648 42356
rect 2780 42236 2832 42288
rect 11796 42304 11848 42356
rect 20996 42304 21048 42356
rect 27068 42347 27120 42356
rect 27068 42313 27077 42347
rect 27077 42313 27111 42347
rect 27111 42313 27120 42347
rect 27068 42304 27120 42313
rect 30656 42347 30708 42356
rect 30656 42313 30665 42347
rect 30665 42313 30699 42347
rect 30699 42313 30708 42347
rect 30656 42304 30708 42313
rect 33324 42347 33376 42356
rect 33324 42313 33333 42347
rect 33333 42313 33367 42347
rect 33367 42313 33376 42347
rect 33324 42304 33376 42313
rect 34152 42304 34204 42356
rect 34888 42304 34940 42356
rect 4988 42168 5040 42220
rect 1860 42143 1912 42152
rect 1860 42109 1869 42143
rect 1869 42109 1903 42143
rect 1903 42109 1912 42143
rect 1860 42100 1912 42109
rect 2872 42143 2924 42152
rect 2872 42109 2881 42143
rect 2881 42109 2915 42143
rect 2915 42109 2924 42143
rect 2872 42100 2924 42109
rect 7104 42100 7156 42152
rect 12440 42236 12492 42288
rect 9312 42168 9364 42220
rect 7472 42032 7524 42084
rect 11520 42168 11572 42220
rect 15752 42236 15804 42288
rect 38660 42304 38712 42356
rect 42708 42347 42760 42356
rect 42708 42313 42717 42347
rect 42717 42313 42751 42347
rect 42751 42313 42760 42347
rect 42708 42304 42760 42313
rect 42616 42236 42668 42288
rect 20812 42211 20864 42220
rect 20812 42177 20821 42211
rect 20821 42177 20855 42211
rect 20855 42177 20864 42211
rect 20812 42168 20864 42177
rect 22652 42211 22704 42220
rect 22652 42177 22661 42211
rect 22661 42177 22695 42211
rect 22695 42177 22704 42211
rect 22652 42168 22704 42177
rect 26424 42211 26476 42220
rect 26424 42177 26433 42211
rect 26433 42177 26467 42211
rect 26467 42177 26476 42211
rect 26424 42168 26476 42177
rect 27804 42211 27856 42220
rect 12900 42143 12952 42152
rect 12900 42109 12909 42143
rect 12909 42109 12943 42143
rect 12943 42109 12952 42143
rect 12900 42100 12952 42109
rect 14464 42143 14516 42152
rect 14464 42109 14473 42143
rect 14473 42109 14507 42143
rect 14507 42109 14516 42143
rect 14464 42100 14516 42109
rect 22836 42143 22888 42152
rect 22836 42109 22845 42143
rect 22845 42109 22879 42143
rect 22879 42109 22888 42143
rect 22836 42100 22888 42109
rect 23204 42143 23256 42152
rect 23204 42109 23213 42143
rect 23213 42109 23247 42143
rect 23247 42109 23256 42143
rect 23204 42100 23256 42109
rect 27804 42177 27813 42211
rect 27813 42177 27847 42211
rect 27847 42177 27856 42211
rect 27804 42168 27856 42177
rect 30564 42211 30616 42220
rect 30564 42177 30573 42211
rect 30573 42177 30607 42211
rect 30607 42177 30616 42211
rect 30564 42168 30616 42177
rect 33416 42211 33468 42220
rect 33416 42177 33425 42211
rect 33425 42177 33459 42211
rect 33459 42177 33468 42211
rect 33416 42168 33468 42177
rect 33968 42211 34020 42220
rect 33968 42177 33977 42211
rect 33977 42177 34011 42211
rect 34011 42177 34020 42211
rect 33968 42168 34020 42177
rect 36452 42211 36504 42220
rect 36452 42177 36461 42211
rect 36461 42177 36495 42211
rect 36495 42177 36504 42211
rect 36452 42168 36504 42177
rect 42800 42211 42852 42220
rect 42800 42177 42809 42211
rect 42809 42177 42843 42211
rect 42843 42177 42852 42211
rect 42800 42168 42852 42177
rect 14004 42032 14056 42084
rect 20812 42032 20864 42084
rect 27068 42032 27120 42084
rect 6368 41964 6420 42016
rect 28080 42100 28132 42152
rect 28356 42143 28408 42152
rect 28356 42109 28365 42143
rect 28365 42109 28399 42143
rect 28399 42109 28408 42143
rect 28356 42100 28408 42109
rect 34796 42100 34848 42152
rect 34888 42143 34940 42152
rect 34888 42109 34897 42143
rect 34897 42109 34931 42143
rect 34931 42109 34940 42143
rect 34888 42100 34940 42109
rect 35348 42032 35400 42084
rect 38384 42100 38436 42152
rect 35624 41964 35676 42016
rect 42800 42032 42852 42084
rect 43536 42168 43588 42220
rect 43904 42211 43956 42220
rect 43904 42177 43913 42211
rect 43913 42177 43947 42211
rect 43947 42177 43956 42211
rect 43904 42168 43956 42177
rect 43352 42007 43404 42016
rect 43352 41973 43361 42007
rect 43361 41973 43395 42007
rect 43395 41973 43404 42007
rect 43352 41964 43404 41973
rect 43996 42007 44048 42016
rect 43996 41973 44005 42007
rect 44005 41973 44039 42007
rect 44039 41973 44048 42007
rect 43996 41964 44048 41973
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 3976 41760 4028 41812
rect 4988 41760 5040 41812
rect 10048 41803 10100 41812
rect 2964 41692 3016 41744
rect 10048 41769 10057 41803
rect 10057 41769 10091 41803
rect 10091 41769 10100 41803
rect 10048 41760 10100 41769
rect 14556 41803 14608 41812
rect 14556 41769 14565 41803
rect 14565 41769 14599 41803
rect 14599 41769 14608 41803
rect 14556 41760 14608 41769
rect 22836 41760 22888 41812
rect 23480 41760 23532 41812
rect 24584 41760 24636 41812
rect 28080 41803 28132 41812
rect 28080 41769 28089 41803
rect 28089 41769 28123 41803
rect 28123 41769 28132 41803
rect 28080 41760 28132 41769
rect 34796 41803 34848 41812
rect 34796 41769 34805 41803
rect 34805 41769 34839 41803
rect 34839 41769 34848 41803
rect 34796 41760 34848 41769
rect 37832 41803 37884 41812
rect 37832 41769 37841 41803
rect 37841 41769 37875 41803
rect 37875 41769 37884 41803
rect 37832 41760 37884 41769
rect 38384 41803 38436 41812
rect 38384 41769 38393 41803
rect 38393 41769 38427 41803
rect 38427 41769 38436 41803
rect 38384 41760 38436 41769
rect 39948 41803 40000 41812
rect 39948 41769 39957 41803
rect 39957 41769 39991 41803
rect 39991 41769 40000 41803
rect 39948 41760 40000 41769
rect 12164 41692 12216 41744
rect 14372 41692 14424 41744
rect 30564 41692 30616 41744
rect 42892 41692 42944 41744
rect 43904 41692 43956 41744
rect 2872 41624 2924 41676
rect 5172 41667 5224 41676
rect 5172 41633 5181 41667
rect 5181 41633 5215 41667
rect 5215 41633 5224 41667
rect 5172 41624 5224 41633
rect 6368 41667 6420 41676
rect 6368 41633 6377 41667
rect 6377 41633 6411 41667
rect 6411 41633 6420 41667
rect 6368 41624 6420 41633
rect 6552 41667 6604 41676
rect 6552 41633 6561 41667
rect 6561 41633 6595 41667
rect 6595 41633 6604 41667
rect 6552 41624 6604 41633
rect 27068 41624 27120 41676
rect 35256 41624 35308 41676
rect 35440 41667 35492 41676
rect 35440 41633 35449 41667
rect 35449 41633 35483 41667
rect 35483 41633 35492 41667
rect 35440 41624 35492 41633
rect 35624 41667 35676 41676
rect 35624 41633 35633 41667
rect 35633 41633 35667 41667
rect 35667 41633 35676 41667
rect 35624 41624 35676 41633
rect 36084 41667 36136 41676
rect 36084 41633 36093 41667
rect 36093 41633 36127 41667
rect 36127 41633 36136 41667
rect 36084 41624 36136 41633
rect 42524 41667 42576 41676
rect 42524 41633 42533 41667
rect 42533 41633 42567 41667
rect 42567 41633 42576 41667
rect 42524 41624 42576 41633
rect 43996 41667 44048 41676
rect 43996 41633 44005 41667
rect 44005 41633 44039 41667
rect 44039 41633 44048 41667
rect 43996 41624 44048 41633
rect 44180 41667 44232 41676
rect 44180 41633 44189 41667
rect 44189 41633 44223 41667
rect 44223 41633 44232 41667
rect 44180 41624 44232 41633
rect 4620 41556 4672 41608
rect 12072 41599 12124 41608
rect 3056 41531 3108 41540
rect 3056 41497 3065 41531
rect 3065 41497 3099 41531
rect 3099 41497 3108 41531
rect 3056 41488 3108 41497
rect 12072 41565 12081 41599
rect 12081 41565 12115 41599
rect 12115 41565 12124 41599
rect 12072 41556 12124 41565
rect 14648 41556 14700 41608
rect 22560 41556 22612 41608
rect 22836 41556 22888 41608
rect 24400 41599 24452 41608
rect 24400 41565 24409 41599
rect 24409 41565 24443 41599
rect 24443 41565 24452 41599
rect 24400 41556 24452 41565
rect 28172 41599 28224 41608
rect 10968 41531 11020 41540
rect 10968 41497 10977 41531
rect 10977 41497 11011 41531
rect 11011 41497 11020 41531
rect 10968 41488 11020 41497
rect 12992 41488 13044 41540
rect 28172 41565 28181 41599
rect 28181 41565 28215 41599
rect 28215 41565 28224 41599
rect 28172 41556 28224 41565
rect 34520 41556 34572 41608
rect 37924 41599 37976 41608
rect 37924 41565 37933 41599
rect 37933 41565 37967 41599
rect 37967 41565 37976 41599
rect 37924 41556 37976 41565
rect 39856 41599 39908 41608
rect 39856 41565 39865 41599
rect 39865 41565 39899 41599
rect 39899 41565 39908 41599
rect 39856 41556 39908 41565
rect 43260 41420 43312 41472
rect 44456 41420 44508 41472
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 3056 41216 3108 41268
rect 6460 41259 6512 41268
rect 6460 41225 6469 41259
rect 6469 41225 6503 41259
rect 6503 41225 6512 41259
rect 6460 41216 6512 41225
rect 3148 41148 3200 41200
rect 12532 41216 12584 41268
rect 14464 41216 14516 41268
rect 1860 41080 1912 41132
rect 2320 41012 2372 41064
rect 3240 41080 3292 41132
rect 5632 41080 5684 41132
rect 9312 41148 9364 41200
rect 39856 41216 39908 41268
rect 10692 41123 10744 41132
rect 10692 41089 10701 41123
rect 10701 41089 10735 41123
rect 10735 41089 10744 41123
rect 10692 41080 10744 41089
rect 11060 41080 11112 41132
rect 12072 41080 12124 41132
rect 14004 41080 14056 41132
rect 14648 41080 14700 41132
rect 32496 41123 32548 41132
rect 32496 41089 32505 41123
rect 32505 41089 32539 41123
rect 32539 41089 32548 41123
rect 32496 41080 32548 41089
rect 32588 41123 32640 41132
rect 32588 41089 32597 41123
rect 32597 41089 32631 41123
rect 32631 41089 32640 41123
rect 32588 41080 32640 41089
rect 33048 41080 33100 41132
rect 33416 41123 33468 41132
rect 33416 41089 33425 41123
rect 33425 41089 33459 41123
rect 33459 41089 33468 41123
rect 33416 41080 33468 41089
rect 4712 41055 4764 41064
rect 4712 41021 4721 41055
rect 4721 41021 4755 41055
rect 4755 41021 4764 41055
rect 4712 41012 4764 41021
rect 6644 41012 6696 41064
rect 9588 41055 9640 41064
rect 4804 40944 4856 40996
rect 9588 41021 9597 41055
rect 9597 41021 9631 41055
rect 9631 41021 9640 41055
rect 9588 41012 9640 41021
rect 36452 41012 36504 41064
rect 41512 41012 41564 41064
rect 43444 41012 43496 41064
rect 11060 40944 11112 40996
rect 9588 40876 9640 40928
rect 30564 40944 30616 40996
rect 13268 40876 13320 40928
rect 22836 40876 22888 40928
rect 23388 40876 23440 40928
rect 33324 40876 33376 40928
rect 33600 40919 33652 40928
rect 33600 40885 33609 40919
rect 33609 40885 33643 40919
rect 33643 40885 33652 40919
rect 33600 40876 33652 40885
rect 44180 40919 44232 40928
rect 44180 40885 44189 40919
rect 44189 40885 44223 40919
rect 44223 40885 44232 40919
rect 44180 40876 44232 40885
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 2872 40715 2924 40724
rect 2872 40681 2881 40715
rect 2881 40681 2915 40715
rect 2915 40681 2924 40715
rect 2872 40672 2924 40681
rect 14096 40672 14148 40724
rect 32312 40715 32364 40724
rect 32312 40681 32321 40715
rect 32321 40681 32355 40715
rect 32355 40681 32364 40715
rect 32312 40672 32364 40681
rect 32496 40672 32548 40724
rect 2320 40604 2372 40656
rect 10692 40536 10744 40588
rect 37372 40604 37424 40656
rect 40684 40604 40736 40656
rect 28908 40536 28960 40588
rect 43260 40579 43312 40588
rect 43260 40545 43269 40579
rect 43269 40545 43303 40579
rect 43303 40545 43312 40579
rect 43260 40536 43312 40545
rect 43352 40536 43404 40588
rect 44180 40579 44232 40588
rect 44180 40545 44189 40579
rect 44189 40545 44223 40579
rect 44223 40545 44232 40579
rect 44180 40536 44232 40545
rect 1952 40468 2004 40520
rect 3608 40468 3660 40520
rect 3884 40511 3936 40520
rect 3884 40477 3893 40511
rect 3893 40477 3927 40511
rect 3927 40477 3936 40511
rect 3884 40468 3936 40477
rect 5632 40468 5684 40520
rect 8852 40468 8904 40520
rect 9312 40511 9364 40520
rect 9312 40477 9321 40511
rect 9321 40477 9355 40511
rect 9355 40477 9364 40511
rect 9312 40468 9364 40477
rect 7472 40443 7524 40452
rect 7472 40409 7481 40443
rect 7481 40409 7515 40443
rect 7515 40409 7524 40443
rect 7472 40400 7524 40409
rect 10140 40443 10192 40452
rect 10140 40409 10149 40443
rect 10149 40409 10183 40443
rect 10183 40409 10192 40443
rect 12072 40468 12124 40520
rect 31116 40511 31168 40520
rect 10140 40400 10192 40409
rect 5908 40375 5960 40384
rect 5908 40341 5917 40375
rect 5917 40341 5951 40375
rect 5951 40341 5960 40375
rect 5908 40332 5960 40341
rect 14648 40400 14700 40452
rect 26424 40400 26476 40452
rect 31116 40477 31125 40511
rect 31125 40477 31159 40511
rect 31159 40477 31168 40511
rect 31116 40468 31168 40477
rect 32128 40511 32180 40520
rect 32128 40477 32137 40511
rect 32137 40477 32171 40511
rect 32171 40477 32180 40511
rect 32128 40468 32180 40477
rect 30748 40400 30800 40452
rect 35348 40468 35400 40520
rect 37740 40468 37792 40520
rect 39948 40468 40000 40520
rect 40040 40511 40092 40520
rect 40040 40477 40049 40511
rect 40049 40477 40083 40511
rect 40083 40477 40092 40511
rect 40500 40511 40552 40520
rect 40040 40468 40092 40477
rect 40500 40477 40509 40511
rect 40509 40477 40543 40511
rect 40543 40477 40552 40511
rect 40500 40468 40552 40477
rect 33600 40400 33652 40452
rect 37280 40443 37332 40452
rect 37280 40409 37289 40443
rect 37289 40409 37323 40443
rect 37323 40409 37332 40443
rect 37280 40400 37332 40409
rect 40776 40443 40828 40452
rect 20812 40332 20864 40384
rect 28080 40332 28132 40384
rect 31024 40332 31076 40384
rect 33048 40332 33100 40384
rect 35256 40375 35308 40384
rect 35256 40341 35265 40375
rect 35265 40341 35299 40375
rect 35299 40341 35308 40375
rect 35256 40332 35308 40341
rect 37648 40332 37700 40384
rect 39212 40332 39264 40384
rect 40776 40409 40785 40443
rect 40785 40409 40819 40443
rect 40819 40409 40828 40443
rect 40776 40400 40828 40409
rect 40592 40375 40644 40384
rect 40592 40341 40601 40375
rect 40601 40341 40635 40375
rect 40635 40341 40644 40375
rect 40592 40332 40644 40341
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 4620 40128 4672 40180
rect 13084 40128 13136 40180
rect 27436 40128 27488 40180
rect 31116 40171 31168 40180
rect 31116 40137 31125 40171
rect 31125 40137 31159 40171
rect 31159 40137 31168 40171
rect 31116 40128 31168 40137
rect 2872 40060 2924 40112
rect 1952 40035 2004 40044
rect 1952 40001 1961 40035
rect 1961 40001 1995 40035
rect 1995 40001 2004 40035
rect 1952 39992 2004 40001
rect 5632 40060 5684 40112
rect 12072 40060 12124 40112
rect 29828 40103 29880 40112
rect 29828 40069 29837 40103
rect 29837 40069 29871 40103
rect 29871 40069 29880 40103
rect 29828 40060 29880 40069
rect 31300 40060 31352 40112
rect 32588 40128 32640 40180
rect 33416 40128 33468 40180
rect 37648 40128 37700 40180
rect 33048 40060 33100 40112
rect 34520 40060 34572 40112
rect 35256 40060 35308 40112
rect 39488 40103 39540 40112
rect 39488 40069 39497 40103
rect 39497 40069 39531 40103
rect 39531 40069 39540 40103
rect 39488 40060 39540 40069
rect 40684 40060 40736 40112
rect 19248 39992 19300 40044
rect 20536 40035 20588 40044
rect 20536 40001 20545 40035
rect 20545 40001 20579 40035
rect 20579 40001 20588 40035
rect 20536 39992 20588 40001
rect 24584 39992 24636 40044
rect 27068 39992 27120 40044
rect 30288 39992 30340 40044
rect 37372 39992 37424 40044
rect 2780 39967 2832 39976
rect 2780 39933 2789 39967
rect 2789 39933 2823 39967
rect 2823 39933 2832 39967
rect 2780 39924 2832 39933
rect 4620 39924 4672 39976
rect 12164 39967 12216 39976
rect 12164 39933 12173 39967
rect 12173 39933 12207 39967
rect 12207 39933 12216 39967
rect 12164 39924 12216 39933
rect 16396 39924 16448 39976
rect 18696 39967 18748 39976
rect 18696 39933 18705 39967
rect 18705 39933 18739 39967
rect 18739 39933 18748 39967
rect 18696 39924 18748 39933
rect 26976 39967 27028 39976
rect 19984 39788 20036 39840
rect 20720 39831 20772 39840
rect 20720 39797 20729 39831
rect 20729 39797 20763 39831
rect 20763 39797 20772 39831
rect 20720 39788 20772 39797
rect 26976 39933 26985 39967
rect 26985 39933 27019 39967
rect 27019 39933 27028 39967
rect 26976 39924 27028 39933
rect 31760 39924 31812 39976
rect 32312 39924 32364 39976
rect 36084 39924 36136 39976
rect 24308 39788 24360 39840
rect 31484 39856 31536 39908
rect 32956 39899 33008 39908
rect 32956 39865 32965 39899
rect 32965 39865 32999 39899
rect 32999 39865 33008 39899
rect 32956 39856 33008 39865
rect 25320 39788 25372 39840
rect 30012 39831 30064 39840
rect 30012 39797 30021 39831
rect 30021 39797 30055 39831
rect 30055 39797 30064 39831
rect 30012 39788 30064 39797
rect 30104 39788 30156 39840
rect 32312 39831 32364 39840
rect 32312 39797 32321 39831
rect 32321 39797 32355 39831
rect 32355 39797 32364 39831
rect 32312 39788 32364 39797
rect 33324 39831 33376 39840
rect 33324 39797 33333 39831
rect 33333 39797 33367 39831
rect 33367 39797 33376 39831
rect 33324 39788 33376 39797
rect 33968 39788 34020 39840
rect 39948 39924 40000 39976
rect 38936 39856 38988 39908
rect 40040 39856 40092 39908
rect 39396 39788 39448 39840
rect 41880 39831 41932 39840
rect 41880 39797 41889 39831
rect 41889 39797 41923 39831
rect 41923 39797 41932 39831
rect 41880 39788 41932 39797
rect 44180 39788 44232 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 2872 39627 2924 39636
rect 2872 39593 2881 39627
rect 2881 39593 2915 39627
rect 2915 39593 2924 39627
rect 2872 39584 2924 39593
rect 3792 39627 3844 39636
rect 3792 39593 3801 39627
rect 3801 39593 3835 39627
rect 3835 39593 3844 39627
rect 3792 39584 3844 39593
rect 19248 39627 19300 39636
rect 19248 39593 19257 39627
rect 19257 39593 19291 39627
rect 19291 39593 19300 39627
rect 19248 39584 19300 39593
rect 24584 39627 24636 39636
rect 24584 39593 24593 39627
rect 24593 39593 24627 39627
rect 24627 39593 24636 39627
rect 24584 39584 24636 39593
rect 27068 39627 27120 39636
rect 27068 39593 27077 39627
rect 27077 39593 27111 39627
rect 27111 39593 27120 39627
rect 27068 39584 27120 39593
rect 28908 39627 28960 39636
rect 28908 39593 28917 39627
rect 28917 39593 28951 39627
rect 28951 39593 28960 39627
rect 28908 39584 28960 39593
rect 32128 39627 32180 39636
rect 32128 39593 32137 39627
rect 32137 39593 32171 39627
rect 32171 39593 32180 39627
rect 32128 39584 32180 39593
rect 35348 39584 35400 39636
rect 37280 39584 37332 39636
rect 38936 39627 38988 39636
rect 38936 39593 38945 39627
rect 38945 39593 38979 39627
rect 38979 39593 38988 39627
rect 38936 39584 38988 39593
rect 39212 39584 39264 39636
rect 39488 39584 39540 39636
rect 40776 39584 40828 39636
rect 32588 39516 32640 39568
rect 34520 39516 34572 39568
rect 39396 39516 39448 39568
rect 10140 39448 10192 39500
rect 18696 39448 18748 39500
rect 26424 39491 26476 39500
rect 4804 39423 4856 39432
rect 4804 39389 4813 39423
rect 4813 39389 4847 39423
rect 4847 39389 4856 39423
rect 4804 39380 4856 39389
rect 5632 39423 5684 39432
rect 5632 39389 5641 39423
rect 5641 39389 5675 39423
rect 5675 39389 5684 39423
rect 5632 39380 5684 39389
rect 19984 39380 20036 39432
rect 26424 39457 26433 39491
rect 26433 39457 26467 39491
rect 26467 39457 26476 39491
rect 26424 39448 26476 39457
rect 27436 39448 27488 39500
rect 30748 39491 30800 39500
rect 30748 39457 30757 39491
rect 30757 39457 30791 39491
rect 30791 39457 30800 39491
rect 30748 39448 30800 39457
rect 21640 39380 21692 39432
rect 22928 39380 22980 39432
rect 25504 39423 25556 39432
rect 25504 39389 25513 39423
rect 25513 39389 25547 39423
rect 25547 39389 25556 39423
rect 25504 39380 25556 39389
rect 25596 39423 25648 39432
rect 25596 39389 25605 39423
rect 25605 39389 25639 39423
rect 25639 39389 25648 39423
rect 25596 39380 25648 39389
rect 26884 39423 26936 39432
rect 20444 39312 20496 39364
rect 20720 39355 20772 39364
rect 20720 39321 20754 39355
rect 20754 39321 20772 39355
rect 20720 39312 20772 39321
rect 24492 39355 24544 39364
rect 24492 39321 24501 39355
rect 24501 39321 24535 39355
rect 24535 39321 24544 39355
rect 24492 39312 24544 39321
rect 25412 39312 25464 39364
rect 26884 39389 26893 39423
rect 26893 39389 26927 39423
rect 26927 39389 26936 39423
rect 26884 39380 26936 39389
rect 26976 39380 27028 39432
rect 29460 39380 29512 39432
rect 30288 39423 30340 39432
rect 30288 39389 30297 39423
rect 30297 39389 30331 39423
rect 30331 39389 30340 39423
rect 30288 39380 30340 39389
rect 31024 39423 31076 39432
rect 31024 39389 31058 39423
rect 31058 39389 31076 39423
rect 31024 39380 31076 39389
rect 31484 39380 31536 39432
rect 32128 39380 32180 39432
rect 32956 39380 33008 39432
rect 33968 39423 34020 39432
rect 33968 39389 33977 39423
rect 33977 39389 34011 39423
rect 34011 39389 34020 39423
rect 33968 39380 34020 39389
rect 34704 39423 34756 39432
rect 34704 39389 34713 39423
rect 34713 39389 34747 39423
rect 34747 39389 34756 39423
rect 34704 39380 34756 39389
rect 27896 39312 27948 39364
rect 30840 39312 30892 39364
rect 20076 39244 20128 39296
rect 20812 39244 20864 39296
rect 30012 39244 30064 39296
rect 31852 39244 31904 39296
rect 33324 39312 33376 39364
rect 33048 39287 33100 39296
rect 33048 39253 33057 39287
rect 33057 39253 33091 39287
rect 33091 39253 33100 39287
rect 33232 39287 33284 39296
rect 33048 39244 33100 39253
rect 33232 39253 33241 39287
rect 33241 39253 33275 39287
rect 33275 39253 33284 39287
rect 33232 39244 33284 39253
rect 34520 39244 34572 39296
rect 37740 39448 37792 39500
rect 40776 39491 40828 39500
rect 37648 39380 37700 39432
rect 39212 39380 39264 39432
rect 39672 39380 39724 39432
rect 40776 39457 40785 39491
rect 40785 39457 40819 39491
rect 40819 39457 40828 39491
rect 40776 39448 40828 39457
rect 40500 39380 40552 39432
rect 41052 39516 41104 39568
rect 42708 39491 42760 39500
rect 42708 39457 42717 39491
rect 42717 39457 42751 39491
rect 42751 39457 42760 39491
rect 42708 39448 42760 39457
rect 44180 39491 44232 39500
rect 44180 39457 44189 39491
rect 44189 39457 44223 39491
rect 44223 39457 44232 39491
rect 44180 39448 44232 39457
rect 39304 39355 39356 39364
rect 39304 39321 39313 39355
rect 39313 39321 39347 39355
rect 39347 39321 39356 39355
rect 39304 39312 39356 39321
rect 40592 39312 40644 39364
rect 41880 39380 41932 39432
rect 37556 39244 37608 39296
rect 40776 39244 40828 39296
rect 43444 39312 43496 39364
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 20536 39040 20588 39092
rect 24492 39040 24544 39092
rect 26884 39040 26936 39092
rect 27896 39083 27948 39092
rect 27896 39049 27905 39083
rect 27905 39049 27939 39083
rect 27939 39049 27948 39083
rect 27896 39040 27948 39049
rect 30840 39083 30892 39092
rect 30840 39049 30849 39083
rect 30849 39049 30883 39083
rect 30883 39049 30892 39083
rect 30840 39040 30892 39049
rect 31300 39083 31352 39092
rect 31300 39049 31309 39083
rect 31309 39049 31343 39083
rect 31343 39049 31352 39083
rect 31300 39040 31352 39049
rect 43444 39083 43496 39092
rect 16764 38836 16816 38888
rect 16948 38947 17000 38956
rect 16948 38913 16957 38947
rect 16957 38913 16991 38947
rect 16991 38913 17000 38947
rect 16948 38904 17000 38913
rect 18420 38904 18472 38956
rect 25412 38972 25464 39024
rect 25596 38972 25648 39024
rect 28172 38972 28224 39024
rect 20076 38904 20128 38956
rect 22192 38947 22244 38956
rect 22192 38913 22226 38947
rect 22226 38913 22244 38947
rect 24400 38947 24452 38956
rect 22192 38904 22244 38913
rect 24400 38913 24409 38947
rect 24409 38913 24443 38947
rect 24443 38913 24452 38947
rect 24400 38904 24452 38913
rect 25320 38947 25372 38956
rect 25320 38913 25329 38947
rect 25329 38913 25363 38947
rect 25363 38913 25372 38947
rect 25320 38904 25372 38913
rect 25872 38904 25924 38956
rect 27160 38947 27212 38956
rect 27160 38913 27169 38947
rect 27169 38913 27203 38947
rect 27203 38913 27212 38947
rect 27160 38904 27212 38913
rect 28080 38947 28132 38956
rect 28080 38913 28089 38947
rect 28089 38913 28123 38947
rect 28123 38913 28132 38947
rect 28080 38904 28132 38913
rect 29460 38947 29512 38956
rect 29460 38913 29469 38947
rect 29469 38913 29503 38947
rect 29503 38913 29512 38947
rect 29460 38904 29512 38913
rect 29736 38947 29788 38956
rect 29736 38913 29770 38947
rect 29770 38913 29788 38947
rect 29736 38904 29788 38913
rect 16856 38743 16908 38752
rect 16856 38709 16865 38743
rect 16865 38709 16899 38743
rect 16899 38709 16908 38743
rect 16856 38700 16908 38709
rect 19340 38700 19392 38752
rect 20812 38836 20864 38888
rect 21640 38836 21692 38888
rect 27436 38879 27488 38888
rect 27436 38845 27445 38879
rect 27445 38845 27479 38879
rect 27479 38845 27488 38879
rect 27436 38836 27488 38845
rect 32588 38972 32640 39024
rect 33416 38972 33468 39024
rect 31760 38904 31812 38956
rect 31852 38904 31904 38956
rect 33324 38947 33376 38956
rect 33324 38913 33333 38947
rect 33333 38913 33367 38947
rect 33367 38913 33376 38947
rect 33324 38904 33376 38913
rect 34060 38947 34112 38956
rect 34060 38913 34069 38947
rect 34069 38913 34103 38947
rect 34103 38913 34112 38947
rect 34060 38904 34112 38913
rect 37280 38904 37332 38956
rect 37372 38904 37424 38956
rect 37648 38947 37700 38956
rect 37648 38913 37657 38947
rect 37657 38913 37691 38947
rect 37691 38913 37700 38947
rect 37648 38904 37700 38913
rect 37740 38947 37792 38956
rect 37740 38913 37749 38947
rect 37749 38913 37783 38947
rect 37783 38913 37792 38947
rect 38844 38947 38896 38956
rect 37740 38904 37792 38913
rect 38844 38913 38853 38947
rect 38853 38913 38887 38947
rect 38887 38913 38896 38947
rect 38844 38904 38896 38913
rect 38936 38947 38988 38956
rect 38936 38913 38945 38947
rect 38945 38913 38979 38947
rect 38979 38913 38988 38947
rect 38936 38904 38988 38913
rect 39304 38904 39356 38956
rect 39672 38904 39724 38956
rect 43444 39049 43453 39083
rect 43453 39049 43487 39083
rect 43487 39049 43496 39083
rect 43444 39040 43496 39049
rect 39120 38879 39172 38888
rect 39120 38845 39129 38879
rect 39129 38845 39163 38879
rect 39163 38845 39172 38879
rect 39120 38836 39172 38845
rect 43168 38904 43220 38956
rect 40776 38879 40828 38888
rect 40776 38845 40785 38879
rect 40785 38845 40819 38879
rect 40819 38845 40828 38879
rect 40776 38836 40828 38845
rect 41052 38879 41104 38888
rect 41052 38845 41061 38879
rect 41061 38845 41095 38879
rect 41095 38845 41104 38879
rect 41052 38836 41104 38845
rect 27804 38768 27856 38820
rect 37740 38768 37792 38820
rect 40040 38768 40092 38820
rect 22928 38700 22980 38752
rect 25044 38700 25096 38752
rect 33048 38743 33100 38752
rect 33048 38709 33057 38743
rect 33057 38709 33091 38743
rect 33091 38709 33100 38743
rect 33048 38700 33100 38709
rect 33508 38743 33560 38752
rect 33508 38709 33517 38743
rect 33517 38709 33551 38743
rect 33551 38709 33560 38743
rect 33508 38700 33560 38709
rect 34152 38700 34204 38752
rect 36360 38700 36412 38752
rect 37464 38700 37516 38752
rect 39856 38700 39908 38752
rect 44180 38743 44232 38752
rect 44180 38709 44189 38743
rect 44189 38709 44223 38743
rect 44223 38709 44232 38743
rect 44180 38700 44232 38709
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 19340 38539 19392 38548
rect 19340 38505 19349 38539
rect 19349 38505 19383 38539
rect 19383 38505 19392 38539
rect 19340 38496 19392 38505
rect 22192 38539 22244 38548
rect 22192 38505 22201 38539
rect 22201 38505 22235 38539
rect 22235 38505 22244 38539
rect 22192 38496 22244 38505
rect 29736 38496 29788 38548
rect 34980 38471 35032 38480
rect 34980 38437 34989 38471
rect 34989 38437 35023 38471
rect 35023 38437 35032 38471
rect 34980 38428 35032 38437
rect 20260 38360 20312 38412
rect 21640 38403 21692 38412
rect 21640 38369 21649 38403
rect 21649 38369 21683 38403
rect 21683 38369 21692 38403
rect 21640 38360 21692 38369
rect 25320 38360 25372 38412
rect 15844 38292 15896 38344
rect 16396 38292 16448 38344
rect 16856 38292 16908 38344
rect 19432 38224 19484 38276
rect 20076 38292 20128 38344
rect 21548 38292 21600 38344
rect 20352 38224 20404 38276
rect 21272 38224 21324 38276
rect 23020 38292 23072 38344
rect 25872 38335 25924 38344
rect 24768 38224 24820 38276
rect 25872 38301 25881 38335
rect 25881 38301 25915 38335
rect 25915 38301 25924 38335
rect 25872 38292 25924 38301
rect 33232 38360 33284 38412
rect 36084 38403 36136 38412
rect 36084 38369 36093 38403
rect 36093 38369 36127 38403
rect 36127 38369 36136 38403
rect 36084 38360 36136 38369
rect 37648 38360 37700 38412
rect 38660 38360 38712 38412
rect 38844 38360 38896 38412
rect 39948 38360 40000 38412
rect 42708 38403 42760 38412
rect 42708 38369 42717 38403
rect 42717 38369 42751 38403
rect 42751 38369 42760 38403
rect 42708 38360 42760 38369
rect 44180 38403 44232 38412
rect 44180 38369 44189 38403
rect 44189 38369 44223 38403
rect 44223 38369 44232 38403
rect 44180 38360 44232 38369
rect 30104 38335 30156 38344
rect 30104 38301 30113 38335
rect 30113 38301 30147 38335
rect 30147 38301 30156 38335
rect 30104 38292 30156 38301
rect 34704 38335 34756 38344
rect 34704 38301 34713 38335
rect 34713 38301 34747 38335
rect 34747 38301 34756 38335
rect 34704 38292 34756 38301
rect 34796 38292 34848 38344
rect 36360 38335 36412 38344
rect 36360 38301 36394 38335
rect 36394 38301 36412 38335
rect 36360 38292 36412 38301
rect 26240 38224 26292 38276
rect 17316 38156 17368 38208
rect 20260 38199 20312 38208
rect 20260 38165 20269 38199
rect 20269 38165 20303 38199
rect 20303 38165 20312 38199
rect 20260 38156 20312 38165
rect 22928 38156 22980 38208
rect 24952 38156 25004 38208
rect 25504 38156 25556 38208
rect 26148 38156 26200 38208
rect 27160 38224 27212 38276
rect 27988 38156 28040 38208
rect 28816 38156 28868 38208
rect 34152 38156 34204 38208
rect 37372 38156 37424 38208
rect 39856 38335 39908 38344
rect 39856 38301 39865 38335
rect 39865 38301 39899 38335
rect 39899 38301 39908 38335
rect 39856 38292 39908 38301
rect 40040 38335 40092 38344
rect 40040 38301 40049 38335
rect 40049 38301 40083 38335
rect 40083 38301 40092 38335
rect 40040 38292 40092 38301
rect 39672 38224 39724 38276
rect 41144 38224 41196 38276
rect 43628 38224 43680 38276
rect 38844 38199 38896 38208
rect 38844 38165 38853 38199
rect 38853 38165 38887 38199
rect 38887 38165 38896 38199
rect 38844 38156 38896 38165
rect 39580 38156 39632 38208
rect 41604 38156 41656 38208
rect 42432 38156 42484 38208
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 16948 37952 17000 38004
rect 18420 37995 18472 38004
rect 18420 37961 18429 37995
rect 18429 37961 18463 37995
rect 18463 37961 18472 37995
rect 18420 37952 18472 37961
rect 19340 37952 19392 38004
rect 20444 37952 20496 38004
rect 21272 37995 21324 38004
rect 21272 37961 21281 37995
rect 21281 37961 21315 37995
rect 21315 37961 21324 37995
rect 21272 37952 21324 37961
rect 33232 37952 33284 38004
rect 34060 37952 34112 38004
rect 37280 37995 37332 38004
rect 37280 37961 37289 37995
rect 37289 37961 37323 37995
rect 37323 37961 37332 37995
rect 37280 37952 37332 37961
rect 4804 37884 4856 37936
rect 17592 37816 17644 37868
rect 18604 37859 18656 37868
rect 18604 37825 18613 37859
rect 18613 37825 18647 37859
rect 18647 37825 18656 37859
rect 18604 37816 18656 37825
rect 17316 37791 17368 37800
rect 17316 37757 17325 37791
rect 17325 37757 17359 37791
rect 17359 37757 17368 37791
rect 17316 37748 17368 37757
rect 18880 37859 18932 37868
rect 18880 37825 18889 37859
rect 18889 37825 18923 37859
rect 18923 37825 18932 37859
rect 18880 37816 18932 37825
rect 19340 37791 19392 37800
rect 19340 37757 19349 37791
rect 19349 37757 19383 37791
rect 19383 37757 19392 37791
rect 19340 37748 19392 37757
rect 19524 37859 19576 37868
rect 19524 37825 19533 37859
rect 19533 37825 19567 37859
rect 19567 37825 19576 37859
rect 19524 37816 19576 37825
rect 20260 37791 20312 37800
rect 20260 37757 20269 37791
rect 20269 37757 20303 37791
rect 20303 37757 20312 37791
rect 20260 37748 20312 37757
rect 19432 37680 19484 37732
rect 21640 37816 21692 37868
rect 23204 37859 23256 37868
rect 23204 37825 23238 37859
rect 23238 37825 23256 37859
rect 23204 37816 23256 37825
rect 25504 37816 25556 37868
rect 26240 37816 26292 37868
rect 27804 37816 27856 37868
rect 32036 37816 32088 37868
rect 21456 37748 21508 37800
rect 24400 37748 24452 37800
rect 24676 37748 24728 37800
rect 27712 37748 27764 37800
rect 28908 37748 28960 37800
rect 32220 37859 32272 37868
rect 32220 37825 32229 37859
rect 32229 37825 32263 37859
rect 32263 37825 32272 37859
rect 32404 37859 32456 37868
rect 32220 37816 32272 37825
rect 32404 37825 32413 37859
rect 32413 37825 32447 37859
rect 32447 37825 32456 37859
rect 32404 37816 32456 37825
rect 33416 37816 33468 37868
rect 33600 37859 33652 37868
rect 33600 37825 33609 37859
rect 33609 37825 33643 37859
rect 33643 37825 33652 37859
rect 33600 37816 33652 37825
rect 34060 37816 34112 37868
rect 34980 37816 35032 37868
rect 37280 37816 37332 37868
rect 32496 37748 32548 37800
rect 36084 37748 36136 37800
rect 27436 37723 27488 37732
rect 27436 37689 27445 37723
rect 27445 37689 27479 37723
rect 27479 37689 27488 37723
rect 27436 37680 27488 37689
rect 32680 37680 32732 37732
rect 38660 37952 38712 38004
rect 41144 37995 41196 38004
rect 41144 37961 41153 37995
rect 41153 37961 41187 37995
rect 41187 37961 41196 37995
rect 41144 37952 41196 37961
rect 39580 37927 39632 37936
rect 39580 37893 39598 37927
rect 39598 37893 39632 37927
rect 39580 37884 39632 37893
rect 39948 37816 40000 37868
rect 41052 37859 41104 37868
rect 41052 37825 41061 37859
rect 41061 37825 41095 37859
rect 41095 37825 41104 37859
rect 41052 37816 41104 37825
rect 43628 37995 43680 38004
rect 43628 37961 43637 37995
rect 43637 37961 43671 37995
rect 43671 37961 43680 37995
rect 43628 37952 43680 37961
rect 43260 37884 43312 37936
rect 42432 37859 42484 37868
rect 42432 37825 42441 37859
rect 42441 37825 42475 37859
rect 42475 37825 42484 37859
rect 42432 37816 42484 37825
rect 43720 37816 43772 37868
rect 3240 37612 3292 37664
rect 17132 37655 17184 37664
rect 17132 37621 17141 37655
rect 17141 37621 17175 37655
rect 17175 37621 17184 37655
rect 17132 37612 17184 37621
rect 19524 37612 19576 37664
rect 20260 37612 20312 37664
rect 24860 37655 24912 37664
rect 24860 37621 24869 37655
rect 24869 37621 24903 37655
rect 24903 37621 24912 37655
rect 24860 37612 24912 37621
rect 25044 37612 25096 37664
rect 26332 37612 26384 37664
rect 27528 37612 27580 37664
rect 31300 37655 31352 37664
rect 31300 37621 31309 37655
rect 31309 37621 31343 37655
rect 31343 37621 31352 37655
rect 31300 37612 31352 37621
rect 32588 37655 32640 37664
rect 32588 37621 32597 37655
rect 32597 37621 32631 37655
rect 32631 37621 32640 37655
rect 32588 37612 32640 37621
rect 33048 37612 33100 37664
rect 42708 37791 42760 37800
rect 42708 37757 42717 37791
rect 42717 37757 42751 37791
rect 42751 37757 42760 37791
rect 42708 37748 42760 37757
rect 42892 37748 42944 37800
rect 37464 37655 37516 37664
rect 37464 37621 37473 37655
rect 37473 37621 37507 37655
rect 37507 37621 37516 37655
rect 37464 37612 37516 37621
rect 42248 37612 42300 37664
rect 42432 37680 42484 37732
rect 43720 37612 43772 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 18880 37408 18932 37460
rect 23204 37408 23256 37460
rect 19524 37315 19576 37324
rect 19524 37281 19533 37315
rect 19533 37281 19567 37315
rect 19567 37281 19576 37315
rect 19524 37272 19576 37281
rect 25228 37408 25280 37460
rect 25596 37408 25648 37460
rect 32036 37408 32088 37460
rect 32680 37451 32732 37460
rect 32680 37417 32689 37451
rect 32689 37417 32723 37451
rect 32723 37417 32732 37451
rect 32680 37408 32732 37417
rect 33416 37408 33468 37460
rect 34796 37408 34848 37460
rect 37280 37451 37332 37460
rect 37280 37417 37289 37451
rect 37289 37417 37323 37451
rect 37323 37417 37332 37451
rect 37280 37408 37332 37417
rect 41696 37451 41748 37460
rect 41696 37417 41705 37451
rect 41705 37417 41739 37451
rect 41739 37417 41748 37451
rect 41696 37408 41748 37417
rect 25044 37340 25096 37392
rect 24860 37272 24912 37324
rect 24952 37315 25004 37324
rect 24952 37281 24961 37315
rect 24961 37281 24995 37315
rect 24995 37281 25004 37315
rect 27436 37340 27488 37392
rect 42708 37408 42760 37460
rect 24952 37272 25004 37281
rect 27528 37272 27580 37324
rect 1400 37247 1452 37256
rect 1400 37213 1409 37247
rect 1409 37213 1443 37247
rect 1443 37213 1452 37247
rect 1400 37204 1452 37213
rect 3240 37247 3292 37256
rect 3240 37213 3249 37247
rect 3249 37213 3283 37247
rect 3283 37213 3292 37247
rect 3240 37204 3292 37213
rect 17316 37204 17368 37256
rect 17776 37204 17828 37256
rect 18604 37204 18656 37256
rect 20168 37204 20220 37256
rect 20536 37204 20588 37256
rect 24676 37204 24728 37256
rect 24768 37247 24820 37256
rect 24768 37213 24777 37247
rect 24777 37213 24811 37247
rect 24811 37213 24820 37247
rect 24768 37204 24820 37213
rect 27988 37272 28040 37324
rect 33048 37315 33100 37324
rect 33048 37281 33057 37315
rect 33057 37281 33091 37315
rect 33091 37281 33100 37315
rect 33048 37272 33100 37281
rect 2688 37136 2740 37188
rect 17592 37136 17644 37188
rect 25872 37179 25924 37188
rect 25872 37145 25881 37179
rect 25881 37145 25915 37179
rect 25915 37145 25924 37179
rect 25872 37136 25924 37145
rect 27528 37179 27580 37188
rect 27528 37145 27537 37179
rect 27537 37145 27571 37179
rect 27571 37145 27580 37179
rect 27528 37136 27580 37145
rect 21180 37068 21232 37120
rect 27252 37111 27304 37120
rect 27252 37077 27261 37111
rect 27261 37077 27295 37111
rect 27295 37077 27304 37111
rect 27252 37068 27304 37077
rect 27620 37068 27672 37120
rect 28448 37204 28500 37256
rect 30748 37204 30800 37256
rect 31300 37204 31352 37256
rect 35348 37272 35400 37324
rect 39120 37272 39172 37324
rect 41604 37315 41656 37324
rect 41604 37281 41613 37315
rect 41613 37281 41647 37315
rect 41647 37281 41656 37315
rect 41604 37272 41656 37281
rect 32588 37136 32640 37188
rect 28724 37068 28776 37120
rect 32404 37068 32456 37120
rect 32956 37136 33008 37188
rect 34152 37204 34204 37256
rect 34796 37247 34848 37256
rect 34796 37213 34805 37247
rect 34805 37213 34839 37247
rect 34839 37213 34848 37247
rect 34796 37204 34848 37213
rect 37372 37204 37424 37256
rect 39304 37247 39356 37256
rect 39304 37213 39313 37247
rect 39313 37213 39347 37247
rect 39347 37213 39356 37247
rect 39304 37204 39356 37213
rect 41420 37247 41472 37256
rect 41420 37213 41429 37247
rect 41429 37213 41463 37247
rect 41463 37213 41472 37247
rect 41420 37204 41472 37213
rect 37648 37136 37700 37188
rect 39948 37136 40000 37188
rect 41880 37179 41932 37188
rect 41880 37145 41889 37179
rect 41889 37145 41923 37179
rect 41923 37145 41932 37179
rect 41880 37136 41932 37145
rect 42248 37136 42300 37188
rect 37740 37068 37792 37120
rect 38936 37068 38988 37120
rect 40224 37068 40276 37120
rect 43812 37111 43864 37120
rect 43812 37077 43821 37111
rect 43821 37077 43855 37111
rect 43855 37077 43864 37111
rect 43812 37068 43864 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 2688 36907 2740 36916
rect 2688 36873 2697 36907
rect 2697 36873 2731 36907
rect 2731 36873 2740 36907
rect 2688 36864 2740 36873
rect 20260 36864 20312 36916
rect 20352 36864 20404 36916
rect 24308 36907 24360 36916
rect 7932 36728 7984 36780
rect 18880 36796 18932 36848
rect 19340 36796 19392 36848
rect 21180 36796 21232 36848
rect 22008 36796 22060 36848
rect 24308 36873 24317 36907
rect 24317 36873 24351 36907
rect 24351 36873 24360 36907
rect 24308 36864 24360 36873
rect 18420 36728 18472 36780
rect 20260 36728 20312 36780
rect 20444 36771 20496 36780
rect 20444 36737 20453 36771
rect 20453 36737 20487 36771
rect 20487 36737 20496 36771
rect 20444 36728 20496 36737
rect 20628 36771 20680 36780
rect 20628 36737 20637 36771
rect 20637 36737 20671 36771
rect 20671 36737 20680 36771
rect 20628 36728 20680 36737
rect 20720 36771 20772 36780
rect 20720 36737 20729 36771
rect 20729 36737 20763 36771
rect 20763 36737 20772 36771
rect 20720 36728 20772 36737
rect 17592 36703 17644 36712
rect 17592 36669 17601 36703
rect 17601 36669 17635 36703
rect 17635 36669 17644 36703
rect 17592 36660 17644 36669
rect 20812 36660 20864 36712
rect 21732 36728 21784 36780
rect 23756 36796 23808 36848
rect 30748 36864 30800 36916
rect 30932 36864 30984 36916
rect 16856 36592 16908 36644
rect 17132 36592 17184 36644
rect 19432 36592 19484 36644
rect 19892 36592 19944 36644
rect 22376 36660 22428 36712
rect 21916 36592 21968 36644
rect 23664 36728 23716 36780
rect 25044 36771 25096 36780
rect 25044 36737 25053 36771
rect 25053 36737 25087 36771
rect 25087 36737 25096 36771
rect 25044 36728 25096 36737
rect 26332 36771 26384 36780
rect 26332 36737 26341 36771
rect 26341 36737 26375 36771
rect 26375 36737 26384 36771
rect 26332 36728 26384 36737
rect 26424 36771 26476 36780
rect 26424 36737 26433 36771
rect 26433 36737 26467 36771
rect 26467 36737 26476 36771
rect 27712 36771 27764 36780
rect 26424 36728 26476 36737
rect 27712 36737 27716 36771
rect 27716 36737 27750 36771
rect 27750 36737 27764 36771
rect 27712 36728 27764 36737
rect 24676 36660 24728 36712
rect 26056 36660 26108 36712
rect 26332 36592 26384 36644
rect 16672 36567 16724 36576
rect 16672 36533 16681 36567
rect 16681 36533 16715 36567
rect 16715 36533 16724 36567
rect 16672 36524 16724 36533
rect 18420 36524 18472 36576
rect 20812 36567 20864 36576
rect 20812 36533 20821 36567
rect 20821 36533 20855 36567
rect 20855 36533 20864 36567
rect 20812 36524 20864 36533
rect 22192 36524 22244 36576
rect 26148 36524 26200 36576
rect 27436 36524 27488 36576
rect 27896 36771 27948 36780
rect 27896 36737 27905 36771
rect 27905 36737 27939 36771
rect 27939 36737 27948 36771
rect 28080 36771 28132 36780
rect 27896 36728 27948 36737
rect 28080 36737 28088 36771
rect 28088 36737 28122 36771
rect 28122 36737 28132 36771
rect 28080 36728 28132 36737
rect 28724 36796 28776 36848
rect 28816 36771 28868 36780
rect 28816 36737 28825 36771
rect 28825 36737 28859 36771
rect 28859 36737 28868 36771
rect 28816 36728 28868 36737
rect 32312 36771 32364 36780
rect 32312 36737 32321 36771
rect 32321 36737 32355 36771
rect 32355 36737 32364 36771
rect 32312 36728 32364 36737
rect 28356 36524 28408 36576
rect 28908 36524 28960 36576
rect 31300 36524 31352 36576
rect 32220 36592 32272 36644
rect 32956 36660 33008 36712
rect 34152 36864 34204 36916
rect 40776 36864 40828 36916
rect 41604 36907 41656 36916
rect 41604 36873 41613 36907
rect 41613 36873 41647 36907
rect 41647 36873 41656 36907
rect 41604 36864 41656 36873
rect 41696 36907 41748 36916
rect 41696 36873 41705 36907
rect 41705 36873 41739 36907
rect 41739 36873 41748 36907
rect 42432 36907 42484 36916
rect 41696 36864 41748 36873
rect 42432 36873 42441 36907
rect 42441 36873 42475 36907
rect 42475 36873 42484 36907
rect 42432 36864 42484 36873
rect 43260 36907 43312 36916
rect 43260 36873 43269 36907
rect 43269 36873 43303 36907
rect 43303 36873 43312 36907
rect 43260 36864 43312 36873
rect 34520 36796 34572 36848
rect 35992 36796 36044 36848
rect 39948 36796 40000 36848
rect 41420 36796 41472 36848
rect 34704 36728 34756 36780
rect 35440 36728 35492 36780
rect 38660 36771 38712 36780
rect 38660 36737 38669 36771
rect 38669 36737 38703 36771
rect 38703 36737 38712 36771
rect 38660 36728 38712 36737
rect 38936 36771 38988 36780
rect 38936 36737 38970 36771
rect 38970 36737 38988 36771
rect 38936 36728 38988 36737
rect 41972 36796 42024 36848
rect 36176 36660 36228 36712
rect 43812 36728 43864 36780
rect 41972 36660 42024 36712
rect 42892 36660 42944 36712
rect 32496 36567 32548 36576
rect 32496 36533 32505 36567
rect 32505 36533 32539 36567
rect 32539 36533 32548 36567
rect 42064 36592 42116 36644
rect 32496 36524 32548 36533
rect 34796 36524 34848 36576
rect 40040 36567 40092 36576
rect 40040 36533 40049 36567
rect 40049 36533 40083 36567
rect 40083 36533 40092 36567
rect 40040 36524 40092 36533
rect 41696 36524 41748 36576
rect 44180 36567 44232 36576
rect 44180 36533 44189 36567
rect 44189 36533 44223 36567
rect 44223 36533 44232 36567
rect 44180 36524 44232 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 18604 36363 18656 36372
rect 18604 36329 18613 36363
rect 18613 36329 18647 36363
rect 18647 36329 18656 36363
rect 18604 36320 18656 36329
rect 20076 36295 20128 36304
rect 20076 36261 20085 36295
rect 20085 36261 20119 36295
rect 20119 36261 20128 36295
rect 20076 36252 20128 36261
rect 20536 36320 20588 36372
rect 21548 36320 21600 36372
rect 21732 36320 21784 36372
rect 22100 36363 22152 36372
rect 22100 36329 22109 36363
rect 22109 36329 22143 36363
rect 22143 36329 22152 36363
rect 26240 36363 26292 36372
rect 22100 36320 22152 36329
rect 26240 36329 26249 36363
rect 26249 36329 26283 36363
rect 26283 36329 26292 36363
rect 26240 36320 26292 36329
rect 27252 36320 27304 36372
rect 27804 36320 27856 36372
rect 32312 36320 32364 36372
rect 33600 36320 33652 36372
rect 34244 36320 34296 36372
rect 35440 36320 35492 36372
rect 40040 36320 40092 36372
rect 40224 36363 40276 36372
rect 40224 36329 40233 36363
rect 40233 36329 40267 36363
rect 40267 36329 40276 36363
rect 40224 36320 40276 36329
rect 18696 36227 18748 36236
rect 18696 36193 18705 36227
rect 18705 36193 18739 36227
rect 18739 36193 18748 36227
rect 18696 36184 18748 36193
rect 15844 36116 15896 36168
rect 16672 36116 16724 36168
rect 17776 36159 17828 36168
rect 17776 36125 17785 36159
rect 17785 36125 17819 36159
rect 17819 36125 17828 36159
rect 17776 36116 17828 36125
rect 18420 36159 18472 36168
rect 18420 36125 18429 36159
rect 18429 36125 18463 36159
rect 18463 36125 18472 36159
rect 18420 36116 18472 36125
rect 19892 36116 19944 36168
rect 21824 36252 21876 36304
rect 26332 36252 26384 36304
rect 20812 36184 20864 36236
rect 20996 36159 21048 36168
rect 20996 36125 21005 36159
rect 21005 36125 21039 36159
rect 21039 36125 21048 36159
rect 20996 36116 21048 36125
rect 17592 36048 17644 36100
rect 18604 36048 18656 36100
rect 20720 36048 20772 36100
rect 21180 36116 21232 36168
rect 22008 36116 22060 36168
rect 22376 36159 22428 36168
rect 22376 36125 22385 36159
rect 22385 36125 22419 36159
rect 22419 36125 22428 36159
rect 22652 36159 22704 36168
rect 22376 36116 22428 36125
rect 22652 36125 22660 36159
rect 22660 36125 22694 36159
rect 22694 36125 22704 36159
rect 22652 36116 22704 36125
rect 23480 36159 23532 36168
rect 23480 36125 23489 36159
rect 23489 36125 23523 36159
rect 23523 36125 23532 36159
rect 23480 36116 23532 36125
rect 26148 36159 26200 36168
rect 20628 35980 20680 36032
rect 21916 36048 21968 36100
rect 26148 36125 26157 36159
rect 26157 36125 26191 36159
rect 26191 36125 26200 36159
rect 26148 36116 26200 36125
rect 26332 36159 26384 36168
rect 26332 36125 26341 36159
rect 26341 36125 26375 36159
rect 26375 36125 26384 36159
rect 26332 36116 26384 36125
rect 27528 36252 27580 36304
rect 27712 36252 27764 36304
rect 21548 35980 21600 36032
rect 26056 36048 26108 36100
rect 27436 36156 27488 36206
rect 27436 36154 27448 36156
rect 27448 36154 27482 36156
rect 27482 36154 27488 36156
rect 27804 36116 27856 36168
rect 32496 36252 32548 36304
rect 38752 36252 38804 36304
rect 34520 36184 34572 36236
rect 36176 36227 36228 36236
rect 36176 36193 36185 36227
rect 36185 36193 36219 36227
rect 36219 36193 36228 36227
rect 36176 36184 36228 36193
rect 38844 36184 38896 36236
rect 31024 36116 31076 36168
rect 31300 36159 31352 36168
rect 31300 36125 31309 36159
rect 31309 36125 31343 36159
rect 31343 36125 31352 36159
rect 31300 36116 31352 36125
rect 32496 36116 32548 36168
rect 38936 36116 38988 36168
rect 40500 36252 40552 36304
rect 40040 36159 40092 36168
rect 40040 36125 40049 36159
rect 40049 36125 40083 36159
rect 40083 36125 40092 36159
rect 40040 36116 40092 36125
rect 42708 36227 42760 36236
rect 42708 36193 42717 36227
rect 42717 36193 42751 36227
rect 42751 36193 42760 36227
rect 42708 36184 42760 36193
rect 44180 36227 44232 36236
rect 44180 36193 44189 36227
rect 44189 36193 44223 36227
rect 44223 36193 44232 36227
rect 44180 36184 44232 36193
rect 40868 36159 40920 36168
rect 40868 36125 40877 36159
rect 40877 36125 40911 36159
rect 40911 36125 40920 36159
rect 40868 36116 40920 36125
rect 41512 36159 41564 36168
rect 41512 36125 41521 36159
rect 41521 36125 41555 36159
rect 41555 36125 41564 36159
rect 41512 36116 41564 36125
rect 42064 36116 42116 36168
rect 33324 36048 33376 36100
rect 33692 36048 33744 36100
rect 34152 36091 34204 36100
rect 34152 36057 34161 36091
rect 34161 36057 34195 36091
rect 34195 36057 34204 36091
rect 34152 36048 34204 36057
rect 35900 36091 35952 36100
rect 35900 36057 35918 36091
rect 35918 36057 35952 36091
rect 35900 36048 35952 36057
rect 36728 36048 36780 36100
rect 43996 36091 44048 36100
rect 43996 36057 44005 36091
rect 44005 36057 44039 36091
rect 44039 36057 44048 36091
rect 43996 36048 44048 36057
rect 23848 35980 23900 36032
rect 25596 36023 25648 36032
rect 25596 35989 25605 36023
rect 25605 35989 25639 36023
rect 25639 35989 25648 36023
rect 25596 35980 25648 35989
rect 27436 35980 27488 36032
rect 28080 35980 28132 36032
rect 29552 35980 29604 36032
rect 34704 35980 34756 36032
rect 39856 36023 39908 36032
rect 39856 35989 39865 36023
rect 39865 35989 39899 36023
rect 39899 35989 39908 36023
rect 39856 35980 39908 35989
rect 40684 36023 40736 36032
rect 40684 35989 40693 36023
rect 40693 35989 40727 36023
rect 40727 35989 40736 36023
rect 40684 35980 40736 35989
rect 41604 36023 41656 36032
rect 41604 35989 41613 36023
rect 41613 35989 41647 36023
rect 41647 35989 41656 36023
rect 41604 35980 41656 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 20444 35776 20496 35828
rect 21916 35776 21968 35828
rect 22744 35776 22796 35828
rect 23388 35776 23440 35828
rect 21640 35708 21692 35760
rect 23664 35708 23716 35760
rect 23848 35751 23900 35760
rect 23848 35717 23866 35751
rect 23866 35717 23900 35751
rect 31024 35776 31076 35828
rect 31484 35819 31536 35828
rect 31484 35785 31493 35819
rect 31493 35785 31527 35819
rect 31527 35785 31536 35819
rect 31484 35776 31536 35785
rect 39304 35819 39356 35828
rect 23848 35708 23900 35717
rect 34704 35708 34756 35760
rect 18604 35615 18656 35624
rect 18604 35581 18613 35615
rect 18613 35581 18647 35615
rect 18647 35581 18656 35615
rect 18604 35572 18656 35581
rect 20812 35640 20864 35692
rect 24308 35640 24360 35692
rect 25044 35640 25096 35692
rect 25688 35640 25740 35692
rect 27160 35683 27212 35692
rect 27160 35649 27169 35683
rect 27169 35649 27203 35683
rect 27203 35649 27212 35683
rect 27160 35640 27212 35649
rect 27620 35640 27672 35692
rect 27804 35683 27856 35692
rect 27804 35649 27813 35683
rect 27813 35649 27847 35683
rect 27847 35649 27856 35683
rect 27804 35640 27856 35649
rect 31392 35683 31444 35692
rect 31392 35649 31401 35683
rect 31401 35649 31435 35683
rect 31435 35649 31444 35683
rect 31392 35640 31444 35649
rect 33324 35640 33376 35692
rect 33692 35683 33744 35692
rect 33692 35649 33701 35683
rect 33701 35649 33735 35683
rect 33735 35649 33744 35683
rect 33692 35640 33744 35649
rect 20076 35572 20128 35624
rect 20996 35572 21048 35624
rect 33508 35615 33560 35624
rect 33508 35581 33517 35615
rect 33517 35581 33551 35615
rect 33551 35581 33560 35615
rect 33508 35572 33560 35581
rect 21272 35504 21324 35556
rect 32772 35547 32824 35556
rect 32772 35513 32781 35547
rect 32781 35513 32815 35547
rect 32815 35513 32824 35547
rect 32772 35504 32824 35513
rect 34796 35640 34848 35692
rect 34060 35572 34112 35624
rect 35900 35504 35952 35556
rect 22744 35479 22796 35488
rect 22744 35445 22753 35479
rect 22753 35445 22787 35479
rect 22787 35445 22796 35479
rect 22744 35436 22796 35445
rect 27528 35436 27580 35488
rect 28632 35436 28684 35488
rect 32956 35436 33008 35488
rect 34428 35479 34480 35488
rect 34428 35445 34437 35479
rect 34437 35445 34471 35479
rect 34471 35445 34480 35479
rect 34428 35436 34480 35445
rect 34520 35436 34572 35488
rect 38476 35640 38528 35692
rect 38752 35640 38804 35692
rect 39304 35785 39313 35819
rect 39313 35785 39347 35819
rect 39347 35785 39356 35819
rect 39304 35776 39356 35785
rect 40040 35776 40092 35828
rect 40868 35776 40920 35828
rect 40500 35683 40552 35692
rect 37464 35572 37516 35624
rect 36728 35547 36780 35556
rect 36728 35513 36737 35547
rect 36737 35513 36771 35547
rect 36771 35513 36780 35547
rect 36728 35504 36780 35513
rect 37648 35436 37700 35488
rect 39396 35436 39448 35488
rect 40500 35649 40509 35683
rect 40509 35649 40543 35683
rect 40543 35649 40552 35683
rect 40500 35640 40552 35649
rect 41696 35776 41748 35828
rect 42064 35776 42116 35828
rect 43996 35776 44048 35828
rect 39764 35572 39816 35624
rect 39672 35504 39724 35556
rect 41972 35640 42024 35692
rect 43260 35683 43312 35692
rect 43260 35649 43269 35683
rect 43269 35649 43303 35683
rect 43303 35649 43312 35683
rect 43260 35640 43312 35649
rect 43260 35436 43312 35488
rect 44180 35436 44232 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 22284 35232 22336 35284
rect 22652 35232 22704 35284
rect 22836 35232 22888 35284
rect 23480 35232 23532 35284
rect 23664 35275 23716 35284
rect 23664 35241 23673 35275
rect 23673 35241 23707 35275
rect 23707 35241 23716 35275
rect 23664 35232 23716 35241
rect 28080 35232 28132 35284
rect 28448 35232 28500 35284
rect 29184 35232 29236 35284
rect 34060 35275 34112 35284
rect 34060 35241 34069 35275
rect 34069 35241 34103 35275
rect 34103 35241 34112 35275
rect 34060 35232 34112 35241
rect 34428 35232 34480 35284
rect 35992 35275 36044 35284
rect 26424 35164 26476 35216
rect 19984 35071 20036 35080
rect 19984 35037 19993 35071
rect 19993 35037 20027 35071
rect 20027 35037 20036 35071
rect 19984 35028 20036 35037
rect 22744 35096 22796 35148
rect 23020 35096 23072 35148
rect 22652 35028 22704 35080
rect 17224 35003 17276 35012
rect 17224 34969 17233 35003
rect 17233 34969 17267 35003
rect 17267 34969 17276 35003
rect 17224 34960 17276 34969
rect 17408 35003 17460 35012
rect 17408 34969 17417 35003
rect 17417 34969 17451 35003
rect 17451 34969 17460 35003
rect 17408 34960 17460 34969
rect 23112 34960 23164 35012
rect 24492 34960 24544 35012
rect 24860 35028 24912 35080
rect 25596 35071 25648 35080
rect 25596 35037 25605 35071
rect 25605 35037 25639 35071
rect 25639 35037 25648 35071
rect 25596 35028 25648 35037
rect 25964 35071 26016 35080
rect 25964 35037 25973 35071
rect 25973 35037 26007 35071
rect 26007 35037 26016 35071
rect 25964 35028 26016 35037
rect 25136 34960 25188 35012
rect 26792 35139 26844 35148
rect 26792 35105 26801 35139
rect 26801 35105 26835 35139
rect 26835 35105 26844 35139
rect 26792 35096 26844 35105
rect 27712 35139 27764 35148
rect 27712 35105 27721 35139
rect 27721 35105 27755 35139
rect 27755 35105 27764 35139
rect 27712 35096 27764 35105
rect 28908 35096 28960 35148
rect 30932 35139 30984 35148
rect 30932 35105 30941 35139
rect 30941 35105 30975 35139
rect 30975 35105 30984 35139
rect 30932 35096 30984 35105
rect 33232 35164 33284 35216
rect 35348 35207 35400 35216
rect 35348 35173 35357 35207
rect 35357 35173 35391 35207
rect 35391 35173 35400 35207
rect 35348 35164 35400 35173
rect 35992 35241 36001 35275
rect 36001 35241 36035 35275
rect 36035 35241 36044 35275
rect 35992 35232 36044 35241
rect 39856 35232 39908 35284
rect 41696 35232 41748 35284
rect 38476 35207 38528 35216
rect 38476 35173 38485 35207
rect 38485 35173 38519 35207
rect 38519 35173 38528 35207
rect 38476 35164 38528 35173
rect 39672 35164 39724 35216
rect 32772 35096 32824 35148
rect 36084 35096 36136 35148
rect 38660 35096 38712 35148
rect 39948 35096 40000 35148
rect 42708 35139 42760 35148
rect 42708 35105 42717 35139
rect 42717 35105 42751 35139
rect 42751 35105 42760 35139
rect 42708 35096 42760 35105
rect 44180 35139 44232 35148
rect 44180 35105 44189 35139
rect 44189 35105 44223 35139
rect 44223 35105 44232 35139
rect 44180 35096 44232 35105
rect 27620 35028 27672 35080
rect 28264 35028 28316 35080
rect 26884 34960 26936 35012
rect 29828 35028 29880 35080
rect 32496 35071 32548 35080
rect 32496 35037 32505 35071
rect 32505 35037 32539 35071
rect 32539 35037 32548 35071
rect 32496 35028 32548 35037
rect 33140 35028 33192 35080
rect 34244 35028 34296 35080
rect 41604 35028 41656 35080
rect 17592 34935 17644 34944
rect 17592 34901 17601 34935
rect 17601 34901 17635 34935
rect 17635 34901 17644 34935
rect 17592 34892 17644 34901
rect 19432 34892 19484 34944
rect 23848 34892 23900 34944
rect 24952 34935 25004 34944
rect 24952 34901 24961 34935
rect 24961 34901 24995 34935
rect 24995 34901 25004 34935
rect 24952 34892 25004 34901
rect 26148 34892 26200 34944
rect 29644 34960 29696 35012
rect 30380 34960 30432 35012
rect 33324 35003 33376 35012
rect 33324 34969 33333 35003
rect 33333 34969 33367 35003
rect 33367 34969 33376 35003
rect 33324 34960 33376 34969
rect 35900 35003 35952 35012
rect 35900 34969 35909 35003
rect 35909 34969 35943 35003
rect 35943 34969 35952 35003
rect 35900 34960 35952 34969
rect 38568 34960 38620 35012
rect 40684 34960 40736 35012
rect 43628 34960 43680 35012
rect 29460 34892 29512 34944
rect 32312 34935 32364 34944
rect 32312 34901 32321 34935
rect 32321 34901 32355 34935
rect 32355 34901 32364 34935
rect 32312 34892 32364 34901
rect 38936 34892 38988 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 17408 34688 17460 34740
rect 19984 34688 20036 34740
rect 22652 34688 22704 34740
rect 22836 34731 22888 34740
rect 22836 34697 22845 34731
rect 22845 34697 22879 34731
rect 22879 34697 22888 34731
rect 22836 34688 22888 34697
rect 23020 34688 23072 34740
rect 23848 34731 23900 34740
rect 18696 34595 18748 34604
rect 18696 34561 18705 34595
rect 18705 34561 18739 34595
rect 18739 34561 18748 34595
rect 18696 34552 18748 34561
rect 20720 34620 20772 34672
rect 21272 34663 21324 34672
rect 21272 34629 21281 34663
rect 21281 34629 21315 34663
rect 21315 34629 21324 34663
rect 21272 34620 21324 34629
rect 22192 34663 22244 34672
rect 22192 34629 22201 34663
rect 22201 34629 22235 34663
rect 22235 34629 22244 34663
rect 22192 34620 22244 34629
rect 22744 34620 22796 34672
rect 23848 34697 23857 34731
rect 23857 34697 23891 34731
rect 23891 34697 23900 34731
rect 23848 34688 23900 34697
rect 25872 34688 25924 34740
rect 27160 34688 27212 34740
rect 27620 34688 27672 34740
rect 29184 34731 29236 34740
rect 24952 34663 25004 34672
rect 19708 34595 19760 34604
rect 19708 34561 19717 34595
rect 19717 34561 19751 34595
rect 19751 34561 19760 34595
rect 19708 34552 19760 34561
rect 22836 34552 22888 34604
rect 23020 34595 23072 34604
rect 23020 34561 23029 34595
rect 23029 34561 23063 34595
rect 23063 34561 23072 34595
rect 23020 34552 23072 34561
rect 23204 34595 23256 34604
rect 23204 34561 23213 34595
rect 23213 34561 23247 34595
rect 23247 34561 23256 34595
rect 23388 34595 23440 34604
rect 23204 34552 23256 34561
rect 23388 34561 23397 34595
rect 23397 34561 23431 34595
rect 23431 34561 23440 34595
rect 23388 34552 23440 34561
rect 24032 34595 24084 34604
rect 15384 34484 15436 34536
rect 15844 34484 15896 34536
rect 24032 34561 24041 34595
rect 24041 34561 24075 34595
rect 24075 34561 24084 34595
rect 24032 34552 24084 34561
rect 24308 34552 24360 34604
rect 24952 34629 24986 34663
rect 24986 34629 25004 34663
rect 24952 34620 25004 34629
rect 28908 34663 28960 34672
rect 25780 34552 25832 34604
rect 27436 34552 27488 34604
rect 27988 34552 28040 34604
rect 28632 34595 28684 34604
rect 28632 34561 28641 34595
rect 28641 34561 28675 34595
rect 28675 34561 28684 34595
rect 28632 34552 28684 34561
rect 28908 34629 28917 34663
rect 28917 34629 28951 34663
rect 28951 34629 28960 34663
rect 28908 34620 28960 34629
rect 29184 34697 29193 34731
rect 29193 34697 29227 34731
rect 29227 34697 29236 34731
rect 29184 34688 29236 34697
rect 29644 34731 29696 34740
rect 29644 34697 29653 34731
rect 29653 34697 29687 34731
rect 29687 34697 29696 34731
rect 29644 34688 29696 34697
rect 31392 34688 31444 34740
rect 32588 34688 32640 34740
rect 33048 34688 33100 34740
rect 38200 34688 38252 34740
rect 38476 34688 38528 34740
rect 41512 34688 41564 34740
rect 43628 34731 43680 34740
rect 43628 34697 43637 34731
rect 43637 34697 43671 34731
rect 43671 34697 43680 34731
rect 43628 34688 43680 34697
rect 29000 34595 29052 34604
rect 29000 34561 29009 34595
rect 29009 34561 29043 34595
rect 29043 34561 29052 34595
rect 29644 34595 29696 34604
rect 29000 34552 29052 34561
rect 29644 34561 29653 34595
rect 29653 34561 29687 34595
rect 29687 34561 29696 34595
rect 29644 34552 29696 34561
rect 30472 34595 30524 34604
rect 30472 34561 30481 34595
rect 30481 34561 30515 34595
rect 30515 34561 30524 34595
rect 30472 34552 30524 34561
rect 32772 34620 32824 34672
rect 34520 34552 34572 34604
rect 37372 34595 37424 34604
rect 37372 34561 37381 34595
rect 37381 34561 37415 34595
rect 37415 34561 37424 34595
rect 37372 34552 37424 34561
rect 38568 34552 38620 34604
rect 38936 34595 38988 34604
rect 37648 34527 37700 34536
rect 22284 34416 22336 34468
rect 27528 34416 27580 34468
rect 37648 34493 37657 34527
rect 37657 34493 37691 34527
rect 37691 34493 37700 34527
rect 37648 34484 37700 34493
rect 38384 34484 38436 34536
rect 38936 34561 38945 34595
rect 38945 34561 38979 34595
rect 38979 34561 38988 34595
rect 38936 34552 38988 34561
rect 39764 34552 39816 34604
rect 40132 34595 40184 34604
rect 40132 34561 40141 34595
rect 40141 34561 40175 34595
rect 40175 34561 40184 34595
rect 40132 34552 40184 34561
rect 41696 34552 41748 34604
rect 43628 34552 43680 34604
rect 40040 34484 40092 34536
rect 41236 34527 41288 34536
rect 41236 34493 41245 34527
rect 41245 34493 41279 34527
rect 41279 34493 41288 34527
rect 41236 34484 41288 34493
rect 20996 34348 21048 34400
rect 33140 34416 33192 34468
rect 41972 34416 42024 34468
rect 33048 34391 33100 34400
rect 33048 34357 33057 34391
rect 33057 34357 33091 34391
rect 33091 34357 33100 34391
rect 33048 34348 33100 34357
rect 38752 34348 38804 34400
rect 40224 34348 40276 34400
rect 42340 34348 42392 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 16948 34144 17000 34196
rect 17224 34144 17276 34196
rect 19708 34144 19760 34196
rect 15384 34051 15436 34060
rect 15384 34017 15393 34051
rect 15393 34017 15427 34051
rect 15427 34017 15436 34051
rect 15384 34008 15436 34017
rect 17408 34008 17460 34060
rect 22836 34144 22888 34196
rect 23388 34144 23440 34196
rect 24860 34187 24912 34196
rect 24860 34153 24869 34187
rect 24869 34153 24903 34187
rect 24903 34153 24912 34187
rect 24860 34144 24912 34153
rect 26884 34144 26936 34196
rect 27804 34144 27856 34196
rect 28356 34187 28408 34196
rect 28356 34153 28365 34187
rect 28365 34153 28399 34187
rect 28399 34153 28408 34187
rect 28356 34144 28408 34153
rect 30380 34144 30432 34196
rect 20812 34076 20864 34128
rect 20720 34008 20772 34060
rect 17868 33940 17920 33992
rect 19984 33983 20036 33992
rect 19984 33949 19993 33983
rect 19993 33949 20027 33983
rect 20027 33949 20036 33983
rect 19984 33940 20036 33949
rect 16212 33872 16264 33924
rect 20260 33983 20312 33992
rect 20260 33949 20295 33983
rect 20295 33949 20312 33983
rect 22376 34076 22428 34128
rect 23296 34076 23348 34128
rect 20260 33940 20312 33949
rect 20996 33915 21048 33924
rect 12164 33804 12216 33856
rect 18880 33804 18932 33856
rect 20996 33881 21005 33915
rect 21005 33881 21039 33915
rect 21039 33881 21048 33915
rect 20996 33872 21048 33881
rect 22100 33940 22152 33992
rect 24032 34008 24084 34060
rect 22284 33940 22336 33992
rect 22376 33983 22428 33992
rect 22376 33949 22385 33983
rect 22385 33949 22419 33983
rect 22419 33949 22428 33983
rect 22376 33940 22428 33949
rect 21824 33872 21876 33924
rect 25136 33983 25188 33992
rect 25136 33949 25145 33983
rect 25145 33949 25179 33983
rect 25179 33949 25188 33983
rect 25136 33940 25188 33949
rect 25504 33940 25556 33992
rect 25688 33983 25740 33992
rect 25688 33949 25697 33983
rect 25697 33949 25731 33983
rect 25731 33949 25740 33983
rect 25688 33940 25740 33949
rect 25872 33983 25924 33992
rect 25872 33949 25881 33983
rect 25881 33949 25915 33983
rect 25915 33949 25924 33983
rect 25872 33940 25924 33949
rect 26884 33983 26936 33992
rect 26884 33949 26893 33983
rect 26893 33949 26927 33983
rect 26927 33949 26936 33983
rect 26884 33940 26936 33949
rect 27160 33983 27212 33992
rect 27160 33949 27169 33983
rect 27169 33949 27203 33983
rect 27203 33949 27212 33983
rect 27160 33940 27212 33949
rect 27528 33940 27580 33992
rect 29644 34008 29696 34060
rect 30932 34144 30984 34196
rect 31668 34144 31720 34196
rect 32496 34144 32548 34196
rect 37372 34144 37424 34196
rect 31944 34119 31996 34128
rect 31944 34085 31953 34119
rect 31953 34085 31987 34119
rect 31987 34085 31996 34119
rect 31944 34076 31996 34085
rect 32956 34076 33008 34128
rect 34336 34076 34388 34128
rect 35348 34051 35400 34060
rect 35348 34017 35357 34051
rect 35357 34017 35391 34051
rect 35391 34017 35400 34051
rect 35348 34008 35400 34017
rect 36084 34076 36136 34128
rect 38568 34076 38620 34128
rect 41236 34144 41288 34196
rect 39948 34051 40000 34060
rect 39948 34017 39957 34051
rect 39957 34017 39991 34051
rect 39991 34017 40000 34051
rect 39948 34008 40000 34017
rect 42340 34051 42392 34060
rect 42340 34017 42349 34051
rect 42349 34017 42383 34051
rect 42383 34017 42392 34051
rect 42340 34008 42392 34017
rect 44088 34051 44140 34060
rect 44088 34017 44097 34051
rect 44097 34017 44131 34051
rect 44131 34017 44140 34051
rect 44088 34008 44140 34017
rect 28264 33983 28316 33992
rect 28264 33949 28273 33983
rect 28273 33949 28307 33983
rect 28307 33949 28316 33983
rect 28264 33940 28316 33949
rect 29460 33940 29512 33992
rect 32128 33940 32180 33992
rect 32588 33983 32640 33992
rect 32588 33949 32597 33983
rect 32597 33949 32631 33983
rect 32631 33949 32640 33983
rect 32588 33940 32640 33949
rect 33140 33940 33192 33992
rect 33416 33940 33468 33992
rect 34244 33940 34296 33992
rect 35440 33940 35492 33992
rect 36912 33940 36964 33992
rect 22192 33804 22244 33856
rect 26976 33872 27028 33924
rect 29000 33872 29052 33924
rect 31484 33872 31536 33924
rect 27436 33804 27488 33856
rect 33968 33872 34020 33924
rect 36176 33872 36228 33924
rect 34060 33847 34112 33856
rect 34060 33813 34069 33847
rect 34069 33813 34103 33847
rect 34103 33813 34112 33847
rect 34060 33804 34112 33813
rect 34796 33847 34848 33856
rect 34796 33813 34805 33847
rect 34805 33813 34839 33847
rect 34839 33813 34848 33847
rect 34796 33804 34848 33813
rect 35624 33804 35676 33856
rect 36268 33847 36320 33856
rect 36268 33813 36277 33847
rect 36277 33813 36311 33847
rect 36311 33813 36320 33847
rect 36268 33804 36320 33813
rect 36360 33847 36412 33856
rect 36360 33813 36369 33847
rect 36369 33813 36403 33847
rect 36403 33813 36412 33847
rect 37188 33983 37240 33992
rect 37188 33949 37197 33983
rect 37197 33949 37231 33983
rect 37231 33949 37240 33983
rect 37188 33940 37240 33949
rect 38844 33940 38896 33992
rect 40224 33983 40276 33992
rect 40224 33949 40258 33983
rect 40258 33949 40276 33983
rect 40224 33940 40276 33949
rect 38752 33915 38804 33924
rect 38752 33881 38761 33915
rect 38761 33881 38795 33915
rect 38795 33881 38804 33915
rect 38752 33872 38804 33881
rect 43536 33872 43588 33924
rect 36360 33804 36412 33813
rect 37280 33804 37332 33856
rect 39120 33804 39172 33856
rect 40040 33804 40092 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 18604 33600 18656 33652
rect 18696 33600 18748 33652
rect 18880 33600 18932 33652
rect 35992 33600 36044 33652
rect 36268 33600 36320 33652
rect 37556 33600 37608 33652
rect 38384 33643 38436 33652
rect 38384 33609 38409 33643
rect 38409 33609 38436 33643
rect 38384 33600 38436 33609
rect 19340 33532 19392 33584
rect 19432 33532 19484 33584
rect 19984 33532 20036 33584
rect 22376 33532 22428 33584
rect 23296 33532 23348 33584
rect 24492 33575 24544 33584
rect 24492 33541 24501 33575
rect 24501 33541 24535 33575
rect 24535 33541 24544 33575
rect 24492 33532 24544 33541
rect 31484 33575 31536 33584
rect 16948 33507 17000 33516
rect 16948 33473 16957 33507
rect 16957 33473 16991 33507
rect 16991 33473 17000 33507
rect 16948 33464 17000 33473
rect 17592 33464 17644 33516
rect 17776 33464 17828 33516
rect 16488 33328 16540 33380
rect 17868 33396 17920 33448
rect 20260 33464 20312 33516
rect 20720 33464 20772 33516
rect 21272 33507 21324 33516
rect 21272 33473 21281 33507
rect 21281 33473 21315 33507
rect 21315 33473 21324 33507
rect 21272 33464 21324 33473
rect 19248 33439 19300 33448
rect 19248 33405 19257 33439
rect 19257 33405 19291 33439
rect 19291 33405 19300 33439
rect 19248 33396 19300 33405
rect 20812 33396 20864 33448
rect 22468 33464 22520 33516
rect 23664 33507 23716 33516
rect 23664 33473 23673 33507
rect 23673 33473 23707 33507
rect 23707 33473 23716 33507
rect 23664 33464 23716 33473
rect 25964 33507 26016 33516
rect 25964 33473 25973 33507
rect 25973 33473 26007 33507
rect 26007 33473 26016 33507
rect 25964 33464 26016 33473
rect 27160 33507 27212 33516
rect 22192 33396 22244 33448
rect 22744 33439 22796 33448
rect 22744 33405 22753 33439
rect 22753 33405 22787 33439
rect 22787 33405 22796 33439
rect 22744 33396 22796 33405
rect 23204 33396 23256 33448
rect 25688 33396 25740 33448
rect 26056 33396 26108 33448
rect 27160 33473 27169 33507
rect 27169 33473 27203 33507
rect 27203 33473 27212 33507
rect 27160 33464 27212 33473
rect 27804 33464 27856 33516
rect 28080 33507 28132 33516
rect 28080 33473 28089 33507
rect 28089 33473 28123 33507
rect 28123 33473 28132 33507
rect 28080 33464 28132 33473
rect 29460 33507 29512 33516
rect 29460 33473 29469 33507
rect 29469 33473 29503 33507
rect 29503 33473 29512 33507
rect 29460 33464 29512 33473
rect 27988 33439 28040 33448
rect 27988 33405 27997 33439
rect 27997 33405 28031 33439
rect 28031 33405 28040 33439
rect 27988 33396 28040 33405
rect 28264 33396 28316 33448
rect 28632 33396 28684 33448
rect 17960 33328 18012 33380
rect 20720 33328 20772 33380
rect 21824 33328 21876 33380
rect 24768 33328 24820 33380
rect 25780 33371 25832 33380
rect 25780 33337 25789 33371
rect 25789 33337 25823 33371
rect 25823 33337 25832 33371
rect 25780 33328 25832 33337
rect 26976 33328 27028 33380
rect 31484 33541 31493 33575
rect 31493 33541 31527 33575
rect 31527 33541 31536 33575
rect 31484 33532 31536 33541
rect 32496 33532 32548 33584
rect 34244 33575 34296 33584
rect 34244 33541 34253 33575
rect 34253 33541 34287 33575
rect 34287 33541 34296 33575
rect 34244 33532 34296 33541
rect 35440 33532 35492 33584
rect 31668 33464 31720 33516
rect 32680 33464 32732 33516
rect 33968 33507 34020 33516
rect 33968 33473 33977 33507
rect 33977 33473 34011 33507
rect 34011 33473 34020 33507
rect 33968 33464 34020 33473
rect 34060 33464 34112 33516
rect 36176 33464 36228 33516
rect 38200 33575 38252 33584
rect 38200 33541 38209 33575
rect 38209 33541 38243 33575
rect 38243 33541 38252 33575
rect 38200 33532 38252 33541
rect 40132 33600 40184 33652
rect 43536 33643 43588 33652
rect 43536 33609 43545 33643
rect 43545 33609 43579 33643
rect 43579 33609 43588 33643
rect 43536 33600 43588 33609
rect 38844 33532 38896 33584
rect 40040 33532 40092 33584
rect 37556 33507 37608 33516
rect 32036 33396 32088 33448
rect 33140 33396 33192 33448
rect 16672 33260 16724 33312
rect 18604 33260 18656 33312
rect 21364 33260 21416 33312
rect 22376 33260 22428 33312
rect 27068 33303 27120 33312
rect 27068 33269 27077 33303
rect 27077 33269 27111 33303
rect 27111 33269 27120 33303
rect 27068 33260 27120 33269
rect 27896 33260 27948 33312
rect 33416 33328 33468 33380
rect 33140 33260 33192 33312
rect 33232 33260 33284 33312
rect 34336 33396 34388 33448
rect 35440 33396 35492 33448
rect 36452 33396 36504 33448
rect 37188 33396 37240 33448
rect 35992 33328 36044 33380
rect 36084 33260 36136 33312
rect 36636 33303 36688 33312
rect 36636 33269 36645 33303
rect 36645 33269 36679 33303
rect 36679 33269 36688 33303
rect 36636 33260 36688 33269
rect 36912 33328 36964 33380
rect 37556 33473 37565 33507
rect 37565 33473 37599 33507
rect 37599 33473 37608 33507
rect 37556 33464 37608 33473
rect 38568 33464 38620 33516
rect 39764 33464 39816 33516
rect 43076 33464 43128 33516
rect 43444 33507 43496 33516
rect 43444 33473 43453 33507
rect 43453 33473 43487 33507
rect 43487 33473 43496 33507
rect 43444 33464 43496 33473
rect 38936 33328 38988 33380
rect 42892 33303 42944 33312
rect 42892 33269 42901 33303
rect 42901 33269 42935 33303
rect 42935 33269 42944 33303
rect 42892 33260 42944 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 16212 33099 16264 33108
rect 16212 33065 16221 33099
rect 16221 33065 16255 33099
rect 16255 33065 16264 33099
rect 16212 33056 16264 33065
rect 19340 33056 19392 33108
rect 23664 33056 23716 33108
rect 26056 33099 26108 33108
rect 26056 33065 26065 33099
rect 26065 33065 26099 33099
rect 26099 33065 26108 33099
rect 26056 33056 26108 33065
rect 32036 33056 32088 33108
rect 32680 33099 32732 33108
rect 32680 33065 32689 33099
rect 32689 33065 32723 33099
rect 32723 33065 32732 33099
rect 32680 33056 32732 33065
rect 34704 33056 34756 33108
rect 36268 33056 36320 33108
rect 36452 33099 36504 33108
rect 36452 33065 36461 33099
rect 36461 33065 36495 33099
rect 36495 33065 36504 33099
rect 36452 33056 36504 33065
rect 37556 33056 37608 33108
rect 13912 32988 13964 33040
rect 19248 32988 19300 33040
rect 27252 33031 27304 33040
rect 27252 32997 27261 33031
rect 27261 32997 27295 33031
rect 27295 32997 27304 33031
rect 27252 32988 27304 32997
rect 27620 32988 27672 33040
rect 28080 32988 28132 33040
rect 33968 32988 34020 33040
rect 16396 32920 16448 32972
rect 17868 32963 17920 32972
rect 15752 32895 15804 32904
rect 15752 32861 15761 32895
rect 15761 32861 15795 32895
rect 15795 32861 15804 32895
rect 15752 32852 15804 32861
rect 16488 32895 16540 32904
rect 16488 32861 16497 32895
rect 16497 32861 16531 32895
rect 16531 32861 16540 32895
rect 16488 32852 16540 32861
rect 17868 32929 17877 32963
rect 17877 32929 17911 32963
rect 17911 32929 17920 32963
rect 17868 32920 17920 32929
rect 17960 32920 18012 32972
rect 16672 32895 16724 32904
rect 16672 32861 16681 32895
rect 16681 32861 16715 32895
rect 16715 32861 16724 32895
rect 18512 32920 18564 32972
rect 16672 32852 16724 32861
rect 18420 32852 18472 32904
rect 19156 32784 19208 32836
rect 21180 32852 21232 32904
rect 25688 32852 25740 32904
rect 27804 32920 27856 32972
rect 32128 32920 32180 32972
rect 33232 32920 33284 32972
rect 35348 32988 35400 33040
rect 35900 32988 35952 33040
rect 36360 32988 36412 33040
rect 38660 32963 38712 32972
rect 27620 32852 27672 32904
rect 27712 32895 27764 32904
rect 27712 32861 27721 32895
rect 27721 32861 27755 32895
rect 27755 32861 27764 32895
rect 27896 32895 27948 32904
rect 27712 32852 27764 32861
rect 27896 32861 27905 32895
rect 27905 32861 27939 32895
rect 27939 32861 27948 32895
rect 27896 32852 27948 32861
rect 22836 32784 22888 32836
rect 24952 32827 25004 32836
rect 24952 32793 24986 32827
rect 24986 32793 25004 32827
rect 24952 32784 25004 32793
rect 27344 32784 27396 32836
rect 28356 32852 28408 32904
rect 31944 32895 31996 32904
rect 31944 32861 31953 32895
rect 31953 32861 31987 32895
rect 31987 32861 31996 32895
rect 31944 32852 31996 32861
rect 32312 32852 32364 32904
rect 33048 32852 33100 32904
rect 33140 32852 33192 32904
rect 35716 32852 35768 32904
rect 38660 32929 38669 32963
rect 38669 32929 38703 32963
rect 38703 32929 38712 32963
rect 38660 32920 38712 32929
rect 42892 32920 42944 32972
rect 44088 32963 44140 32972
rect 44088 32929 44097 32963
rect 44097 32929 44131 32963
rect 44131 32929 44140 32963
rect 44088 32920 44140 32929
rect 36360 32852 36412 32904
rect 39120 32895 39172 32904
rect 39120 32861 39129 32895
rect 39129 32861 39163 32895
rect 39163 32861 39172 32895
rect 39120 32852 39172 32861
rect 42340 32895 42392 32904
rect 42340 32861 42349 32895
rect 42349 32861 42383 32895
rect 42383 32861 42392 32895
rect 42340 32852 42392 32861
rect 19432 32716 19484 32768
rect 21364 32716 21416 32768
rect 23848 32716 23900 32768
rect 26884 32759 26936 32768
rect 26884 32725 26893 32759
rect 26893 32725 26927 32759
rect 26927 32725 26936 32759
rect 26884 32716 26936 32725
rect 27712 32716 27764 32768
rect 30932 32784 30984 32836
rect 35532 32784 35584 32836
rect 36912 32784 36964 32836
rect 37372 32784 37424 32836
rect 28356 32759 28408 32768
rect 28356 32725 28365 32759
rect 28365 32725 28399 32759
rect 28399 32725 28408 32759
rect 28356 32716 28408 32725
rect 39948 32716 40000 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 16764 32512 16816 32564
rect 15568 32419 15620 32428
rect 15568 32385 15577 32419
rect 15577 32385 15611 32419
rect 15611 32385 15620 32419
rect 15568 32376 15620 32385
rect 15936 32419 15988 32428
rect 15936 32385 15945 32419
rect 15945 32385 15979 32419
rect 15979 32385 15988 32419
rect 15936 32376 15988 32385
rect 16396 32444 16448 32496
rect 16212 32376 16264 32428
rect 16028 32308 16080 32360
rect 16396 32308 16448 32360
rect 16488 32308 16540 32360
rect 18144 32376 18196 32428
rect 18420 32376 18472 32428
rect 19432 32444 19484 32496
rect 20628 32444 20680 32496
rect 18328 32351 18380 32360
rect 14372 32172 14424 32224
rect 16212 32172 16264 32224
rect 16764 32172 16816 32224
rect 18328 32317 18337 32351
rect 18337 32317 18371 32351
rect 18371 32317 18380 32351
rect 18328 32308 18380 32317
rect 19156 32240 19208 32292
rect 18972 32172 19024 32224
rect 21272 32512 21324 32564
rect 22836 32555 22888 32564
rect 22836 32521 22845 32555
rect 22845 32521 22879 32555
rect 22879 32521 22888 32555
rect 22836 32512 22888 32521
rect 24952 32555 25004 32564
rect 24952 32521 24961 32555
rect 24961 32521 24995 32555
rect 24995 32521 25004 32555
rect 24952 32512 25004 32521
rect 22744 32444 22796 32496
rect 24492 32444 24544 32496
rect 26884 32512 26936 32564
rect 27988 32512 28040 32564
rect 28632 32555 28684 32564
rect 28632 32521 28641 32555
rect 28641 32521 28675 32555
rect 28675 32521 28684 32555
rect 28632 32512 28684 32521
rect 33968 32512 34020 32564
rect 36912 32512 36964 32564
rect 37372 32555 37424 32564
rect 37372 32521 37381 32555
rect 37381 32521 37415 32555
rect 37415 32521 37424 32555
rect 37372 32512 37424 32521
rect 38936 32512 38988 32564
rect 21364 32376 21416 32428
rect 22376 32419 22428 32428
rect 22376 32385 22385 32419
rect 22385 32385 22419 32419
rect 22419 32385 22428 32419
rect 22376 32376 22428 32385
rect 22284 32308 22336 32360
rect 23204 32376 23256 32428
rect 23296 32351 23348 32360
rect 23296 32317 23305 32351
rect 23305 32317 23339 32351
rect 23339 32317 23348 32351
rect 23296 32308 23348 32317
rect 24676 32376 24728 32428
rect 27068 32444 27120 32496
rect 25136 32308 25188 32360
rect 26056 32308 26108 32360
rect 26332 32376 26384 32428
rect 26884 32376 26936 32428
rect 27712 32444 27764 32496
rect 28356 32444 28408 32496
rect 34796 32444 34848 32496
rect 35624 32444 35676 32496
rect 36084 32444 36136 32496
rect 27804 32376 27856 32428
rect 28080 32419 28132 32428
rect 28080 32385 28089 32419
rect 28089 32385 28123 32419
rect 28123 32385 28132 32419
rect 28080 32376 28132 32385
rect 30656 32419 30708 32428
rect 30656 32385 30665 32419
rect 30665 32385 30699 32419
rect 30699 32385 30708 32419
rect 30656 32376 30708 32385
rect 35532 32419 35584 32428
rect 35532 32385 35541 32419
rect 35541 32385 35575 32419
rect 35575 32385 35584 32419
rect 35532 32376 35584 32385
rect 35716 32376 35768 32428
rect 37280 32419 37332 32428
rect 37280 32385 37289 32419
rect 37289 32385 37323 32419
rect 37323 32385 37332 32419
rect 37280 32376 37332 32385
rect 38384 32376 38436 32428
rect 39948 32419 40000 32428
rect 39948 32385 39966 32419
rect 39966 32385 40000 32419
rect 39948 32376 40000 32385
rect 42340 32376 42392 32428
rect 24216 32283 24268 32292
rect 24216 32249 24225 32283
rect 24225 32249 24259 32283
rect 24259 32249 24268 32283
rect 24216 32240 24268 32249
rect 20352 32172 20404 32224
rect 20720 32172 20772 32224
rect 22100 32172 22152 32224
rect 22284 32172 22336 32224
rect 31760 32308 31812 32360
rect 34796 32351 34848 32360
rect 34796 32317 34805 32351
rect 34805 32317 34839 32351
rect 34839 32317 34848 32351
rect 34796 32308 34848 32317
rect 26976 32283 27028 32292
rect 26976 32249 26985 32283
rect 26985 32249 27019 32283
rect 27019 32249 27028 32283
rect 26976 32240 27028 32249
rect 27344 32240 27396 32292
rect 30472 32283 30524 32292
rect 30472 32249 30481 32283
rect 30481 32249 30515 32283
rect 30515 32249 30524 32283
rect 30472 32240 30524 32249
rect 26424 32215 26476 32224
rect 26424 32181 26433 32215
rect 26433 32181 26467 32215
rect 26467 32181 26476 32215
rect 26424 32172 26476 32181
rect 35440 32172 35492 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 16672 31968 16724 32020
rect 17868 31968 17920 32020
rect 24676 32011 24728 32020
rect 15568 31900 15620 31952
rect 18328 31943 18380 31952
rect 16120 31875 16172 31884
rect 16120 31841 16129 31875
rect 16129 31841 16163 31875
rect 16163 31841 16172 31875
rect 18328 31909 18337 31943
rect 18337 31909 18371 31943
rect 18371 31909 18380 31943
rect 18328 31900 18380 31909
rect 22192 31900 22244 31952
rect 16120 31832 16172 31841
rect 13912 31764 13964 31816
rect 14372 31739 14424 31748
rect 14372 31705 14406 31739
rect 14406 31705 14424 31739
rect 16488 31764 16540 31816
rect 17776 31807 17828 31816
rect 14372 31696 14424 31705
rect 16580 31696 16632 31748
rect 16672 31696 16724 31748
rect 17776 31773 17785 31807
rect 17785 31773 17819 31807
rect 17819 31773 17828 31807
rect 17776 31764 17828 31773
rect 19248 31764 19300 31816
rect 21180 31807 21232 31816
rect 21180 31773 21189 31807
rect 21189 31773 21223 31807
rect 21223 31773 21232 31807
rect 21180 31764 21232 31773
rect 24216 31832 24268 31884
rect 24676 31977 24685 32011
rect 24685 31977 24719 32011
rect 24719 31977 24728 32011
rect 24676 31968 24728 31977
rect 25136 31968 25188 32020
rect 26884 31968 26936 32020
rect 28172 31968 28224 32020
rect 35716 31968 35768 32020
rect 30380 31900 30432 31952
rect 30656 31900 30708 31952
rect 22192 31807 22244 31816
rect 22192 31773 22201 31807
rect 22201 31773 22235 31807
rect 22235 31773 22244 31807
rect 22468 31807 22520 31816
rect 22192 31764 22244 31773
rect 22468 31773 22477 31807
rect 22477 31773 22511 31807
rect 22511 31773 22520 31807
rect 22468 31764 22520 31773
rect 23388 31764 23440 31816
rect 25688 31832 25740 31884
rect 25044 31764 25096 31816
rect 15936 31671 15988 31680
rect 15936 31637 15945 31671
rect 15945 31637 15979 31671
rect 15979 31637 15988 31671
rect 15936 31628 15988 31637
rect 17500 31628 17552 31680
rect 18512 31671 18564 31680
rect 18512 31637 18539 31671
rect 18539 31637 18564 31671
rect 18512 31628 18564 31637
rect 18972 31696 19024 31748
rect 20352 31739 20404 31748
rect 20352 31705 20370 31739
rect 20370 31705 20404 31739
rect 20352 31696 20404 31705
rect 22744 31696 22796 31748
rect 23296 31739 23348 31748
rect 23296 31705 23318 31739
rect 23318 31705 23348 31739
rect 23296 31696 23348 31705
rect 26424 31764 26476 31816
rect 29644 31807 29696 31816
rect 29644 31773 29653 31807
rect 29653 31773 29687 31807
rect 29687 31773 29696 31807
rect 29644 31764 29696 31773
rect 30288 31764 30340 31816
rect 32128 31832 32180 31884
rect 31760 31764 31812 31816
rect 32772 31764 32824 31816
rect 34796 31807 34848 31816
rect 34796 31773 34805 31807
rect 34805 31773 34839 31807
rect 34839 31773 34848 31807
rect 34796 31764 34848 31773
rect 35440 31764 35492 31816
rect 36636 31764 36688 31816
rect 25964 31739 26016 31748
rect 19156 31628 19208 31680
rect 23112 31671 23164 31680
rect 23112 31637 23121 31671
rect 23121 31637 23155 31671
rect 23155 31637 23164 31671
rect 23112 31628 23164 31637
rect 25964 31705 25973 31739
rect 25973 31705 26007 31739
rect 26007 31705 26016 31739
rect 25964 31696 26016 31705
rect 26148 31696 26200 31748
rect 30472 31696 30524 31748
rect 30840 31628 30892 31680
rect 36636 31671 36688 31680
rect 36636 31637 36645 31671
rect 36645 31637 36679 31671
rect 36679 31637 36688 31671
rect 36636 31628 36688 31637
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 15568 31424 15620 31476
rect 18604 31424 18656 31476
rect 15476 31288 15528 31340
rect 15752 31288 15804 31340
rect 13912 31263 13964 31272
rect 13912 31229 13921 31263
rect 13921 31229 13955 31263
rect 13955 31229 13964 31263
rect 13912 31220 13964 31229
rect 16120 31331 16172 31340
rect 16120 31297 16129 31331
rect 16129 31297 16163 31331
rect 16163 31297 16172 31331
rect 16672 31331 16724 31340
rect 16120 31288 16172 31297
rect 16672 31297 16681 31331
rect 16681 31297 16715 31331
rect 16715 31297 16724 31331
rect 16672 31288 16724 31297
rect 19248 31356 19300 31408
rect 22284 31424 22336 31476
rect 23388 31467 23440 31476
rect 23388 31433 23397 31467
rect 23397 31433 23431 31467
rect 23431 31433 23440 31467
rect 23388 31424 23440 31433
rect 25228 31424 25280 31476
rect 26976 31424 27028 31476
rect 32128 31467 32180 31476
rect 24216 31356 24268 31408
rect 25780 31356 25832 31408
rect 28172 31356 28224 31408
rect 20168 31331 20220 31340
rect 20168 31297 20202 31331
rect 20202 31297 20220 31331
rect 20168 31288 20220 31297
rect 22284 31331 22336 31340
rect 22284 31297 22318 31331
rect 22318 31297 22336 31331
rect 22284 31288 22336 31297
rect 25872 31288 25924 31340
rect 26332 31331 26384 31340
rect 26332 31297 26341 31331
rect 26341 31297 26375 31331
rect 26375 31297 26384 31331
rect 26332 31288 26384 31297
rect 28448 31288 28500 31340
rect 31300 31356 31352 31408
rect 32128 31433 32137 31467
rect 32137 31433 32171 31467
rect 32171 31433 32180 31467
rect 32128 31424 32180 31433
rect 35348 31356 35400 31408
rect 16396 31220 16448 31272
rect 18972 31263 19024 31272
rect 18972 31229 18981 31263
rect 18981 31229 19015 31263
rect 19015 31229 19024 31263
rect 18972 31220 19024 31229
rect 19156 31220 19208 31272
rect 21180 31220 21232 31272
rect 21824 31220 21876 31272
rect 29644 31220 29696 31272
rect 30380 31220 30432 31272
rect 30748 31220 30800 31272
rect 15844 31195 15896 31204
rect 15844 31161 15853 31195
rect 15853 31161 15887 31195
rect 15887 31161 15896 31195
rect 15844 31152 15896 31161
rect 25688 31152 25740 31204
rect 26424 31152 26476 31204
rect 34796 31152 34848 31204
rect 16488 31084 16540 31136
rect 21272 31127 21324 31136
rect 21272 31093 21281 31127
rect 21281 31093 21315 31127
rect 21315 31093 21324 31127
rect 21272 31084 21324 31093
rect 25320 31127 25372 31136
rect 25320 31093 25329 31127
rect 25329 31093 25363 31127
rect 25363 31093 25372 31127
rect 25320 31084 25372 31093
rect 25964 31084 26016 31136
rect 27252 31127 27304 31136
rect 27252 31093 27261 31127
rect 27261 31093 27295 31127
rect 27295 31093 27304 31127
rect 27252 31084 27304 31093
rect 28080 31127 28132 31136
rect 28080 31093 28089 31127
rect 28089 31093 28123 31127
rect 28123 31093 28132 31127
rect 28080 31084 28132 31093
rect 31116 31084 31168 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 15476 30923 15528 30932
rect 15476 30889 15485 30923
rect 15485 30889 15519 30923
rect 15519 30889 15528 30923
rect 15476 30880 15528 30889
rect 16672 30923 16724 30932
rect 1768 30719 1820 30728
rect 1768 30685 1777 30719
rect 1777 30685 1811 30719
rect 1811 30685 1820 30719
rect 1768 30676 1820 30685
rect 16672 30889 16681 30923
rect 16681 30889 16715 30923
rect 16715 30889 16724 30923
rect 16672 30880 16724 30889
rect 15844 30855 15896 30864
rect 15844 30821 15853 30855
rect 15853 30821 15887 30855
rect 15887 30821 15896 30855
rect 15844 30812 15896 30821
rect 16396 30812 16448 30864
rect 18144 30880 18196 30932
rect 20168 30880 20220 30932
rect 22284 30880 22336 30932
rect 23756 30923 23808 30932
rect 23756 30889 23765 30923
rect 23765 30889 23799 30923
rect 23799 30889 23808 30923
rect 23756 30880 23808 30889
rect 25228 30880 25280 30932
rect 28264 30923 28316 30932
rect 28264 30889 28273 30923
rect 28273 30889 28307 30923
rect 28307 30889 28316 30923
rect 28264 30880 28316 30889
rect 28448 30923 28500 30932
rect 28448 30889 28457 30923
rect 28457 30889 28491 30923
rect 28491 30889 28500 30923
rect 28448 30880 28500 30889
rect 31116 30923 31168 30932
rect 31116 30889 31125 30923
rect 31125 30889 31159 30923
rect 31159 30889 31168 30923
rect 31116 30880 31168 30889
rect 37556 30880 37608 30932
rect 16028 30744 16080 30796
rect 15936 30719 15988 30728
rect 15936 30685 15945 30719
rect 15945 30685 15979 30719
rect 15979 30685 15988 30719
rect 16856 30744 16908 30796
rect 18604 30812 18656 30864
rect 17960 30787 18012 30796
rect 17960 30753 17969 30787
rect 17969 30753 18003 30787
rect 18003 30753 18012 30787
rect 17960 30744 18012 30753
rect 18144 30787 18196 30796
rect 18144 30753 18153 30787
rect 18153 30753 18187 30787
rect 18187 30753 18196 30787
rect 18144 30744 18196 30753
rect 15936 30676 15988 30685
rect 16488 30676 16540 30728
rect 17316 30676 17368 30728
rect 18052 30719 18104 30728
rect 18052 30685 18061 30719
rect 18061 30685 18095 30719
rect 18095 30685 18104 30719
rect 18052 30676 18104 30685
rect 18512 30676 18564 30728
rect 21272 30812 21324 30864
rect 22744 30744 22796 30796
rect 23848 30812 23900 30864
rect 24768 30787 24820 30796
rect 24768 30753 24777 30787
rect 24777 30753 24811 30787
rect 24811 30753 24820 30787
rect 24768 30744 24820 30753
rect 20720 30719 20772 30728
rect 20720 30685 20729 30719
rect 20729 30685 20763 30719
rect 20763 30685 20772 30719
rect 20720 30676 20772 30685
rect 20904 30719 20956 30728
rect 20904 30685 20913 30719
rect 20913 30685 20947 30719
rect 20947 30685 20956 30719
rect 20904 30676 20956 30685
rect 23112 30676 23164 30728
rect 27160 30812 27212 30864
rect 30472 30812 30524 30864
rect 25780 30719 25832 30728
rect 8024 30608 8076 30660
rect 24308 30608 24360 30660
rect 25780 30685 25789 30719
rect 25789 30685 25823 30719
rect 25823 30685 25832 30719
rect 25780 30676 25832 30685
rect 27436 30719 27488 30728
rect 27436 30685 27445 30719
rect 27445 30685 27479 30719
rect 27479 30685 27488 30719
rect 27436 30676 27488 30685
rect 25596 30608 25648 30660
rect 26424 30651 26476 30660
rect 26424 30617 26433 30651
rect 26433 30617 26467 30651
rect 26467 30617 26476 30651
rect 26424 30608 26476 30617
rect 19340 30583 19392 30592
rect 19340 30549 19349 30583
rect 19349 30549 19383 30583
rect 19383 30549 19392 30583
rect 19340 30540 19392 30549
rect 25412 30540 25464 30592
rect 27068 30583 27120 30592
rect 27068 30549 27077 30583
rect 27077 30549 27111 30583
rect 27111 30549 27120 30583
rect 27068 30540 27120 30549
rect 30656 30719 30708 30728
rect 30656 30685 30665 30719
rect 30665 30685 30699 30719
rect 30699 30685 30708 30719
rect 30656 30676 30708 30685
rect 30840 30676 30892 30728
rect 31024 30676 31076 30728
rect 31852 30812 31904 30864
rect 28172 30608 28224 30660
rect 30012 30608 30064 30660
rect 31668 30608 31720 30660
rect 31852 30682 31864 30706
rect 31864 30682 31898 30706
rect 31898 30682 31904 30706
rect 31852 30654 31904 30682
rect 32772 30719 32824 30728
rect 32772 30685 32781 30719
rect 32781 30685 32815 30719
rect 32815 30685 32824 30719
rect 32772 30676 32824 30685
rect 35992 30719 36044 30728
rect 35992 30685 36001 30719
rect 36001 30685 36035 30719
rect 36035 30685 36044 30719
rect 35992 30676 36044 30685
rect 36636 30676 36688 30728
rect 43720 30651 43772 30660
rect 43720 30617 43729 30651
rect 43729 30617 43763 30651
rect 43763 30617 43772 30651
rect 43720 30608 43772 30617
rect 44088 30651 44140 30660
rect 44088 30617 44097 30651
rect 44097 30617 44131 30651
rect 44131 30617 44140 30651
rect 44088 30608 44140 30617
rect 28816 30540 28868 30592
rect 30840 30540 30892 30592
rect 33692 30540 33744 30592
rect 33876 30540 33928 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 26332 30379 26384 30388
rect 26332 30345 26341 30379
rect 26341 30345 26375 30379
rect 26375 30345 26384 30379
rect 26332 30336 26384 30345
rect 30472 30379 30524 30388
rect 30472 30345 30481 30379
rect 30481 30345 30515 30379
rect 30515 30345 30524 30379
rect 30472 30336 30524 30345
rect 16672 30268 16724 30320
rect 17592 30268 17644 30320
rect 1768 30243 1820 30252
rect 1768 30209 1777 30243
rect 1777 30209 1811 30243
rect 1811 30209 1820 30243
rect 1768 30200 1820 30209
rect 16764 30200 16816 30252
rect 2228 30132 2280 30184
rect 2780 30175 2832 30184
rect 2780 30141 2789 30175
rect 2789 30141 2823 30175
rect 2823 30141 2832 30175
rect 2780 30132 2832 30141
rect 15844 30132 15896 30184
rect 17316 30107 17368 30116
rect 17316 30073 17325 30107
rect 17325 30073 17359 30107
rect 17359 30073 17368 30107
rect 17316 30064 17368 30073
rect 17684 29996 17736 30048
rect 18236 30243 18288 30252
rect 18236 30209 18245 30243
rect 18245 30209 18279 30243
rect 18279 30209 18288 30243
rect 18236 30200 18288 30209
rect 19340 30268 19392 30320
rect 22100 30268 22152 30320
rect 19248 30200 19300 30252
rect 20444 30200 20496 30252
rect 19064 30132 19116 30184
rect 24308 30243 24360 30252
rect 24308 30209 24317 30243
rect 24317 30209 24351 30243
rect 24351 30209 24360 30243
rect 24308 30200 24360 30209
rect 24768 30200 24820 30252
rect 25228 30200 25280 30252
rect 25780 30268 25832 30320
rect 27068 30268 27120 30320
rect 28080 30311 28132 30320
rect 28080 30277 28114 30311
rect 28114 30277 28132 30311
rect 28080 30268 28132 30277
rect 34796 30268 34848 30320
rect 24860 30064 24912 30116
rect 26516 30200 26568 30252
rect 29000 30200 29052 30252
rect 30012 30243 30064 30252
rect 30012 30209 30021 30243
rect 30021 30209 30055 30243
rect 30055 30209 30064 30243
rect 30012 30200 30064 30209
rect 30656 30200 30708 30252
rect 30932 30243 30984 30252
rect 30932 30209 30941 30243
rect 30941 30209 30975 30243
rect 30975 30209 30984 30243
rect 30932 30200 30984 30209
rect 25688 30132 25740 30184
rect 31208 30243 31260 30252
rect 31208 30209 31217 30243
rect 31217 30209 31251 30243
rect 31251 30209 31260 30243
rect 31208 30200 31260 30209
rect 31484 30200 31536 30252
rect 31852 30200 31904 30252
rect 32312 30243 32364 30252
rect 32312 30209 32321 30243
rect 32321 30209 32355 30243
rect 32355 30209 32364 30243
rect 32312 30200 32364 30209
rect 34520 30200 34572 30252
rect 37464 30243 37516 30252
rect 37464 30209 37473 30243
rect 37473 30209 37507 30243
rect 37507 30209 37516 30243
rect 37464 30200 37516 30209
rect 43352 30243 43404 30252
rect 43352 30209 43361 30243
rect 43361 30209 43395 30243
rect 43395 30209 43404 30243
rect 43352 30200 43404 30209
rect 32772 30175 32824 30184
rect 25596 30064 25648 30116
rect 32772 30141 32781 30175
rect 32781 30141 32815 30175
rect 32815 30141 32824 30175
rect 32772 30132 32824 30141
rect 33876 30132 33928 30184
rect 35992 30064 36044 30116
rect 37188 30064 37240 30116
rect 24676 30039 24728 30048
rect 24676 30005 24685 30039
rect 24685 30005 24719 30039
rect 24719 30005 24728 30039
rect 24676 29996 24728 30005
rect 25412 29996 25464 30048
rect 26056 29996 26108 30048
rect 28908 29996 28960 30048
rect 29552 29996 29604 30048
rect 30472 29996 30524 30048
rect 33968 29996 34020 30048
rect 36820 29996 36872 30048
rect 43996 29996 44048 30048
rect 44180 30039 44232 30048
rect 44180 30005 44189 30039
rect 44189 30005 44223 30039
rect 44223 30005 44232 30039
rect 44180 29996 44232 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 2228 29835 2280 29844
rect 2228 29801 2237 29835
rect 2237 29801 2271 29835
rect 2271 29801 2280 29835
rect 2228 29792 2280 29801
rect 15844 29835 15896 29844
rect 15844 29801 15853 29835
rect 15853 29801 15887 29835
rect 15887 29801 15896 29835
rect 15844 29792 15896 29801
rect 16764 29835 16816 29844
rect 16764 29801 16773 29835
rect 16773 29801 16807 29835
rect 16807 29801 16816 29835
rect 16764 29792 16816 29801
rect 18052 29792 18104 29844
rect 19248 29835 19300 29844
rect 19248 29801 19257 29835
rect 19257 29801 19291 29835
rect 19291 29801 19300 29835
rect 19248 29792 19300 29801
rect 19984 29792 20036 29844
rect 21456 29792 21508 29844
rect 24676 29792 24728 29844
rect 28264 29835 28316 29844
rect 28264 29801 28273 29835
rect 28273 29801 28307 29835
rect 28307 29801 28316 29835
rect 28264 29792 28316 29801
rect 28816 29835 28868 29844
rect 28816 29801 28825 29835
rect 28825 29801 28859 29835
rect 28859 29801 28868 29835
rect 28816 29792 28868 29801
rect 31300 29792 31352 29844
rect 31392 29792 31444 29844
rect 33600 29792 33652 29844
rect 28540 29724 28592 29776
rect 15568 29656 15620 29708
rect 2412 29588 2464 29640
rect 14464 29631 14516 29640
rect 14464 29597 14473 29631
rect 14473 29597 14507 29631
rect 14507 29597 14516 29631
rect 14464 29588 14516 29597
rect 16488 29656 16540 29708
rect 17684 29699 17736 29708
rect 17684 29665 17693 29699
rect 17693 29665 17727 29699
rect 17727 29665 17736 29699
rect 17684 29656 17736 29665
rect 17592 29631 17644 29640
rect 17592 29597 17601 29631
rect 17601 29597 17635 29631
rect 17635 29597 17644 29631
rect 17592 29588 17644 29597
rect 17868 29631 17920 29640
rect 17868 29597 17877 29631
rect 17877 29597 17911 29631
rect 17911 29597 17920 29631
rect 17868 29588 17920 29597
rect 16396 29563 16448 29572
rect 16396 29529 16405 29563
rect 16405 29529 16439 29563
rect 16439 29529 16448 29563
rect 16396 29520 16448 29529
rect 14188 29452 14240 29504
rect 17408 29452 17460 29504
rect 18328 29588 18380 29640
rect 30656 29656 30708 29708
rect 31852 29656 31904 29708
rect 20444 29631 20496 29640
rect 20444 29597 20453 29631
rect 20453 29597 20487 29631
rect 20487 29597 20496 29631
rect 20444 29588 20496 29597
rect 25688 29631 25740 29640
rect 25688 29597 25697 29631
rect 25697 29597 25731 29631
rect 25731 29597 25740 29631
rect 25688 29588 25740 29597
rect 25964 29631 26016 29640
rect 25964 29597 25998 29631
rect 25998 29597 26016 29631
rect 25964 29588 26016 29597
rect 27712 29588 27764 29640
rect 28908 29631 28960 29640
rect 28908 29597 28917 29631
rect 28917 29597 28951 29631
rect 28951 29597 28960 29631
rect 28908 29588 28960 29597
rect 30472 29631 30524 29640
rect 30472 29597 30481 29631
rect 30481 29597 30515 29631
rect 30515 29597 30524 29631
rect 30472 29588 30524 29597
rect 30564 29631 30616 29640
rect 30564 29597 30573 29631
rect 30573 29597 30607 29631
rect 30607 29597 30616 29631
rect 30564 29588 30616 29597
rect 31024 29588 31076 29640
rect 34796 29588 34848 29640
rect 43352 29792 43404 29844
rect 42708 29699 42760 29708
rect 42708 29665 42717 29699
rect 42717 29665 42751 29699
rect 42751 29665 42760 29699
rect 42708 29656 42760 29665
rect 43996 29699 44048 29708
rect 43996 29665 44005 29699
rect 44005 29665 44039 29699
rect 44039 29665 44048 29699
rect 43996 29656 44048 29665
rect 44180 29699 44232 29708
rect 44180 29665 44189 29699
rect 44189 29665 44223 29699
rect 44223 29665 44232 29699
rect 44180 29656 44232 29665
rect 36820 29588 36872 29640
rect 37188 29588 37240 29640
rect 18420 29520 18472 29572
rect 18972 29520 19024 29572
rect 25228 29520 25280 29572
rect 26424 29520 26476 29572
rect 30380 29520 30432 29572
rect 33324 29563 33376 29572
rect 33324 29529 33333 29563
rect 33333 29529 33367 29563
rect 33367 29529 33376 29563
rect 33324 29520 33376 29529
rect 33876 29520 33928 29572
rect 35624 29520 35676 29572
rect 27436 29452 27488 29504
rect 32772 29452 32824 29504
rect 33232 29452 33284 29504
rect 33692 29452 33744 29504
rect 35808 29452 35860 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 13912 29248 13964 29300
rect 17960 29248 18012 29300
rect 18144 29248 18196 29300
rect 18972 29248 19024 29300
rect 19432 29248 19484 29300
rect 29552 29291 29604 29300
rect 14280 29180 14332 29232
rect 14188 29112 14240 29164
rect 17040 29155 17092 29164
rect 17040 29121 17049 29155
rect 17049 29121 17083 29155
rect 17083 29121 17092 29155
rect 17040 29112 17092 29121
rect 19340 29180 19392 29232
rect 21272 29180 21324 29232
rect 24584 29223 24636 29232
rect 24584 29189 24593 29223
rect 24593 29189 24627 29223
rect 24627 29189 24636 29223
rect 24584 29180 24636 29189
rect 25320 29180 25372 29232
rect 29552 29257 29561 29291
rect 29561 29257 29595 29291
rect 29595 29257 29604 29291
rect 29552 29248 29604 29257
rect 30472 29248 30524 29300
rect 32312 29248 32364 29300
rect 43720 29248 43772 29300
rect 35992 29223 36044 29232
rect 35992 29189 36001 29223
rect 36001 29189 36035 29223
rect 36035 29189 36044 29223
rect 35992 29180 36044 29189
rect 18420 29155 18472 29164
rect 17316 29087 17368 29096
rect 17316 29053 17325 29087
rect 17325 29053 17359 29087
rect 17359 29053 17368 29087
rect 17316 29044 17368 29053
rect 18420 29121 18429 29155
rect 18429 29121 18463 29155
rect 18463 29121 18472 29155
rect 18420 29112 18472 29121
rect 18880 29155 18932 29164
rect 18880 29121 18889 29155
rect 18889 29121 18923 29155
rect 18923 29121 18932 29155
rect 18880 29112 18932 29121
rect 19064 29155 19116 29164
rect 19064 29121 19073 29155
rect 19073 29121 19107 29155
rect 19107 29121 19116 29155
rect 19064 29112 19116 29121
rect 20444 29112 20496 29164
rect 21732 29112 21784 29164
rect 28908 29112 28960 29164
rect 18236 29044 18288 29096
rect 19248 29044 19300 29096
rect 21824 29087 21876 29096
rect 21824 29053 21833 29087
rect 21833 29053 21867 29087
rect 21867 29053 21876 29087
rect 21824 29044 21876 29053
rect 15200 28976 15252 29028
rect 16672 28976 16724 29028
rect 17868 28976 17920 29028
rect 18328 29019 18380 29028
rect 18328 28985 18337 29019
rect 18337 28985 18371 29019
rect 18371 28985 18380 29019
rect 18328 28976 18380 28985
rect 20536 28976 20588 29028
rect 20904 28976 20956 29028
rect 24216 29019 24268 29028
rect 24216 28985 24225 29019
rect 24225 28985 24259 29019
rect 24259 28985 24268 29019
rect 24216 28976 24268 28985
rect 24860 28976 24912 29028
rect 30472 29112 30524 29164
rect 31484 29112 31536 29164
rect 31668 29112 31720 29164
rect 32588 29112 32640 29164
rect 33324 29112 33376 29164
rect 33876 29155 33928 29164
rect 33876 29121 33885 29155
rect 33885 29121 33919 29155
rect 33919 29121 33928 29155
rect 33876 29112 33928 29121
rect 33968 29155 34020 29164
rect 33968 29121 33977 29155
rect 33977 29121 34011 29155
rect 34011 29121 34020 29155
rect 33968 29112 34020 29121
rect 35532 29112 35584 29164
rect 35808 29155 35860 29164
rect 35808 29121 35817 29155
rect 35817 29121 35851 29155
rect 35851 29121 35860 29155
rect 35808 29112 35860 29121
rect 28724 29019 28776 29028
rect 28724 28985 28733 29019
rect 28733 28985 28767 29019
rect 28767 28985 28776 29019
rect 28724 28976 28776 28985
rect 30380 29019 30432 29028
rect 17224 28951 17276 28960
rect 17224 28917 17233 28951
rect 17233 28917 17267 28951
rect 17267 28917 17276 28951
rect 17224 28908 17276 28917
rect 23204 28951 23256 28960
rect 23204 28917 23213 28951
rect 23213 28917 23247 28951
rect 23247 28917 23256 28951
rect 23204 28908 23256 28917
rect 25412 28951 25464 28960
rect 25412 28917 25421 28951
rect 25421 28917 25455 28951
rect 25455 28917 25464 28951
rect 25412 28908 25464 28917
rect 30380 28985 30389 29019
rect 30389 28985 30423 29019
rect 30423 28985 30432 29019
rect 30380 28976 30432 28985
rect 30472 28908 30524 28960
rect 30748 29044 30800 29096
rect 31300 29087 31352 29096
rect 31300 29053 31309 29087
rect 31309 29053 31343 29087
rect 31343 29053 31352 29087
rect 31300 29044 31352 29053
rect 33232 29044 33284 29096
rect 31576 28976 31628 29028
rect 32588 28976 32640 29028
rect 33968 28976 34020 29028
rect 34796 28976 34848 29028
rect 32128 28951 32180 28960
rect 32128 28917 32137 28951
rect 32137 28917 32171 28951
rect 32171 28917 32180 28951
rect 32128 28908 32180 28917
rect 32312 28908 32364 28960
rect 33692 28908 33744 28960
rect 35716 28908 35768 28960
rect 36544 28951 36596 28960
rect 36544 28917 36553 28951
rect 36553 28917 36587 28951
rect 36587 28917 36596 28951
rect 36544 28908 36596 28917
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 15200 28704 15252 28756
rect 16488 28704 16540 28756
rect 21272 28747 21324 28756
rect 16396 28636 16448 28688
rect 17316 28636 17368 28688
rect 16856 28568 16908 28620
rect 17224 28568 17276 28620
rect 14280 28543 14332 28552
rect 14280 28509 14289 28543
rect 14289 28509 14323 28543
rect 14323 28509 14332 28543
rect 14280 28500 14332 28509
rect 16580 28543 16632 28552
rect 16580 28509 16589 28543
rect 16589 28509 16623 28543
rect 16623 28509 16632 28543
rect 17500 28543 17552 28552
rect 16580 28500 16632 28509
rect 17500 28509 17509 28543
rect 17509 28509 17543 28543
rect 17543 28509 17552 28543
rect 17500 28500 17552 28509
rect 21272 28713 21281 28747
rect 21281 28713 21315 28747
rect 21315 28713 21324 28747
rect 21272 28704 21324 28713
rect 22192 28704 22244 28756
rect 27712 28747 27764 28756
rect 27712 28713 27721 28747
rect 27721 28713 27755 28747
rect 27755 28713 27764 28747
rect 27712 28704 27764 28713
rect 27896 28747 27948 28756
rect 27896 28713 27905 28747
rect 27905 28713 27939 28747
rect 27939 28713 27948 28747
rect 27896 28704 27948 28713
rect 30472 28704 30524 28756
rect 31300 28704 31352 28756
rect 31668 28704 31720 28756
rect 35532 28704 35584 28756
rect 35716 28747 35768 28756
rect 35716 28713 35725 28747
rect 35725 28713 35759 28747
rect 35759 28713 35768 28747
rect 35716 28704 35768 28713
rect 37464 28704 37516 28756
rect 25412 28636 25464 28688
rect 25780 28679 25832 28688
rect 25780 28645 25789 28679
rect 25789 28645 25823 28679
rect 25823 28645 25832 28679
rect 25780 28636 25832 28645
rect 34888 28636 34940 28688
rect 19064 28568 19116 28620
rect 22652 28568 22704 28620
rect 18328 28500 18380 28552
rect 21824 28500 21876 28552
rect 22284 28543 22336 28552
rect 22284 28509 22293 28543
rect 22293 28509 22327 28543
rect 22327 28509 22336 28543
rect 22284 28500 22336 28509
rect 23020 28543 23072 28552
rect 20720 28432 20772 28484
rect 23020 28509 23029 28543
rect 23029 28509 23063 28543
rect 23063 28509 23072 28543
rect 23020 28500 23072 28509
rect 24216 28568 24268 28620
rect 24860 28568 24912 28620
rect 27988 28568 28040 28620
rect 28540 28568 28592 28620
rect 23296 28500 23348 28552
rect 26056 28500 26108 28552
rect 27068 28543 27120 28552
rect 27068 28509 27077 28543
rect 27077 28509 27111 28543
rect 27111 28509 27120 28543
rect 27068 28500 27120 28509
rect 27344 28500 27396 28552
rect 30748 28568 30800 28620
rect 31208 28568 31260 28620
rect 32128 28568 32180 28620
rect 33600 28611 33652 28620
rect 33600 28577 33609 28611
rect 33609 28577 33643 28611
rect 33643 28577 33652 28611
rect 33600 28568 33652 28577
rect 34796 28568 34848 28620
rect 30564 28500 30616 28552
rect 31576 28500 31628 28552
rect 16120 28407 16172 28416
rect 16120 28373 16129 28407
rect 16129 28373 16163 28407
rect 16163 28373 16172 28407
rect 16120 28364 16172 28373
rect 18052 28364 18104 28416
rect 21640 28364 21692 28416
rect 21916 28407 21968 28416
rect 21916 28373 21925 28407
rect 21925 28373 21959 28407
rect 21959 28373 21968 28407
rect 21916 28364 21968 28373
rect 23388 28364 23440 28416
rect 27528 28364 27580 28416
rect 27988 28432 28040 28484
rect 28908 28432 28960 28484
rect 31760 28432 31812 28484
rect 31944 28432 31996 28484
rect 32312 28543 32364 28552
rect 32312 28509 32321 28543
rect 32321 28509 32355 28543
rect 32355 28509 32364 28543
rect 33324 28543 33376 28552
rect 32312 28500 32364 28509
rect 33324 28509 33333 28543
rect 33333 28509 33367 28543
rect 33367 28509 33376 28543
rect 33324 28500 33376 28509
rect 34520 28432 34572 28484
rect 37188 28500 37240 28552
rect 43444 28543 43496 28552
rect 43444 28509 43453 28543
rect 43453 28509 43487 28543
rect 43487 28509 43496 28543
rect 43444 28500 43496 28509
rect 35532 28475 35584 28484
rect 28172 28364 28224 28416
rect 31024 28364 31076 28416
rect 31116 28364 31168 28416
rect 32496 28364 32548 28416
rect 32588 28364 32640 28416
rect 34428 28364 34480 28416
rect 35532 28441 35541 28475
rect 35541 28441 35575 28475
rect 35575 28441 35584 28475
rect 35532 28432 35584 28441
rect 36084 28432 36136 28484
rect 36544 28432 36596 28484
rect 36728 28475 36780 28484
rect 36728 28441 36762 28475
rect 36762 28441 36780 28475
rect 36728 28432 36780 28441
rect 36176 28364 36228 28416
rect 37464 28364 37516 28416
rect 43996 28364 44048 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 14464 28160 14516 28212
rect 17868 28160 17920 28212
rect 21272 28160 21324 28212
rect 22192 28203 22244 28212
rect 22192 28169 22201 28203
rect 22201 28169 22235 28203
rect 22235 28169 22244 28203
rect 22192 28160 22244 28169
rect 17040 28092 17092 28144
rect 16028 28024 16080 28076
rect 16856 28024 16908 28076
rect 15200 27999 15252 28008
rect 15200 27965 15209 27999
rect 15209 27965 15243 27999
rect 15243 27965 15252 27999
rect 15200 27956 15252 27965
rect 17684 28024 17736 28076
rect 18052 28067 18104 28076
rect 18052 28033 18061 28067
rect 18061 28033 18095 28067
rect 18095 28033 18104 28067
rect 18052 28024 18104 28033
rect 19432 28024 19484 28076
rect 21916 28092 21968 28144
rect 22284 28024 22336 28076
rect 23204 28160 23256 28212
rect 24216 28160 24268 28212
rect 27344 28203 27396 28212
rect 22744 28092 22796 28144
rect 22652 28067 22704 28076
rect 22652 28033 22661 28067
rect 22661 28033 22695 28067
rect 22695 28033 22704 28067
rect 25688 28092 25740 28144
rect 22652 28024 22704 28033
rect 23388 28067 23440 28076
rect 23388 28033 23422 28067
rect 23422 28033 23440 28067
rect 23388 28024 23440 28033
rect 27344 28169 27353 28203
rect 27353 28169 27387 28203
rect 27387 28169 27396 28203
rect 27344 28160 27396 28169
rect 27528 28203 27580 28212
rect 27528 28169 27537 28203
rect 27537 28169 27571 28203
rect 27571 28169 27580 28203
rect 27528 28160 27580 28169
rect 31208 28160 31260 28212
rect 27068 28024 27120 28076
rect 28540 28067 28592 28076
rect 28540 28033 28549 28067
rect 28549 28033 28583 28067
rect 28583 28033 28592 28067
rect 28540 28024 28592 28033
rect 29552 28067 29604 28076
rect 29552 28033 29561 28067
rect 29561 28033 29595 28067
rect 29595 28033 29604 28067
rect 29552 28024 29604 28033
rect 17960 27888 18012 27940
rect 26056 27956 26108 28008
rect 24860 27888 24912 27940
rect 27712 27956 27764 28008
rect 27988 27956 28040 28008
rect 30564 28024 30616 28076
rect 31300 28067 31352 28076
rect 31300 28033 31309 28067
rect 31309 28033 31343 28067
rect 31343 28033 31352 28067
rect 31300 28024 31352 28033
rect 32588 28160 32640 28212
rect 33324 28160 33376 28212
rect 36084 28160 36136 28212
rect 36728 28203 36780 28212
rect 36728 28169 36737 28203
rect 36737 28169 36771 28203
rect 36771 28169 36780 28203
rect 36728 28160 36780 28169
rect 32772 28092 32824 28144
rect 34060 28092 34112 28144
rect 32680 28067 32732 28076
rect 32680 28033 32714 28067
rect 32714 28033 32732 28067
rect 34428 28067 34480 28076
rect 32680 28024 32732 28033
rect 34428 28033 34437 28067
rect 34437 28033 34471 28067
rect 34471 28033 34480 28067
rect 34428 28024 34480 28033
rect 35532 28024 35584 28076
rect 36268 28067 36320 28076
rect 36268 28033 36277 28067
rect 36277 28033 36311 28067
rect 36311 28033 36320 28067
rect 36268 28024 36320 28033
rect 37464 28067 37516 28076
rect 30748 27956 30800 28008
rect 33600 27956 33652 28008
rect 16764 27820 16816 27872
rect 18328 27820 18380 27872
rect 20904 27820 20956 27872
rect 25320 27863 25372 27872
rect 25320 27829 25329 27863
rect 25329 27829 25363 27863
rect 25363 27829 25372 27863
rect 25320 27820 25372 27829
rect 26608 27820 26660 27872
rect 30656 27888 30708 27940
rect 31024 27931 31076 27940
rect 31024 27897 31033 27931
rect 31033 27897 31067 27931
rect 31067 27897 31076 27931
rect 31024 27888 31076 27897
rect 29828 27820 29880 27872
rect 31852 27820 31904 27872
rect 36176 27820 36228 27872
rect 37464 28033 37473 28067
rect 37473 28033 37507 28067
rect 37507 28033 37516 28067
rect 37464 28024 37516 28033
rect 44180 27820 44232 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 16120 27616 16172 27668
rect 16580 27616 16632 27668
rect 17960 27616 18012 27668
rect 22284 27616 22336 27668
rect 16672 27591 16724 27600
rect 16672 27557 16681 27591
rect 16681 27557 16715 27591
rect 16715 27557 16724 27591
rect 16672 27548 16724 27557
rect 18328 27548 18380 27600
rect 20720 27591 20772 27600
rect 20720 27557 20729 27591
rect 20729 27557 20763 27591
rect 20763 27557 20772 27591
rect 20720 27548 20772 27557
rect 21732 27548 21784 27600
rect 23020 27616 23072 27668
rect 22744 27548 22796 27600
rect 17868 27480 17920 27532
rect 21272 27480 21324 27532
rect 27896 27616 27948 27668
rect 30656 27616 30708 27668
rect 31116 27616 31168 27668
rect 32680 27659 32732 27668
rect 32680 27625 32689 27659
rect 32689 27625 32723 27659
rect 32723 27625 32732 27659
rect 32680 27616 32732 27625
rect 36268 27616 36320 27668
rect 30380 27548 30432 27600
rect 31852 27591 31904 27600
rect 31852 27557 31861 27591
rect 31861 27557 31895 27591
rect 31895 27557 31904 27591
rect 31852 27548 31904 27557
rect 25688 27523 25740 27532
rect 25688 27489 25697 27523
rect 25697 27489 25731 27523
rect 25731 27489 25740 27523
rect 25688 27480 25740 27489
rect 29000 27480 29052 27532
rect 29828 27523 29880 27532
rect 29828 27489 29837 27523
rect 29837 27489 29871 27523
rect 29871 27489 29880 27523
rect 29828 27480 29880 27489
rect 42708 27523 42760 27532
rect 42708 27489 42717 27523
rect 42717 27489 42751 27523
rect 42751 27489 42760 27523
rect 42708 27480 42760 27489
rect 43996 27523 44048 27532
rect 43996 27489 44005 27523
rect 44005 27489 44039 27523
rect 44039 27489 44048 27523
rect 43996 27480 44048 27489
rect 44180 27523 44232 27532
rect 44180 27489 44189 27523
rect 44189 27489 44223 27523
rect 44223 27489 44232 27523
rect 44180 27480 44232 27489
rect 16672 27412 16724 27464
rect 16856 27412 16908 27464
rect 17684 27412 17736 27464
rect 17960 27412 18012 27464
rect 20904 27455 20956 27464
rect 20904 27421 20913 27455
rect 20913 27421 20947 27455
rect 20947 27421 20956 27455
rect 20904 27412 20956 27421
rect 21640 27455 21692 27464
rect 21640 27421 21649 27455
rect 21649 27421 21683 27455
rect 21683 27421 21692 27455
rect 21640 27412 21692 27421
rect 23112 27412 23164 27464
rect 23296 27455 23348 27464
rect 23296 27421 23305 27455
rect 23305 27421 23339 27455
rect 23339 27421 23348 27455
rect 23296 27412 23348 27421
rect 23388 27412 23440 27464
rect 24584 27412 24636 27464
rect 28172 27412 28224 27464
rect 30840 27455 30892 27464
rect 30840 27421 30849 27455
rect 30849 27421 30883 27455
rect 30883 27421 30892 27455
rect 30840 27412 30892 27421
rect 31852 27455 31904 27464
rect 31852 27421 31861 27455
rect 31861 27421 31895 27455
rect 31895 27421 31904 27455
rect 31852 27412 31904 27421
rect 32036 27455 32088 27464
rect 32036 27421 32045 27455
rect 32045 27421 32079 27455
rect 32079 27421 32088 27455
rect 32036 27412 32088 27421
rect 32496 27455 32548 27464
rect 32496 27421 32505 27455
rect 32505 27421 32539 27455
rect 32539 27421 32548 27455
rect 32496 27412 32548 27421
rect 34704 27455 34756 27464
rect 34704 27421 34713 27455
rect 34713 27421 34747 27455
rect 34747 27421 34756 27455
rect 34704 27412 34756 27421
rect 36084 27455 36136 27464
rect 20168 27344 20220 27396
rect 20628 27344 20680 27396
rect 23204 27344 23256 27396
rect 25320 27344 25372 27396
rect 34612 27344 34664 27396
rect 36084 27421 36093 27455
rect 36093 27421 36127 27455
rect 36127 27421 36136 27455
rect 36084 27412 36136 27421
rect 36176 27412 36228 27464
rect 17592 27276 17644 27328
rect 22652 27319 22704 27328
rect 22652 27285 22679 27319
rect 22679 27285 22704 27319
rect 22652 27276 22704 27285
rect 23388 27276 23440 27328
rect 25136 27319 25188 27328
rect 25136 27285 25145 27319
rect 25145 27285 25179 27319
rect 25179 27285 25188 27319
rect 25136 27276 25188 27285
rect 28908 27276 28960 27328
rect 31116 27276 31168 27328
rect 33508 27276 33560 27328
rect 34428 27276 34480 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 16856 27072 16908 27124
rect 28724 27072 28776 27124
rect 29000 27115 29052 27124
rect 29000 27081 29009 27115
rect 29009 27081 29043 27115
rect 29043 27081 29052 27115
rect 29000 27072 29052 27081
rect 16672 27004 16724 27056
rect 17408 27047 17460 27056
rect 17408 27013 17417 27047
rect 17417 27013 17451 27047
rect 17451 27013 17460 27047
rect 17408 27004 17460 27013
rect 24032 27004 24084 27056
rect 28540 27004 28592 27056
rect 32956 27004 33008 27056
rect 34152 27004 34204 27056
rect 14280 26936 14332 26988
rect 15476 26936 15528 26988
rect 17592 26979 17644 26988
rect 17592 26945 17601 26979
rect 17601 26945 17635 26979
rect 17635 26945 17644 26979
rect 17592 26936 17644 26945
rect 17868 26936 17920 26988
rect 17776 26868 17828 26920
rect 23296 26936 23348 26988
rect 23480 26868 23532 26920
rect 28816 26979 28868 26988
rect 28816 26945 28825 26979
rect 28825 26945 28859 26979
rect 28859 26945 28868 26979
rect 28816 26936 28868 26945
rect 30840 26936 30892 26988
rect 33600 26979 33652 26988
rect 33600 26945 33609 26979
rect 33609 26945 33643 26979
rect 33643 26945 33652 26979
rect 33600 26936 33652 26945
rect 33968 26936 34020 26988
rect 34244 26979 34296 26988
rect 34244 26945 34253 26979
rect 34253 26945 34287 26979
rect 34287 26945 34296 26979
rect 34244 26936 34296 26945
rect 34428 26979 34480 26988
rect 34428 26945 34437 26979
rect 34437 26945 34471 26979
rect 34471 26945 34480 26979
rect 34428 26936 34480 26945
rect 34704 27004 34756 27056
rect 34612 26979 34664 26988
rect 34612 26945 34621 26979
rect 34621 26945 34655 26979
rect 34655 26945 34664 26979
rect 34612 26936 34664 26945
rect 28908 26868 28960 26920
rect 31300 26868 31352 26920
rect 37188 26868 37240 26920
rect 27528 26800 27580 26852
rect 28540 26800 28592 26852
rect 29552 26800 29604 26852
rect 31852 26800 31904 26852
rect 16212 26732 16264 26784
rect 23020 26775 23072 26784
rect 23020 26741 23029 26775
rect 23029 26741 23063 26775
rect 23063 26741 23072 26775
rect 23020 26732 23072 26741
rect 35348 26775 35400 26784
rect 35348 26741 35357 26775
rect 35357 26741 35391 26775
rect 35391 26741 35400 26775
rect 35348 26732 35400 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 15476 26571 15528 26580
rect 15476 26537 15485 26571
rect 15485 26537 15519 26571
rect 15519 26537 15528 26571
rect 15476 26528 15528 26537
rect 17408 26528 17460 26580
rect 17684 26528 17736 26580
rect 28816 26528 28868 26580
rect 31852 26528 31904 26580
rect 34612 26528 34664 26580
rect 34704 26528 34756 26580
rect 16120 26460 16172 26512
rect 19984 26460 20036 26512
rect 17868 26392 17920 26444
rect 16212 26324 16264 26376
rect 16764 26367 16816 26376
rect 16764 26333 16773 26367
rect 16773 26333 16807 26367
rect 16807 26333 16816 26367
rect 16764 26324 16816 26333
rect 17040 26256 17092 26308
rect 17960 26324 18012 26376
rect 18328 26367 18380 26376
rect 18328 26333 18337 26367
rect 18337 26333 18371 26367
rect 18371 26333 18380 26367
rect 19248 26367 19300 26376
rect 18328 26324 18380 26333
rect 19248 26333 19257 26367
rect 19257 26333 19291 26367
rect 19291 26333 19300 26367
rect 19248 26324 19300 26333
rect 22376 26460 22428 26512
rect 23756 26460 23808 26512
rect 26792 26460 26844 26512
rect 31024 26503 31076 26512
rect 31024 26469 31033 26503
rect 31033 26469 31067 26503
rect 31067 26469 31076 26503
rect 31024 26460 31076 26469
rect 32036 26460 32088 26512
rect 35348 26460 35400 26512
rect 22100 26367 22152 26376
rect 22100 26333 22123 26367
rect 22123 26333 22152 26367
rect 22100 26324 22152 26333
rect 22284 26367 22336 26376
rect 22284 26333 22293 26367
rect 22293 26333 22327 26367
rect 22327 26333 22336 26367
rect 22284 26324 22336 26333
rect 22928 26324 22980 26376
rect 23388 26324 23440 26376
rect 24492 26324 24544 26376
rect 25504 26367 25556 26376
rect 25504 26333 25513 26367
rect 25513 26333 25547 26367
rect 25547 26333 25556 26367
rect 25504 26324 25556 26333
rect 27896 26324 27948 26376
rect 33324 26392 33376 26444
rect 31484 26324 31536 26376
rect 32128 26367 32180 26376
rect 32128 26333 32137 26367
rect 32137 26333 32171 26367
rect 32171 26333 32180 26367
rect 32128 26324 32180 26333
rect 33600 26367 33652 26376
rect 5172 26188 5224 26240
rect 16580 26188 16632 26240
rect 18052 26231 18104 26240
rect 18052 26197 18061 26231
rect 18061 26197 18095 26231
rect 18095 26197 18104 26231
rect 18052 26188 18104 26197
rect 20812 26231 20864 26240
rect 20812 26197 20821 26231
rect 20821 26197 20855 26231
rect 20855 26197 20864 26231
rect 20812 26188 20864 26197
rect 20996 26188 21048 26240
rect 21272 26188 21324 26240
rect 23020 26256 23072 26308
rect 30288 26256 30340 26308
rect 31944 26256 31996 26308
rect 33600 26333 33609 26367
rect 33609 26333 33643 26367
rect 33643 26333 33652 26367
rect 33600 26324 33652 26333
rect 33784 26324 33836 26376
rect 34520 26324 34572 26376
rect 41420 26392 41472 26444
rect 37188 26367 37240 26376
rect 37188 26333 37197 26367
rect 37197 26333 37231 26367
rect 37231 26333 37240 26367
rect 37188 26324 37240 26333
rect 41604 26367 41656 26376
rect 41604 26333 41613 26367
rect 41613 26333 41647 26367
rect 41647 26333 41656 26367
rect 41604 26324 41656 26333
rect 43904 26367 43956 26376
rect 43904 26333 43913 26367
rect 43913 26333 43947 26367
rect 43947 26333 43956 26367
rect 43904 26324 43956 26333
rect 34244 26256 34296 26308
rect 35992 26256 36044 26308
rect 41788 26299 41840 26308
rect 41788 26265 41797 26299
rect 41797 26265 41831 26299
rect 41831 26265 41840 26299
rect 41788 26256 41840 26265
rect 22192 26188 22244 26240
rect 23480 26188 23532 26240
rect 24492 26188 24544 26240
rect 26332 26231 26384 26240
rect 26332 26197 26341 26231
rect 26341 26197 26375 26231
rect 26375 26197 26384 26231
rect 26332 26188 26384 26197
rect 29828 26188 29880 26240
rect 32956 26231 33008 26240
rect 32956 26197 32991 26231
rect 32991 26197 33008 26231
rect 32956 26188 33008 26197
rect 33324 26188 33376 26240
rect 33876 26188 33928 26240
rect 35716 26188 35768 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 16580 25984 16632 26036
rect 3332 25959 3384 25968
rect 3332 25925 3341 25959
rect 3341 25925 3375 25959
rect 3375 25925 3384 25959
rect 3332 25916 3384 25925
rect 15568 25916 15620 25968
rect 24032 25959 24084 25968
rect 5172 25891 5224 25900
rect 5172 25857 5181 25891
rect 5181 25857 5215 25891
rect 5215 25857 5224 25891
rect 15844 25891 15896 25900
rect 5172 25848 5224 25857
rect 15844 25857 15853 25891
rect 15853 25857 15887 25891
rect 15887 25857 15896 25891
rect 15844 25848 15896 25857
rect 3976 25780 4028 25832
rect 16672 25848 16724 25900
rect 17040 25891 17092 25900
rect 17040 25857 17049 25891
rect 17049 25857 17083 25891
rect 17083 25857 17092 25891
rect 17040 25848 17092 25857
rect 17960 25848 18012 25900
rect 18144 25891 18196 25900
rect 18144 25857 18178 25891
rect 18178 25857 18196 25891
rect 18144 25848 18196 25857
rect 19984 25891 20036 25900
rect 19984 25857 20018 25891
rect 20018 25857 20036 25891
rect 19984 25848 20036 25857
rect 22192 25891 22244 25900
rect 22192 25857 22226 25891
rect 22226 25857 22244 25891
rect 22192 25848 22244 25857
rect 24032 25925 24041 25959
rect 24041 25925 24075 25959
rect 24075 25925 24084 25959
rect 24032 25916 24084 25925
rect 24492 25959 24544 25968
rect 24492 25925 24501 25959
rect 24501 25925 24535 25959
rect 24535 25925 24544 25959
rect 24492 25916 24544 25925
rect 26332 25916 26384 25968
rect 23664 25848 23716 25900
rect 27068 25916 27120 25968
rect 30564 25984 30616 26036
rect 33784 25984 33836 26036
rect 34704 26027 34756 26036
rect 34704 25993 34713 26027
rect 34713 25993 34747 26027
rect 34747 25993 34756 26027
rect 34704 25984 34756 25993
rect 35992 26027 36044 26036
rect 32036 25916 32088 25968
rect 32128 25916 32180 25968
rect 33600 25916 33652 25968
rect 34612 25916 34664 25968
rect 35992 25993 36001 26027
rect 36001 25993 36035 26027
rect 36035 25993 36044 26027
rect 35992 25984 36044 25993
rect 41604 25984 41656 26036
rect 16764 25823 16816 25832
rect 16764 25789 16773 25823
rect 16773 25789 16807 25823
rect 16807 25789 16816 25823
rect 16764 25780 16816 25789
rect 19248 25755 19300 25764
rect 19248 25721 19257 25755
rect 19257 25721 19291 25755
rect 19291 25721 19300 25755
rect 19248 25712 19300 25721
rect 15844 25687 15896 25696
rect 15844 25653 15853 25687
rect 15853 25653 15887 25687
rect 15887 25653 15896 25687
rect 15844 25644 15896 25653
rect 20996 25644 21048 25696
rect 23296 25755 23348 25764
rect 23296 25721 23305 25755
rect 23305 25721 23339 25755
rect 23339 25721 23348 25755
rect 23296 25712 23348 25721
rect 26516 25712 26568 25764
rect 27620 25780 27672 25832
rect 23572 25644 23624 25696
rect 26148 25644 26200 25696
rect 28632 25712 28684 25764
rect 28908 25891 28960 25900
rect 28908 25857 28917 25891
rect 28917 25857 28951 25891
rect 28951 25857 28960 25891
rect 28908 25848 28960 25857
rect 31024 25848 31076 25900
rect 31760 25848 31812 25900
rect 33324 25891 33376 25900
rect 30472 25780 30524 25832
rect 33048 25780 33100 25832
rect 33324 25857 33333 25891
rect 33333 25857 33367 25891
rect 33367 25857 33376 25891
rect 33324 25848 33376 25857
rect 33968 25848 34020 25900
rect 34152 25848 34204 25900
rect 34520 25891 34572 25900
rect 34520 25857 34529 25891
rect 34529 25857 34563 25891
rect 34563 25857 34572 25891
rect 34520 25848 34572 25857
rect 35348 25891 35400 25900
rect 35348 25857 35357 25891
rect 35357 25857 35391 25891
rect 35391 25857 35400 25891
rect 35348 25848 35400 25857
rect 35716 25848 35768 25900
rect 37372 25848 37424 25900
rect 38936 25848 38988 25900
rect 41696 25848 41748 25900
rect 37188 25780 37240 25832
rect 32036 25712 32088 25764
rect 29000 25644 29052 25696
rect 30840 25644 30892 25696
rect 31392 25644 31444 25696
rect 44180 25644 44232 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 3976 25440 4028 25492
rect 16764 25440 16816 25492
rect 17960 25483 18012 25492
rect 17960 25449 17969 25483
rect 17969 25449 18003 25483
rect 18003 25449 18012 25483
rect 17960 25440 18012 25449
rect 18144 25440 18196 25492
rect 21272 25483 21324 25492
rect 21272 25449 21281 25483
rect 21281 25449 21315 25483
rect 21315 25449 21324 25483
rect 21272 25440 21324 25449
rect 22100 25483 22152 25492
rect 22100 25449 22109 25483
rect 22109 25449 22143 25483
rect 22143 25449 22152 25483
rect 22100 25440 22152 25449
rect 24492 25440 24544 25492
rect 27620 25483 27672 25492
rect 27620 25449 27629 25483
rect 27629 25449 27663 25483
rect 27663 25449 27672 25483
rect 27620 25440 27672 25449
rect 28632 25440 28684 25492
rect 30380 25440 30432 25492
rect 30472 25440 30524 25492
rect 38936 25483 38988 25492
rect 38936 25449 38945 25483
rect 38945 25449 38979 25483
rect 38979 25449 38988 25483
rect 38936 25440 38988 25449
rect 15568 25347 15620 25356
rect 15568 25313 15577 25347
rect 15577 25313 15611 25347
rect 15611 25313 15620 25347
rect 15568 25304 15620 25313
rect 18052 25304 18104 25356
rect 20444 25304 20496 25356
rect 23020 25372 23072 25424
rect 23572 25347 23624 25356
rect 3976 25279 4028 25288
rect 3976 25245 3985 25279
rect 3985 25245 4019 25279
rect 4019 25245 4028 25279
rect 3976 25236 4028 25245
rect 15844 25279 15896 25288
rect 15844 25245 15878 25279
rect 15878 25245 15896 25279
rect 15844 25236 15896 25245
rect 17868 25279 17920 25288
rect 17868 25245 17877 25279
rect 17877 25245 17911 25279
rect 17911 25245 17920 25279
rect 17868 25236 17920 25245
rect 18604 25236 18656 25288
rect 19064 25236 19116 25288
rect 20812 25236 20864 25288
rect 20996 25279 21048 25288
rect 20996 25245 21005 25279
rect 21005 25245 21039 25279
rect 21039 25245 21048 25279
rect 20996 25236 21048 25245
rect 23572 25313 23581 25347
rect 23581 25313 23615 25347
rect 23615 25313 23624 25347
rect 23572 25304 23624 25313
rect 25412 25304 25464 25356
rect 26516 25347 26568 25356
rect 23388 25236 23440 25288
rect 24952 25279 25004 25288
rect 22376 25168 22428 25220
rect 24952 25245 24961 25279
rect 24961 25245 24995 25279
rect 24995 25245 25004 25279
rect 24952 25236 25004 25245
rect 26148 25236 26200 25288
rect 26516 25313 26525 25347
rect 26525 25313 26559 25347
rect 26559 25313 26568 25347
rect 26516 25304 26568 25313
rect 27896 25304 27948 25356
rect 28908 25304 28960 25356
rect 27436 25279 27488 25288
rect 25136 25168 25188 25220
rect 20352 25143 20404 25152
rect 20352 25109 20361 25143
rect 20361 25109 20395 25143
rect 20395 25109 20404 25143
rect 20352 25100 20404 25109
rect 23112 25100 23164 25152
rect 27436 25245 27445 25279
rect 27445 25245 27479 25279
rect 27479 25245 27488 25279
rect 27436 25236 27488 25245
rect 27528 25236 27580 25288
rect 28632 25279 28684 25288
rect 28632 25245 28641 25279
rect 28641 25245 28675 25279
rect 28675 25245 28684 25279
rect 28632 25236 28684 25245
rect 29000 25279 29052 25288
rect 29000 25245 29009 25279
rect 29009 25245 29043 25279
rect 29043 25245 29052 25279
rect 32128 25304 32180 25356
rect 41420 25304 41472 25356
rect 43904 25304 43956 25356
rect 44088 25347 44140 25356
rect 44088 25313 44097 25347
rect 44097 25313 44131 25347
rect 44131 25313 44140 25347
rect 44088 25304 44140 25313
rect 29000 25236 29052 25245
rect 31024 25236 31076 25288
rect 31484 25279 31536 25288
rect 31484 25245 31493 25279
rect 31493 25245 31527 25279
rect 31527 25245 31536 25279
rect 31484 25236 31536 25245
rect 30748 25168 30800 25220
rect 31208 25168 31260 25220
rect 33876 25279 33928 25288
rect 33876 25245 33894 25279
rect 33894 25245 33928 25279
rect 33876 25236 33928 25245
rect 34060 25236 34112 25288
rect 39304 25279 39356 25288
rect 39304 25245 39313 25279
rect 39313 25245 39347 25279
rect 39347 25245 39356 25279
rect 39304 25236 39356 25245
rect 42340 25279 42392 25288
rect 42340 25245 42349 25279
rect 42349 25245 42383 25279
rect 42383 25245 42392 25279
rect 42340 25236 42392 25245
rect 40868 25168 40920 25220
rect 42524 25211 42576 25220
rect 30196 25100 30248 25152
rect 30564 25143 30616 25152
rect 30564 25109 30589 25143
rect 30589 25109 30616 25143
rect 30564 25100 30616 25109
rect 31760 25143 31812 25152
rect 31760 25109 31769 25143
rect 31769 25109 31803 25143
rect 31803 25109 31812 25143
rect 42524 25177 42533 25211
rect 42533 25177 42567 25211
rect 42567 25177 42576 25211
rect 42524 25168 42576 25177
rect 31760 25100 31812 25109
rect 43996 25100 44048 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 19984 24896 20036 24948
rect 30380 24896 30432 24948
rect 28632 24828 28684 24880
rect 20352 24803 20404 24812
rect 20352 24769 20361 24803
rect 20361 24769 20395 24803
rect 20395 24769 20404 24803
rect 20352 24760 20404 24769
rect 22376 24760 22428 24812
rect 23296 24803 23348 24812
rect 23296 24769 23305 24803
rect 23305 24769 23339 24803
rect 23339 24769 23348 24803
rect 23296 24760 23348 24769
rect 24952 24760 25004 24812
rect 22284 24692 22336 24744
rect 24032 24692 24084 24744
rect 24492 24624 24544 24676
rect 23204 24556 23256 24608
rect 25596 24803 25648 24812
rect 25596 24769 25605 24803
rect 25605 24769 25639 24803
rect 25639 24769 25648 24803
rect 25596 24760 25648 24769
rect 26148 24760 26200 24812
rect 29092 24803 29144 24812
rect 29092 24769 29101 24803
rect 29101 24769 29135 24803
rect 29135 24769 29144 24803
rect 29092 24760 29144 24769
rect 29552 24803 29604 24812
rect 29552 24769 29561 24803
rect 29561 24769 29595 24803
rect 29595 24769 29604 24803
rect 29552 24760 29604 24769
rect 31024 24803 31076 24812
rect 31024 24769 31033 24803
rect 31033 24769 31067 24803
rect 31067 24769 31076 24803
rect 31024 24760 31076 24769
rect 31760 24828 31812 24880
rect 31300 24760 31352 24812
rect 32312 24803 32364 24812
rect 32312 24769 32321 24803
rect 32321 24769 32355 24803
rect 32355 24769 32364 24803
rect 32312 24760 32364 24769
rect 39304 24896 39356 24948
rect 37188 24828 37240 24880
rect 38568 24803 38620 24812
rect 38568 24769 38602 24803
rect 38602 24769 38620 24803
rect 25412 24735 25464 24744
rect 25412 24701 25421 24735
rect 25421 24701 25455 24735
rect 25455 24701 25464 24735
rect 25412 24692 25464 24701
rect 29000 24692 29052 24744
rect 31116 24735 31168 24744
rect 25872 24667 25924 24676
rect 25872 24633 25881 24667
rect 25881 24633 25915 24667
rect 25915 24633 25924 24667
rect 25872 24624 25924 24633
rect 27620 24624 27672 24676
rect 29460 24624 29512 24676
rect 31116 24701 31125 24735
rect 31125 24701 31159 24735
rect 31159 24701 31168 24735
rect 31116 24692 31168 24701
rect 38568 24760 38620 24769
rect 40040 24760 40092 24812
rect 42432 24803 42484 24812
rect 42432 24769 42441 24803
rect 42441 24769 42475 24803
rect 42475 24769 42484 24803
rect 42432 24760 42484 24769
rect 43260 24803 43312 24812
rect 43260 24769 43269 24803
rect 43269 24769 43303 24803
rect 43303 24769 43312 24803
rect 43260 24760 43312 24769
rect 43720 24760 43772 24812
rect 43996 24803 44048 24812
rect 43996 24769 44005 24803
rect 44005 24769 44039 24803
rect 44039 24769 44048 24803
rect 43996 24760 44048 24769
rect 30564 24624 30616 24676
rect 39948 24692 40000 24744
rect 41788 24692 41840 24744
rect 30288 24556 30340 24608
rect 32404 24624 32456 24676
rect 32036 24556 32088 24608
rect 32312 24556 32364 24608
rect 32956 24599 33008 24608
rect 32956 24565 32965 24599
rect 32965 24565 32999 24599
rect 32999 24565 33008 24599
rect 32956 24556 33008 24565
rect 41512 24599 41564 24608
rect 41512 24565 41521 24599
rect 41521 24565 41555 24599
rect 41555 24565 41564 24599
rect 41512 24556 41564 24565
rect 43352 24599 43404 24608
rect 43352 24565 43361 24599
rect 43361 24565 43395 24599
rect 43395 24565 43404 24599
rect 43352 24556 43404 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 26148 24395 26200 24404
rect 26148 24361 26157 24395
rect 26157 24361 26191 24395
rect 26191 24361 26200 24395
rect 26148 24352 26200 24361
rect 27436 24352 27488 24404
rect 27896 24395 27948 24404
rect 27896 24361 27905 24395
rect 27905 24361 27939 24395
rect 27939 24361 27948 24395
rect 27896 24352 27948 24361
rect 29552 24352 29604 24404
rect 30564 24352 30616 24404
rect 31392 24352 31444 24404
rect 31760 24352 31812 24404
rect 15568 24259 15620 24268
rect 15568 24225 15577 24259
rect 15577 24225 15611 24259
rect 15611 24225 15620 24259
rect 15568 24216 15620 24225
rect 18144 24216 18196 24268
rect 20168 24259 20220 24268
rect 16396 24148 16448 24200
rect 20168 24225 20177 24259
rect 20177 24225 20211 24259
rect 20211 24225 20220 24259
rect 20168 24216 20220 24225
rect 20444 24259 20496 24268
rect 20444 24225 20453 24259
rect 20453 24225 20487 24259
rect 20487 24225 20496 24259
rect 20444 24216 20496 24225
rect 25596 24216 25648 24268
rect 18604 24148 18656 24200
rect 22376 24148 22428 24200
rect 23756 24191 23808 24200
rect 23756 24157 23765 24191
rect 23765 24157 23799 24191
rect 23799 24157 23808 24191
rect 23756 24148 23808 24157
rect 17960 24080 18012 24132
rect 23480 24123 23532 24132
rect 23480 24089 23489 24123
rect 23489 24089 23523 24123
rect 23523 24089 23532 24123
rect 23480 24080 23532 24089
rect 24032 24080 24084 24132
rect 25412 24148 25464 24200
rect 26240 24191 26292 24200
rect 26240 24157 26249 24191
rect 26249 24157 26283 24191
rect 26283 24157 26292 24191
rect 26240 24148 26292 24157
rect 28724 24284 28776 24336
rect 30380 24284 30432 24336
rect 27068 24148 27120 24200
rect 27528 24191 27580 24200
rect 27528 24157 27537 24191
rect 27537 24157 27571 24191
rect 27571 24157 27580 24191
rect 27528 24148 27580 24157
rect 27712 24191 27764 24200
rect 27712 24157 27721 24191
rect 27721 24157 27755 24191
rect 27755 24157 27764 24191
rect 27712 24148 27764 24157
rect 28724 24148 28776 24200
rect 30196 24216 30248 24268
rect 32036 24259 32088 24268
rect 30656 24148 30708 24200
rect 32036 24225 32045 24259
rect 32045 24225 32079 24259
rect 32079 24225 32088 24259
rect 32036 24216 32088 24225
rect 32956 24352 33008 24404
rect 41696 24352 41748 24404
rect 42524 24352 42576 24404
rect 41512 24216 41564 24268
rect 42708 24259 42760 24268
rect 42708 24225 42717 24259
rect 42717 24225 42751 24259
rect 42751 24225 42760 24259
rect 42708 24216 42760 24225
rect 43352 24216 43404 24268
rect 44180 24259 44232 24268
rect 44180 24225 44189 24259
rect 44189 24225 44223 24259
rect 44223 24225 44232 24259
rect 44180 24216 44232 24225
rect 27344 24080 27396 24132
rect 16948 24055 17000 24064
rect 16948 24021 16957 24055
rect 16957 24021 16991 24055
rect 16991 24021 17000 24055
rect 16948 24012 17000 24021
rect 23572 24055 23624 24064
rect 23572 24021 23587 24055
rect 23587 24021 23621 24055
rect 23621 24021 23624 24055
rect 23572 24012 23624 24021
rect 30748 24080 30800 24132
rect 32220 24191 32272 24200
rect 32220 24157 32229 24191
rect 32229 24157 32263 24191
rect 32263 24157 32272 24191
rect 32220 24148 32272 24157
rect 37188 24148 37240 24200
rect 37832 24191 37884 24200
rect 37832 24157 37841 24191
rect 37841 24157 37875 24191
rect 37875 24157 37884 24191
rect 37832 24148 37884 24157
rect 38016 24191 38068 24200
rect 38016 24157 38025 24191
rect 38025 24157 38059 24191
rect 38059 24157 38068 24191
rect 38016 24148 38068 24157
rect 40868 24191 40920 24200
rect 40868 24157 40877 24191
rect 40877 24157 40911 24191
rect 40911 24157 40920 24191
rect 40868 24148 40920 24157
rect 41604 24148 41656 24200
rect 41696 24191 41748 24200
rect 41696 24157 41705 24191
rect 41705 24157 41739 24191
rect 41739 24157 41748 24191
rect 41696 24148 41748 24157
rect 42432 24148 42484 24200
rect 30564 24012 30616 24064
rect 31300 24012 31352 24064
rect 31576 24080 31628 24132
rect 38752 24080 38804 24132
rect 31668 24012 31720 24064
rect 35900 24012 35952 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 17960 23851 18012 23860
rect 17960 23817 17969 23851
rect 17969 23817 18003 23851
rect 18003 23817 18012 23851
rect 17960 23808 18012 23817
rect 19432 23808 19484 23860
rect 23572 23808 23624 23860
rect 25596 23808 25648 23860
rect 26240 23808 26292 23860
rect 27528 23808 27580 23860
rect 19708 23740 19760 23792
rect 2136 23715 2188 23724
rect 2136 23681 2145 23715
rect 2145 23681 2179 23715
rect 2179 23681 2188 23715
rect 2136 23672 2188 23681
rect 10968 23672 11020 23724
rect 15752 23672 15804 23724
rect 16028 23672 16080 23724
rect 17224 23715 17276 23724
rect 17224 23681 17233 23715
rect 17233 23681 17267 23715
rect 17267 23681 17276 23715
rect 17224 23672 17276 23681
rect 18144 23715 18196 23724
rect 18144 23681 18153 23715
rect 18153 23681 18187 23715
rect 18187 23681 18196 23715
rect 18144 23672 18196 23681
rect 18236 23715 18288 23724
rect 18236 23681 18245 23715
rect 18245 23681 18279 23715
rect 18279 23681 18288 23715
rect 18236 23672 18288 23681
rect 16396 23604 16448 23656
rect 19156 23715 19208 23724
rect 19156 23681 19165 23715
rect 19165 23681 19199 23715
rect 19199 23681 19208 23715
rect 19156 23672 19208 23681
rect 20076 23672 20128 23724
rect 20444 23740 20496 23792
rect 22376 23783 22428 23792
rect 22376 23749 22385 23783
rect 22385 23749 22419 23783
rect 22419 23749 22428 23783
rect 22376 23740 22428 23749
rect 27712 23740 27764 23792
rect 28724 23740 28776 23792
rect 23664 23715 23716 23724
rect 23664 23681 23673 23715
rect 23673 23681 23707 23715
rect 23707 23681 23716 23715
rect 23664 23672 23716 23681
rect 27804 23715 27856 23724
rect 27804 23681 27813 23715
rect 27813 23681 27847 23715
rect 27847 23681 27856 23715
rect 27804 23672 27856 23681
rect 27988 23715 28040 23724
rect 27988 23681 27997 23715
rect 27997 23681 28031 23715
rect 28031 23681 28040 23715
rect 27988 23672 28040 23681
rect 18604 23647 18656 23656
rect 3056 23536 3108 23588
rect 18604 23613 18613 23647
rect 18613 23613 18647 23647
rect 18647 23613 18656 23647
rect 18604 23604 18656 23613
rect 30472 23808 30524 23860
rect 30932 23808 30984 23860
rect 31576 23851 31628 23860
rect 30380 23715 30432 23724
rect 30380 23681 30389 23715
rect 30389 23681 30423 23715
rect 30423 23681 30432 23715
rect 30380 23672 30432 23681
rect 30564 23715 30616 23724
rect 30564 23681 30573 23715
rect 30573 23681 30607 23715
rect 30607 23681 30616 23715
rect 30564 23672 30616 23681
rect 31116 23715 31168 23724
rect 31116 23681 31125 23715
rect 31125 23681 31159 23715
rect 31159 23681 31168 23715
rect 31116 23672 31168 23681
rect 31576 23817 31585 23851
rect 31585 23817 31619 23851
rect 31619 23817 31628 23851
rect 31576 23808 31628 23817
rect 37832 23808 37884 23860
rect 38568 23808 38620 23860
rect 42340 23808 42392 23860
rect 42800 23808 42852 23860
rect 43352 23808 43404 23860
rect 31668 23740 31720 23792
rect 31944 23672 31996 23724
rect 22100 23536 22152 23588
rect 28540 23536 28592 23588
rect 31392 23536 31444 23588
rect 31576 23604 31628 23656
rect 32404 23672 32456 23724
rect 34060 23715 34112 23724
rect 33324 23647 33376 23656
rect 33324 23613 33333 23647
rect 33333 23613 33367 23647
rect 33367 23613 33376 23647
rect 33324 23604 33376 23613
rect 34060 23681 34069 23715
rect 34069 23681 34103 23715
rect 34103 23681 34112 23715
rect 34060 23672 34112 23681
rect 34152 23672 34204 23724
rect 33968 23604 34020 23656
rect 33876 23536 33928 23588
rect 36360 23672 36412 23724
rect 37372 23672 37424 23724
rect 39028 23672 39080 23724
rect 41604 23672 41656 23724
rect 41788 23715 41840 23724
rect 41788 23681 41797 23715
rect 41797 23681 41831 23715
rect 41831 23681 41840 23715
rect 41788 23672 41840 23681
rect 42800 23672 42852 23724
rect 43260 23715 43312 23724
rect 43260 23681 43269 23715
rect 43269 23681 43303 23715
rect 43303 23681 43312 23715
rect 43260 23672 43312 23681
rect 35532 23604 35584 23656
rect 38752 23647 38804 23656
rect 38752 23613 38761 23647
rect 38761 23613 38795 23647
rect 38795 23613 38804 23647
rect 38752 23604 38804 23613
rect 38844 23647 38896 23656
rect 38844 23613 38853 23647
rect 38853 23613 38887 23647
rect 38887 23613 38896 23647
rect 38844 23604 38896 23613
rect 2780 23511 2832 23520
rect 2780 23477 2789 23511
rect 2789 23477 2823 23511
rect 2823 23477 2832 23511
rect 2780 23468 2832 23477
rect 15936 23468 15988 23520
rect 19984 23468 20036 23520
rect 21272 23468 21324 23520
rect 27436 23468 27488 23520
rect 29276 23468 29328 23520
rect 30748 23468 30800 23520
rect 31576 23468 31628 23520
rect 33416 23511 33468 23520
rect 33416 23477 33425 23511
rect 33425 23477 33459 23511
rect 33459 23477 33468 23511
rect 33416 23468 33468 23477
rect 42340 23468 42392 23520
rect 42524 23468 42576 23520
rect 44180 23468 44232 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 17224 23264 17276 23316
rect 23480 23264 23532 23316
rect 23756 23264 23808 23316
rect 25044 23264 25096 23316
rect 26700 23264 26752 23316
rect 27804 23264 27856 23316
rect 34152 23264 34204 23316
rect 38016 23264 38068 23316
rect 41788 23264 41840 23316
rect 19432 23196 19484 23248
rect 30656 23196 30708 23248
rect 35900 23196 35952 23248
rect 1400 23171 1452 23180
rect 1400 23137 1409 23171
rect 1409 23137 1443 23171
rect 1443 23137 1452 23171
rect 1400 23128 1452 23137
rect 2780 23128 2832 23180
rect 16948 23128 17000 23180
rect 18052 23128 18104 23180
rect 18604 23128 18656 23180
rect 15476 23060 15528 23112
rect 19340 23060 19392 23112
rect 20444 23128 20496 23180
rect 23848 23128 23900 23180
rect 24584 23128 24636 23180
rect 26424 23128 26476 23180
rect 19708 23103 19760 23112
rect 19708 23069 19743 23103
rect 19743 23069 19760 23103
rect 19708 23060 19760 23069
rect 20076 23060 20128 23112
rect 21272 23103 21324 23112
rect 21272 23069 21306 23103
rect 21306 23069 21324 23103
rect 3056 23035 3108 23044
rect 3056 23001 3065 23035
rect 3065 23001 3099 23035
rect 3099 23001 3108 23035
rect 3056 22992 3108 23001
rect 15660 23035 15712 23044
rect 15660 23001 15694 23035
rect 15694 23001 15712 23035
rect 15660 22992 15712 23001
rect 18236 22992 18288 23044
rect 20352 22992 20404 23044
rect 19248 22967 19300 22976
rect 19248 22933 19257 22967
rect 19257 22933 19291 22967
rect 19291 22933 19300 22967
rect 19248 22924 19300 22933
rect 21272 23060 21324 23069
rect 24032 23060 24084 23112
rect 24400 23103 24452 23112
rect 24400 23069 24409 23103
rect 24409 23069 24443 23103
rect 24443 23069 24452 23103
rect 24400 23060 24452 23069
rect 24860 23060 24912 23112
rect 27344 23128 27396 23180
rect 28080 23103 28132 23112
rect 21456 22924 21508 22976
rect 23572 22992 23624 23044
rect 26240 22992 26292 23044
rect 28080 23069 28089 23103
rect 28089 23069 28123 23103
rect 28123 23069 28132 23103
rect 28080 23060 28132 23069
rect 30380 23128 30432 23180
rect 30932 23128 30984 23180
rect 37832 23128 37884 23180
rect 39948 23171 40000 23180
rect 39948 23137 39957 23171
rect 39957 23137 39991 23171
rect 39991 23137 40000 23171
rect 39948 23128 40000 23137
rect 42708 23171 42760 23180
rect 42708 23137 42717 23171
rect 42717 23137 42751 23171
rect 42751 23137 42760 23171
rect 42708 23128 42760 23137
rect 44180 23171 44232 23180
rect 44180 23137 44189 23171
rect 44189 23137 44223 23171
rect 44223 23137 44232 23171
rect 44180 23128 44232 23137
rect 30012 23035 30064 23044
rect 30012 23001 30021 23035
rect 30021 23001 30055 23035
rect 30055 23001 30064 23035
rect 31024 23103 31076 23112
rect 31024 23069 31033 23103
rect 31033 23069 31067 23103
rect 31067 23069 31076 23103
rect 31024 23060 31076 23069
rect 33416 23060 33468 23112
rect 33876 23103 33928 23112
rect 33876 23069 33885 23103
rect 33885 23069 33919 23103
rect 33919 23069 33928 23103
rect 33876 23060 33928 23069
rect 34428 23060 34480 23112
rect 36360 23103 36412 23112
rect 36360 23069 36369 23103
rect 36369 23069 36403 23103
rect 36403 23069 36412 23103
rect 36360 23060 36412 23069
rect 30012 22992 30064 23001
rect 23296 22924 23348 22976
rect 24584 22967 24636 22976
rect 24584 22933 24593 22967
rect 24593 22933 24627 22967
rect 24627 22933 24636 22967
rect 24584 22924 24636 22933
rect 30196 22924 30248 22976
rect 31392 22992 31444 23044
rect 37648 23060 37700 23112
rect 38752 23060 38804 23112
rect 38844 23103 38896 23112
rect 38844 23069 38853 23103
rect 38853 23069 38887 23103
rect 38887 23069 38896 23103
rect 38844 23060 38896 23069
rect 39028 23060 39080 23112
rect 37372 22992 37424 23044
rect 43444 22992 43496 23044
rect 33968 22924 34020 22976
rect 38200 22924 38252 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 15476 22720 15528 22772
rect 6368 22627 6420 22636
rect 6368 22593 6377 22627
rect 6377 22593 6411 22627
rect 6411 22593 6420 22627
rect 6368 22584 6420 22593
rect 15752 22627 15804 22636
rect 15752 22593 15761 22627
rect 15761 22593 15795 22627
rect 15795 22593 15804 22627
rect 15752 22584 15804 22593
rect 1952 22559 2004 22568
rect 1952 22525 1961 22559
rect 1961 22525 1995 22559
rect 1995 22525 2004 22559
rect 1952 22516 2004 22525
rect 2872 22516 2924 22568
rect 2964 22559 3016 22568
rect 2964 22525 2973 22559
rect 2973 22525 3007 22559
rect 3007 22525 3016 22559
rect 2964 22516 3016 22525
rect 6184 22516 6236 22568
rect 15660 22516 15712 22568
rect 15936 22627 15988 22636
rect 15936 22593 15945 22627
rect 15945 22593 15979 22627
rect 15979 22593 15988 22627
rect 15936 22584 15988 22593
rect 16120 22627 16172 22636
rect 16120 22593 16129 22627
rect 16129 22593 16163 22627
rect 16163 22593 16172 22627
rect 19156 22720 19208 22772
rect 16120 22584 16172 22593
rect 17224 22584 17276 22636
rect 17776 22627 17828 22636
rect 17776 22593 17785 22627
rect 17785 22593 17819 22627
rect 17819 22593 17828 22627
rect 17776 22584 17828 22593
rect 16304 22516 16356 22568
rect 16672 22380 16724 22432
rect 16948 22423 17000 22432
rect 16948 22389 16957 22423
rect 16957 22389 16991 22423
rect 16991 22389 17000 22423
rect 16948 22380 17000 22389
rect 18052 22448 18104 22500
rect 19432 22652 19484 22704
rect 19248 22584 19300 22636
rect 24584 22720 24636 22772
rect 33324 22720 33376 22772
rect 23572 22652 23624 22704
rect 25228 22652 25280 22704
rect 20812 22584 20864 22636
rect 22468 22627 22520 22636
rect 22468 22593 22477 22627
rect 22477 22593 22511 22627
rect 22511 22593 22520 22627
rect 22468 22584 22520 22593
rect 24400 22584 24452 22636
rect 26700 22652 26752 22704
rect 27068 22652 27120 22704
rect 27528 22652 27580 22704
rect 26424 22584 26476 22636
rect 27252 22584 27304 22636
rect 27988 22584 28040 22636
rect 28632 22584 28684 22636
rect 31392 22652 31444 22704
rect 29828 22627 29880 22636
rect 29828 22593 29837 22627
rect 29837 22593 29871 22627
rect 29871 22593 29880 22627
rect 29828 22584 29880 22593
rect 23572 22516 23624 22568
rect 26240 22516 26292 22568
rect 27528 22559 27580 22568
rect 27528 22525 27537 22559
rect 27537 22525 27571 22559
rect 27571 22525 27580 22559
rect 27528 22516 27580 22525
rect 30012 22516 30064 22568
rect 30748 22584 30800 22636
rect 30932 22584 30984 22636
rect 18604 22380 18656 22432
rect 20444 22448 20496 22500
rect 31944 22584 31996 22636
rect 34336 22627 34388 22636
rect 34336 22593 34345 22627
rect 34345 22593 34379 22627
rect 34379 22593 34388 22627
rect 34336 22584 34388 22593
rect 33140 22491 33192 22500
rect 33140 22457 33149 22491
rect 33149 22457 33183 22491
rect 33183 22457 33192 22491
rect 33140 22448 33192 22457
rect 33784 22448 33836 22500
rect 33968 22516 34020 22568
rect 34612 22627 34664 22636
rect 34612 22593 34621 22627
rect 34621 22593 34655 22627
rect 34655 22593 34664 22627
rect 35900 22652 35952 22704
rect 34612 22584 34664 22593
rect 40040 22720 40092 22772
rect 42800 22763 42852 22772
rect 42800 22729 42809 22763
rect 42809 22729 42843 22763
rect 42843 22729 42852 22763
rect 42800 22720 42852 22729
rect 43444 22763 43496 22772
rect 43444 22729 43453 22763
rect 43453 22729 43487 22763
rect 43487 22729 43496 22763
rect 43444 22720 43496 22729
rect 38844 22652 38896 22704
rect 39028 22695 39080 22704
rect 39028 22661 39037 22695
rect 39037 22661 39071 22695
rect 39071 22661 39080 22695
rect 39028 22652 39080 22661
rect 35532 22516 35584 22568
rect 35900 22516 35952 22568
rect 34796 22448 34848 22500
rect 37648 22584 37700 22636
rect 38200 22627 38252 22636
rect 38200 22593 38209 22627
rect 38209 22593 38243 22627
rect 38243 22593 38252 22627
rect 38200 22584 38252 22593
rect 39120 22584 39172 22636
rect 41604 22584 41656 22636
rect 43076 22584 43128 22636
rect 38844 22516 38896 22568
rect 42432 22559 42484 22568
rect 42432 22525 42441 22559
rect 42441 22525 42475 22559
rect 42475 22525 42484 22559
rect 42432 22516 42484 22525
rect 38752 22448 38804 22500
rect 20076 22423 20128 22432
rect 20076 22389 20085 22423
rect 20085 22389 20119 22423
rect 20119 22389 20128 22423
rect 20076 22380 20128 22389
rect 20628 22380 20680 22432
rect 20904 22380 20956 22432
rect 30472 22380 30524 22432
rect 32772 22380 32824 22432
rect 33508 22423 33560 22432
rect 33508 22389 33517 22423
rect 33517 22389 33551 22423
rect 33551 22389 33560 22423
rect 33508 22380 33560 22389
rect 34704 22380 34756 22432
rect 38108 22380 38160 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 1952 22176 2004 22228
rect 6184 22176 6236 22228
rect 25872 22151 25924 22160
rect 25872 22117 25881 22151
rect 25881 22117 25915 22151
rect 25915 22117 25924 22151
rect 25872 22108 25924 22117
rect 28080 22108 28132 22160
rect 2872 22083 2924 22092
rect 2872 22049 2881 22083
rect 2881 22049 2915 22083
rect 2915 22049 2924 22083
rect 2872 22040 2924 22049
rect 3148 22040 3200 22092
rect 6092 22040 6144 22092
rect 16304 22040 16356 22092
rect 18144 22040 18196 22092
rect 19340 22083 19392 22092
rect 19340 22049 19349 22083
rect 19349 22049 19383 22083
rect 19383 22049 19392 22083
rect 19340 22040 19392 22049
rect 25964 22083 26016 22092
rect 25964 22049 25973 22083
rect 25973 22049 26007 22083
rect 26007 22049 26016 22083
rect 25964 22040 26016 22049
rect 27436 22040 27488 22092
rect 30196 22040 30248 22092
rect 3976 21972 4028 22024
rect 6184 21972 6236 22024
rect 6368 21972 6420 22024
rect 15292 21972 15344 22024
rect 15752 21947 15804 21956
rect 15752 21913 15761 21947
rect 15761 21913 15795 21947
rect 15795 21913 15804 21947
rect 15752 21904 15804 21913
rect 16672 21972 16724 22024
rect 18328 21904 18380 21956
rect 18972 21904 19024 21956
rect 19984 21972 20036 22024
rect 20260 22015 20312 22024
rect 19340 21904 19392 21956
rect 20260 21981 20269 22015
rect 20269 21981 20303 22015
rect 20303 21981 20312 22015
rect 20260 21972 20312 21981
rect 20904 22015 20956 22024
rect 20904 21981 20913 22015
rect 20913 21981 20947 22015
rect 20947 21981 20956 22015
rect 20904 21972 20956 21981
rect 21456 21972 21508 22024
rect 26332 21972 26384 22024
rect 26976 22015 27028 22024
rect 14740 21836 14792 21888
rect 16396 21836 16448 21888
rect 19248 21836 19300 21888
rect 26424 21904 26476 21956
rect 26976 21981 26985 22015
rect 26985 21981 27019 22015
rect 27019 21981 27028 22015
rect 26976 21972 27028 21981
rect 27344 21972 27396 22024
rect 27528 21904 27580 21956
rect 30380 22108 30432 22160
rect 31024 22108 31076 22160
rect 33784 22151 33836 22160
rect 33784 22117 33793 22151
rect 33793 22117 33827 22151
rect 33827 22117 33836 22151
rect 33784 22108 33836 22117
rect 33968 22219 34020 22228
rect 33968 22185 33977 22219
rect 33977 22185 34011 22219
rect 34011 22185 34020 22219
rect 33968 22176 34020 22185
rect 41696 22176 41748 22228
rect 42432 22176 42484 22228
rect 38752 22108 38804 22160
rect 31944 22083 31996 22092
rect 31944 22049 31953 22083
rect 31953 22049 31987 22083
rect 31987 22049 31996 22083
rect 31944 22040 31996 22049
rect 42340 22083 42392 22092
rect 22928 21879 22980 21888
rect 22928 21845 22937 21879
rect 22937 21845 22971 21879
rect 22971 21845 22980 21879
rect 22928 21836 22980 21845
rect 26056 21879 26108 21888
rect 26056 21845 26065 21879
rect 26065 21845 26099 21879
rect 26099 21845 26108 21879
rect 26056 21836 26108 21845
rect 27160 21879 27212 21888
rect 27160 21845 27169 21879
rect 27169 21845 27203 21879
rect 27203 21845 27212 21879
rect 27160 21836 27212 21845
rect 27344 21836 27396 21888
rect 29092 21836 29144 21888
rect 32496 22015 32548 22024
rect 32496 21981 32505 22015
rect 32505 21981 32539 22015
rect 32539 21981 32548 22015
rect 32772 22015 32824 22024
rect 32496 21972 32548 21981
rect 32772 21981 32781 22015
rect 32781 21981 32815 22015
rect 32815 21981 32824 22015
rect 32772 21972 32824 21981
rect 34704 22015 34756 22024
rect 34704 21981 34713 22015
rect 34713 21981 34747 22015
rect 34747 21981 34756 22015
rect 34704 21972 34756 21981
rect 35532 21972 35584 22024
rect 35808 22015 35860 22024
rect 35808 21981 35817 22015
rect 35817 21981 35851 22015
rect 35851 21981 35860 22015
rect 35808 21972 35860 21981
rect 35992 22015 36044 22024
rect 35992 21981 36001 22015
rect 36001 21981 36035 22015
rect 36035 21981 36044 22015
rect 35992 21972 36044 21981
rect 37648 22015 37700 22024
rect 37648 21981 37657 22015
rect 37657 21981 37691 22015
rect 37691 21981 37700 22015
rect 37648 21972 37700 21981
rect 38844 22015 38896 22024
rect 38844 21981 38853 22015
rect 38853 21981 38887 22015
rect 38887 21981 38896 22015
rect 38844 21972 38896 21981
rect 39120 22015 39172 22024
rect 39120 21981 39129 22015
rect 39129 21981 39163 22015
rect 39163 21981 39172 22015
rect 39120 21972 39172 21981
rect 40408 22015 40460 22024
rect 40408 21981 40417 22015
rect 40417 21981 40451 22015
rect 40451 21981 40460 22015
rect 40408 21972 40460 21981
rect 42340 22049 42349 22083
rect 42349 22049 42383 22083
rect 42383 22049 42392 22083
rect 42340 22040 42392 22049
rect 42524 22083 42576 22092
rect 42524 22049 42533 22083
rect 42533 22049 42567 22083
rect 42567 22049 42576 22083
rect 42524 22040 42576 22049
rect 42616 22040 42668 22092
rect 41420 21972 41472 22024
rect 31392 21904 31444 21956
rect 31760 21947 31812 21956
rect 31760 21913 31769 21947
rect 31769 21913 31803 21947
rect 31803 21913 31812 21947
rect 31760 21904 31812 21913
rect 31944 21904 31996 21956
rect 34336 21904 34388 21956
rect 38752 21904 38804 21956
rect 40132 21904 40184 21956
rect 30564 21836 30616 21888
rect 31668 21879 31720 21888
rect 31668 21845 31677 21879
rect 31677 21845 31711 21879
rect 31711 21845 31720 21879
rect 31668 21836 31720 21845
rect 32680 21879 32732 21888
rect 32680 21845 32682 21879
rect 32682 21845 32716 21879
rect 32716 21845 32732 21879
rect 32680 21836 32732 21845
rect 34428 21836 34480 21888
rect 34796 21836 34848 21888
rect 36176 21879 36228 21888
rect 36176 21845 36185 21879
rect 36185 21845 36219 21879
rect 36219 21845 36228 21879
rect 36176 21836 36228 21845
rect 38200 21836 38252 21888
rect 39764 21836 39816 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 7932 21632 7984 21684
rect 8208 21632 8260 21684
rect 17776 21632 17828 21684
rect 5540 21496 5592 21548
rect 6368 21564 6420 21616
rect 18144 21607 18196 21616
rect 18144 21573 18153 21607
rect 18153 21573 18187 21607
rect 18187 21573 18196 21607
rect 18144 21564 18196 21573
rect 18236 21539 18288 21548
rect 5172 21428 5224 21480
rect 6552 21428 6604 21480
rect 18236 21505 18245 21539
rect 18245 21505 18279 21539
rect 18279 21505 18288 21539
rect 18236 21496 18288 21505
rect 19248 21607 19300 21616
rect 19248 21573 19257 21607
rect 19257 21573 19291 21607
rect 19291 21573 19300 21607
rect 19248 21564 19300 21573
rect 18972 21539 19024 21548
rect 18972 21505 18981 21539
rect 18981 21505 19015 21539
rect 19015 21505 19024 21539
rect 18972 21496 19024 21505
rect 19064 21539 19116 21548
rect 19064 21505 19073 21539
rect 19073 21505 19107 21539
rect 19107 21505 19116 21539
rect 19432 21632 19484 21684
rect 26332 21632 26384 21684
rect 26976 21632 27028 21684
rect 27252 21675 27304 21684
rect 27252 21641 27261 21675
rect 27261 21641 27295 21675
rect 27295 21641 27304 21675
rect 27252 21632 27304 21641
rect 22284 21564 22336 21616
rect 22468 21564 22520 21616
rect 19064 21496 19116 21505
rect 20076 21496 20128 21548
rect 20260 21496 20312 21548
rect 20812 21496 20864 21548
rect 19524 21428 19576 21480
rect 20628 21428 20680 21480
rect 20352 21360 20404 21412
rect 22376 21496 22428 21548
rect 24584 21539 24636 21548
rect 24584 21505 24618 21539
rect 24618 21505 24636 21539
rect 28080 21564 28132 21616
rect 30932 21632 30984 21684
rect 24584 21496 24636 21505
rect 21456 21428 21508 21480
rect 23664 21428 23716 21480
rect 24308 21471 24360 21480
rect 24308 21437 24317 21471
rect 24317 21437 24351 21471
rect 24351 21437 24360 21471
rect 24308 21428 24360 21437
rect 25964 21428 26016 21480
rect 27344 21428 27396 21480
rect 22100 21360 22152 21412
rect 15476 21292 15528 21344
rect 17500 21292 17552 21344
rect 18236 21292 18288 21344
rect 20444 21292 20496 21344
rect 21732 21292 21784 21344
rect 25872 21292 25924 21344
rect 27528 21292 27580 21344
rect 28632 21471 28684 21480
rect 28632 21437 28641 21471
rect 28641 21437 28675 21471
rect 28675 21437 28684 21471
rect 29828 21564 29880 21616
rect 29368 21496 29420 21548
rect 30748 21564 30800 21616
rect 30840 21564 30892 21616
rect 32496 21632 32548 21684
rect 34336 21632 34388 21684
rect 31668 21564 31720 21616
rect 36084 21632 36136 21684
rect 39120 21632 39172 21684
rect 40132 21675 40184 21684
rect 40132 21641 40141 21675
rect 40141 21641 40175 21675
rect 40175 21641 40184 21675
rect 40132 21632 40184 21641
rect 34796 21607 34848 21616
rect 34796 21573 34814 21607
rect 34814 21573 34848 21607
rect 34796 21564 34848 21573
rect 30564 21539 30616 21548
rect 30564 21505 30573 21539
rect 30573 21505 30607 21539
rect 30607 21505 30616 21539
rect 30564 21496 30616 21505
rect 31944 21496 31996 21548
rect 36176 21496 36228 21548
rect 38200 21496 38252 21548
rect 28632 21428 28684 21437
rect 30196 21428 30248 21480
rect 32312 21428 32364 21480
rect 35348 21428 35400 21480
rect 35900 21428 35952 21480
rect 31576 21360 31628 21412
rect 33048 21360 33100 21412
rect 38752 21428 38804 21480
rect 41696 21496 41748 21548
rect 27896 21292 27948 21344
rect 29368 21292 29420 21344
rect 30380 21292 30432 21344
rect 30840 21292 30892 21344
rect 30932 21335 30984 21344
rect 30932 21301 30941 21335
rect 30941 21301 30975 21335
rect 30975 21301 30984 21335
rect 30932 21292 30984 21301
rect 35440 21292 35492 21344
rect 42064 21292 42116 21344
rect 42616 21292 42668 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 5540 21131 5592 21140
rect 5540 21097 5549 21131
rect 5549 21097 5583 21131
rect 5583 21097 5592 21131
rect 5540 21088 5592 21097
rect 23296 21131 23348 21140
rect 23296 21097 23305 21131
rect 23305 21097 23339 21131
rect 23339 21097 23348 21131
rect 23296 21088 23348 21097
rect 24584 21131 24636 21140
rect 24584 21097 24593 21131
rect 24593 21097 24627 21131
rect 24627 21097 24636 21131
rect 24584 21088 24636 21097
rect 26240 21131 26292 21140
rect 6828 20995 6880 21004
rect 6828 20961 6837 20995
rect 6837 20961 6871 20995
rect 6871 20961 6880 20995
rect 6828 20952 6880 20961
rect 1676 20884 1728 20936
rect 3884 20884 3936 20936
rect 5540 20884 5592 20936
rect 14556 20927 14608 20936
rect 14556 20893 14565 20927
rect 14565 20893 14599 20927
rect 14599 20893 14608 20927
rect 14556 20884 14608 20893
rect 14740 20927 14792 20936
rect 14740 20893 14749 20927
rect 14749 20893 14783 20927
rect 14783 20893 14792 20927
rect 14740 20884 14792 20893
rect 16304 20952 16356 21004
rect 17500 20995 17552 21004
rect 17500 20961 17509 20995
rect 17509 20961 17543 20995
rect 17543 20961 17552 20995
rect 17500 20952 17552 20961
rect 17776 20995 17828 21004
rect 17776 20961 17785 20995
rect 17785 20961 17819 20995
rect 17819 20961 17828 20995
rect 17776 20952 17828 20961
rect 19432 20952 19484 21004
rect 21456 20995 21508 21004
rect 21456 20961 21465 20995
rect 21465 20961 21499 20995
rect 21499 20961 21508 20995
rect 21456 20952 21508 20961
rect 26240 21097 26249 21131
rect 26249 21097 26283 21131
rect 26283 21097 26292 21131
rect 26240 21088 26292 21097
rect 27896 21131 27948 21140
rect 27896 21097 27905 21131
rect 27905 21097 27939 21131
rect 27939 21097 27948 21131
rect 27896 21088 27948 21097
rect 28632 21131 28684 21140
rect 28632 21097 28641 21131
rect 28641 21097 28675 21131
rect 28675 21097 28684 21131
rect 28632 21088 28684 21097
rect 30196 21131 30248 21140
rect 30196 21097 30205 21131
rect 30205 21097 30239 21131
rect 30239 21097 30248 21131
rect 30196 21088 30248 21097
rect 31944 21131 31996 21140
rect 31944 21097 31953 21131
rect 31953 21097 31987 21131
rect 31987 21097 31996 21131
rect 31944 21088 31996 21097
rect 33140 21088 33192 21140
rect 26148 21020 26200 21072
rect 27068 21020 27120 21072
rect 15936 20884 15988 20936
rect 16672 20927 16724 20936
rect 16672 20893 16681 20927
rect 16681 20893 16715 20927
rect 16715 20893 16724 20927
rect 16672 20884 16724 20893
rect 21732 20927 21784 20936
rect 21732 20893 21766 20927
rect 21766 20893 21784 20927
rect 21732 20884 21784 20893
rect 22928 20884 22980 20936
rect 24400 20927 24452 20936
rect 24400 20893 24409 20927
rect 24409 20893 24443 20927
rect 24443 20893 24452 20927
rect 24400 20884 24452 20893
rect 26792 20952 26844 21004
rect 26976 20952 27028 21004
rect 26056 20884 26108 20936
rect 27160 20927 27212 20936
rect 27160 20893 27169 20927
rect 27169 20893 27203 20927
rect 27203 20893 27212 20927
rect 27160 20884 27212 20893
rect 27436 20952 27488 21004
rect 15568 20859 15620 20868
rect 15568 20825 15577 20859
rect 15577 20825 15611 20859
rect 15611 20825 15620 20859
rect 15568 20816 15620 20825
rect 15660 20859 15712 20868
rect 15660 20825 15695 20859
rect 15695 20825 15712 20859
rect 15660 20816 15712 20825
rect 17408 20816 17460 20868
rect 19984 20816 20036 20868
rect 23296 20859 23348 20868
rect 23296 20825 23305 20859
rect 23305 20825 23339 20859
rect 23339 20825 23348 20859
rect 23296 20816 23348 20825
rect 25964 20816 26016 20868
rect 11520 20791 11572 20800
rect 11520 20757 11529 20791
rect 11529 20757 11563 20791
rect 11563 20757 11572 20791
rect 11520 20748 11572 20757
rect 15200 20791 15252 20800
rect 15200 20757 15209 20791
rect 15209 20757 15243 20791
rect 15243 20757 15252 20791
rect 15200 20748 15252 20757
rect 18144 20748 18196 20800
rect 20444 20748 20496 20800
rect 23388 20748 23440 20800
rect 31392 20995 31444 21004
rect 30380 20884 30432 20936
rect 30932 20927 30984 20936
rect 30932 20893 30941 20927
rect 30941 20893 30975 20927
rect 30975 20893 30984 20927
rect 30932 20884 30984 20893
rect 31392 20961 31401 20995
rect 31401 20961 31435 20995
rect 31435 20961 31444 20995
rect 31392 20952 31444 20961
rect 31300 20927 31352 20936
rect 31300 20893 31309 20927
rect 31309 20893 31343 20927
rect 31343 20893 31352 20927
rect 31300 20884 31352 20893
rect 31668 20884 31720 20936
rect 30564 20816 30616 20868
rect 33416 20816 33468 20868
rect 30748 20791 30800 20800
rect 30748 20757 30757 20791
rect 30757 20757 30791 20791
rect 30791 20757 30800 20791
rect 30748 20748 30800 20757
rect 30840 20748 30892 20800
rect 33048 20748 33100 20800
rect 38844 21088 38896 21140
rect 35900 21063 35952 21072
rect 35900 21029 35909 21063
rect 35909 21029 35943 21063
rect 35943 21029 35952 21063
rect 35900 21020 35952 21029
rect 35440 20995 35492 21004
rect 35440 20961 35449 20995
rect 35449 20961 35483 20995
rect 35483 20961 35492 20995
rect 35440 20952 35492 20961
rect 41052 20952 41104 21004
rect 42616 20952 42668 21004
rect 44088 20995 44140 21004
rect 44088 20961 44097 20995
rect 44097 20961 44131 20995
rect 44131 20961 44140 20995
rect 44088 20952 44140 20961
rect 38752 20927 38804 20936
rect 38752 20893 38761 20927
rect 38761 20893 38795 20927
rect 38795 20893 38804 20927
rect 38752 20884 38804 20893
rect 40132 20816 40184 20868
rect 43076 20816 43128 20868
rect 35256 20748 35308 20800
rect 41328 20748 41380 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 16304 20544 16356 20596
rect 16396 20544 16448 20596
rect 1676 20451 1728 20460
rect 1676 20417 1685 20451
rect 1685 20417 1719 20451
rect 1719 20417 1728 20451
rect 1676 20408 1728 20417
rect 11520 20408 11572 20460
rect 12256 20408 12308 20460
rect 15476 20476 15528 20528
rect 14096 20408 14148 20460
rect 15200 20408 15252 20460
rect 15384 20408 15436 20460
rect 2044 20340 2096 20392
rect 2780 20383 2832 20392
rect 2780 20349 2789 20383
rect 2789 20349 2823 20383
rect 2823 20349 2832 20383
rect 2780 20340 2832 20349
rect 12532 20340 12584 20392
rect 17132 20408 17184 20460
rect 17500 20476 17552 20528
rect 18696 20544 18748 20596
rect 19340 20544 19392 20596
rect 19984 20544 20036 20596
rect 19064 20476 19116 20528
rect 37924 20544 37976 20596
rect 41052 20587 41104 20596
rect 17408 20451 17460 20460
rect 17408 20417 17417 20451
rect 17417 20417 17451 20451
rect 17451 20417 17460 20451
rect 18328 20451 18380 20460
rect 17408 20408 17460 20417
rect 17868 20340 17920 20392
rect 18328 20417 18337 20451
rect 18337 20417 18371 20451
rect 18371 20417 18380 20451
rect 18328 20408 18380 20417
rect 19156 20451 19208 20460
rect 19156 20417 19165 20451
rect 19165 20417 19199 20451
rect 19199 20417 19208 20451
rect 19156 20408 19208 20417
rect 19340 20451 19392 20460
rect 19340 20417 19349 20451
rect 19349 20417 19383 20451
rect 19383 20417 19392 20451
rect 19340 20408 19392 20417
rect 19984 20408 20036 20460
rect 20260 20408 20312 20460
rect 20444 20451 20496 20460
rect 20444 20417 20453 20451
rect 20453 20417 20487 20451
rect 20487 20417 20496 20451
rect 20444 20408 20496 20417
rect 20904 20340 20956 20392
rect 22192 20476 22244 20528
rect 26608 20476 26660 20528
rect 29368 20519 29420 20528
rect 29368 20485 29386 20519
rect 29386 20485 29420 20519
rect 29368 20476 29420 20485
rect 32496 20476 32548 20528
rect 22008 20408 22060 20460
rect 24952 20408 25004 20460
rect 29552 20408 29604 20460
rect 30564 20408 30616 20460
rect 31208 20451 31260 20460
rect 31208 20417 31217 20451
rect 31217 20417 31251 20451
rect 31251 20417 31260 20451
rect 31208 20408 31260 20417
rect 31300 20451 31352 20460
rect 31300 20417 31309 20451
rect 31309 20417 31343 20451
rect 31343 20417 31352 20451
rect 31576 20451 31628 20460
rect 31300 20408 31352 20417
rect 31576 20417 31585 20451
rect 31585 20417 31619 20451
rect 31619 20417 31628 20451
rect 31576 20408 31628 20417
rect 31668 20408 31720 20460
rect 32312 20451 32364 20460
rect 32312 20417 32321 20451
rect 32321 20417 32355 20451
rect 32355 20417 32364 20451
rect 32312 20408 32364 20417
rect 33324 20408 33376 20460
rect 35348 20476 35400 20528
rect 23480 20340 23532 20392
rect 24308 20340 24360 20392
rect 24768 20340 24820 20392
rect 33416 20340 33468 20392
rect 38108 20451 38160 20460
rect 38108 20417 38142 20451
rect 38142 20417 38160 20451
rect 38108 20408 38160 20417
rect 40408 20476 40460 20528
rect 39764 20408 39816 20460
rect 41052 20553 41061 20587
rect 41061 20553 41095 20587
rect 41095 20553 41104 20587
rect 41052 20544 41104 20553
rect 43076 20587 43128 20596
rect 43076 20553 43085 20587
rect 43085 20553 43119 20587
rect 43119 20553 43128 20587
rect 43076 20544 43128 20553
rect 8208 20204 8260 20256
rect 22100 20272 22152 20324
rect 23388 20315 23440 20324
rect 23388 20281 23397 20315
rect 23397 20281 23431 20315
rect 23431 20281 23440 20315
rect 23388 20272 23440 20281
rect 26424 20315 26476 20324
rect 26424 20281 26433 20315
rect 26433 20281 26467 20315
rect 26467 20281 26476 20315
rect 26424 20272 26476 20281
rect 35256 20315 35308 20324
rect 35256 20281 35265 20315
rect 35265 20281 35299 20315
rect 35299 20281 35308 20315
rect 35256 20272 35308 20281
rect 15844 20204 15896 20256
rect 22836 20204 22888 20256
rect 24400 20204 24452 20256
rect 31208 20204 31260 20256
rect 39304 20204 39356 20256
rect 43628 20247 43680 20256
rect 43628 20213 43637 20247
rect 43637 20213 43671 20247
rect 43671 20213 43680 20247
rect 43628 20204 43680 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 2044 20043 2096 20052
rect 2044 20009 2053 20043
rect 2053 20009 2087 20043
rect 2087 20009 2096 20043
rect 2044 20000 2096 20009
rect 14556 20000 14608 20052
rect 16396 20000 16448 20052
rect 17408 20000 17460 20052
rect 17868 20000 17920 20052
rect 19340 20000 19392 20052
rect 20076 20043 20128 20052
rect 20076 20009 20085 20043
rect 20085 20009 20119 20043
rect 20119 20009 20128 20043
rect 20076 20000 20128 20009
rect 15568 19932 15620 19984
rect 21824 20000 21876 20052
rect 22284 20043 22336 20052
rect 22284 20009 22293 20043
rect 22293 20009 22327 20043
rect 22327 20009 22336 20043
rect 22284 20000 22336 20009
rect 22744 20000 22796 20052
rect 27436 20043 27488 20052
rect 21180 19932 21232 19984
rect 27436 20009 27445 20043
rect 27445 20009 27479 20043
rect 27479 20009 27488 20043
rect 27436 20000 27488 20009
rect 31576 20000 31628 20052
rect 41420 20000 41472 20052
rect 8852 19864 8904 19916
rect 15844 19907 15896 19916
rect 2136 19839 2188 19848
rect 2136 19805 2145 19839
rect 2145 19805 2179 19839
rect 2179 19805 2188 19839
rect 2136 19796 2188 19805
rect 3976 19796 4028 19848
rect 12256 19839 12308 19848
rect 12256 19805 12265 19839
rect 12265 19805 12299 19839
rect 12299 19805 12308 19839
rect 12256 19796 12308 19805
rect 15844 19873 15853 19907
rect 15853 19873 15887 19907
rect 15887 19873 15896 19907
rect 15844 19864 15896 19873
rect 17132 19839 17184 19848
rect 12808 19728 12860 19780
rect 15292 19728 15344 19780
rect 15936 19728 15988 19780
rect 17132 19805 17141 19839
rect 17141 19805 17175 19839
rect 17175 19805 17184 19839
rect 17132 19796 17184 19805
rect 24768 19864 24820 19916
rect 32496 19907 32548 19916
rect 32496 19873 32505 19907
rect 32505 19873 32539 19907
rect 32539 19873 32548 19907
rect 32496 19864 32548 19873
rect 32956 19907 33008 19916
rect 32956 19873 32965 19907
rect 32965 19873 32999 19907
rect 32999 19873 33008 19907
rect 32956 19864 33008 19873
rect 35348 19864 35400 19916
rect 39304 19907 39356 19916
rect 39304 19873 39313 19907
rect 39313 19873 39347 19907
rect 39347 19873 39356 19907
rect 39304 19864 39356 19873
rect 18144 19771 18196 19780
rect 18144 19737 18153 19771
rect 18153 19737 18187 19771
rect 18187 19737 18196 19771
rect 18144 19728 18196 19737
rect 18328 19771 18380 19780
rect 18328 19737 18358 19771
rect 18358 19737 18380 19771
rect 20076 19796 20128 19848
rect 20904 19839 20956 19848
rect 20904 19805 20913 19839
rect 20913 19805 20947 19839
rect 20947 19805 20956 19839
rect 20904 19796 20956 19805
rect 18328 19728 18380 19737
rect 17500 19660 17552 19712
rect 17684 19660 17736 19712
rect 19064 19660 19116 19712
rect 20260 19660 20312 19712
rect 20352 19660 20404 19712
rect 21640 19660 21692 19712
rect 22836 19839 22888 19848
rect 22836 19805 22845 19839
rect 22845 19805 22879 19839
rect 22879 19805 22888 19839
rect 22836 19796 22888 19805
rect 30564 19796 30616 19848
rect 32680 19796 32732 19848
rect 41604 19864 41656 19916
rect 42064 19907 42116 19916
rect 42064 19873 42073 19907
rect 42073 19873 42107 19907
rect 42107 19873 42116 19907
rect 42064 19864 42116 19873
rect 43076 19907 43128 19916
rect 43076 19873 43085 19907
rect 43085 19873 43119 19907
rect 43119 19873 43128 19907
rect 43076 19864 43128 19873
rect 40132 19839 40184 19848
rect 40132 19805 40141 19839
rect 40141 19805 40175 19839
rect 40175 19805 40184 19839
rect 40132 19796 40184 19805
rect 41512 19796 41564 19848
rect 25320 19728 25372 19780
rect 26332 19771 26384 19780
rect 26332 19737 26366 19771
rect 26366 19737 26384 19771
rect 26332 19728 26384 19737
rect 30380 19728 30432 19780
rect 23020 19703 23072 19712
rect 23020 19669 23029 19703
rect 23029 19669 23063 19703
rect 23063 19669 23072 19703
rect 23020 19660 23072 19669
rect 36912 19660 36964 19712
rect 38936 19703 38988 19712
rect 38936 19669 38945 19703
rect 38945 19669 38979 19703
rect 38979 19669 38988 19703
rect 38936 19660 38988 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 12716 19431 12768 19440
rect 12716 19397 12725 19431
rect 12725 19397 12759 19431
rect 12759 19397 12768 19431
rect 12716 19388 12768 19397
rect 15292 19431 15344 19440
rect 15292 19397 15302 19431
rect 15302 19397 15336 19431
rect 15336 19397 15344 19431
rect 15292 19388 15344 19397
rect 15660 19388 15712 19440
rect 17224 19388 17276 19440
rect 18328 19388 18380 19440
rect 12256 19320 12308 19372
rect 12624 19320 12676 19372
rect 13544 19363 13596 19372
rect 13544 19329 13553 19363
rect 13553 19329 13587 19363
rect 13587 19329 13596 19363
rect 13544 19320 13596 19329
rect 15108 19320 15160 19372
rect 18696 19363 18748 19372
rect 18696 19329 18705 19363
rect 18705 19329 18739 19363
rect 18739 19329 18748 19363
rect 18696 19320 18748 19329
rect 15568 19252 15620 19304
rect 16120 19252 16172 19304
rect 19432 19320 19484 19372
rect 20904 19456 20956 19508
rect 41512 19499 41564 19508
rect 20076 19320 20128 19372
rect 20352 19363 20404 19372
rect 20352 19329 20361 19363
rect 20361 19329 20395 19363
rect 20395 19329 20404 19363
rect 20352 19320 20404 19329
rect 22192 19431 22244 19440
rect 22192 19397 22201 19431
rect 22201 19397 22235 19431
rect 22235 19397 22244 19431
rect 22192 19388 22244 19397
rect 23020 19388 23072 19440
rect 30932 19388 30984 19440
rect 32956 19388 33008 19440
rect 41512 19465 41521 19499
rect 41521 19465 41555 19499
rect 41555 19465 41564 19499
rect 41512 19456 41564 19465
rect 43720 19388 43772 19440
rect 21548 19320 21600 19372
rect 23480 19363 23532 19372
rect 23480 19329 23489 19363
rect 23489 19329 23523 19363
rect 23523 19329 23532 19363
rect 23480 19320 23532 19329
rect 26700 19320 26752 19372
rect 28356 19320 28408 19372
rect 33324 19363 33376 19372
rect 33324 19329 33333 19363
rect 33333 19329 33367 19363
rect 33367 19329 33376 19363
rect 33324 19320 33376 19329
rect 38936 19363 38988 19372
rect 38936 19329 38945 19363
rect 38945 19329 38979 19363
rect 38979 19329 38988 19363
rect 38936 19320 38988 19329
rect 41328 19363 41380 19372
rect 41328 19329 41337 19363
rect 41337 19329 41371 19363
rect 41371 19329 41380 19363
rect 41328 19320 41380 19329
rect 41420 19320 41472 19372
rect 42984 19363 43036 19372
rect 42984 19329 42993 19363
rect 42993 19329 43027 19363
rect 43027 19329 43036 19363
rect 42984 19320 43036 19329
rect 23112 19252 23164 19304
rect 27068 19252 27120 19304
rect 29552 19252 29604 19304
rect 15292 19184 15344 19236
rect 20260 19184 20312 19236
rect 21088 19184 21140 19236
rect 19340 19159 19392 19168
rect 19340 19125 19349 19159
rect 19349 19125 19383 19159
rect 19383 19125 19392 19159
rect 19340 19116 19392 19125
rect 21180 19116 21232 19168
rect 23020 19116 23072 19168
rect 24860 19159 24912 19168
rect 24860 19125 24869 19159
rect 24869 19125 24903 19159
rect 24903 19125 24912 19159
rect 24860 19116 24912 19125
rect 31576 19159 31628 19168
rect 31576 19125 31585 19159
rect 31585 19125 31619 19159
rect 31619 19125 31628 19159
rect 31576 19116 31628 19125
rect 34704 19159 34756 19168
rect 34704 19125 34713 19159
rect 34713 19125 34747 19159
rect 34747 19125 34756 19159
rect 34704 19116 34756 19125
rect 38752 19159 38804 19168
rect 38752 19125 38761 19159
rect 38761 19125 38795 19159
rect 38795 19125 38804 19159
rect 38752 19116 38804 19125
rect 44180 19116 44232 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 13544 18912 13596 18964
rect 16948 18912 17000 18964
rect 19340 18912 19392 18964
rect 26424 18912 26476 18964
rect 15476 18819 15528 18828
rect 15476 18785 15485 18819
rect 15485 18785 15519 18819
rect 15519 18785 15528 18819
rect 15476 18776 15528 18785
rect 17684 18776 17736 18828
rect 2044 18751 2096 18760
rect 2044 18717 2053 18751
rect 2053 18717 2087 18751
rect 2087 18717 2096 18751
rect 2044 18708 2096 18717
rect 12624 18708 12676 18760
rect 15200 18751 15252 18760
rect 15200 18717 15218 18751
rect 15218 18717 15252 18751
rect 15200 18708 15252 18717
rect 16120 18751 16172 18760
rect 11704 18640 11756 18692
rect 14556 18640 14608 18692
rect 16120 18717 16129 18751
rect 16129 18717 16163 18751
rect 16163 18717 16172 18751
rect 16120 18708 16172 18717
rect 17132 18751 17184 18760
rect 17132 18717 17141 18751
rect 17141 18717 17175 18751
rect 17175 18717 17184 18751
rect 17132 18708 17184 18717
rect 17408 18751 17460 18760
rect 17408 18717 17417 18751
rect 17417 18717 17451 18751
rect 17451 18717 17460 18751
rect 17408 18708 17460 18717
rect 18328 18751 18380 18760
rect 18328 18717 18337 18751
rect 18337 18717 18371 18751
rect 18371 18717 18380 18751
rect 18328 18708 18380 18717
rect 18604 18751 18656 18760
rect 18604 18717 18613 18751
rect 18613 18717 18647 18751
rect 18647 18717 18656 18751
rect 18604 18708 18656 18717
rect 21548 18776 21600 18828
rect 21824 18776 21876 18828
rect 23848 18844 23900 18896
rect 26240 18844 26292 18896
rect 34612 18776 34664 18828
rect 34980 18776 35032 18828
rect 35256 18819 35308 18828
rect 35256 18785 35265 18819
rect 35265 18785 35299 18819
rect 35299 18785 35308 18819
rect 35256 18776 35308 18785
rect 23020 18751 23072 18760
rect 23020 18717 23029 18751
rect 23029 18717 23063 18751
rect 23063 18717 23072 18751
rect 23020 18708 23072 18717
rect 24860 18708 24912 18760
rect 25688 18751 25740 18760
rect 25688 18717 25697 18751
rect 25697 18717 25731 18751
rect 25731 18717 25740 18751
rect 25688 18708 25740 18717
rect 16764 18640 16816 18692
rect 17500 18640 17552 18692
rect 19432 18640 19484 18692
rect 25964 18640 26016 18692
rect 26424 18708 26476 18760
rect 26976 18751 27028 18760
rect 26976 18717 26985 18751
rect 26985 18717 27019 18751
rect 27019 18717 27028 18751
rect 26976 18708 27028 18717
rect 28356 18751 28408 18760
rect 28356 18717 28365 18751
rect 28365 18717 28399 18751
rect 28399 18717 28408 18751
rect 28356 18708 28408 18717
rect 29460 18640 29512 18692
rect 29552 18640 29604 18692
rect 31300 18708 31352 18760
rect 34704 18708 34756 18760
rect 34888 18751 34940 18760
rect 34888 18717 34897 18751
rect 34897 18717 34931 18751
rect 34931 18717 34940 18751
rect 34888 18708 34940 18717
rect 30564 18640 30616 18692
rect 34428 18640 34480 18692
rect 36912 18751 36964 18760
rect 36912 18717 36921 18751
rect 36921 18717 36955 18751
rect 36955 18717 36964 18751
rect 36912 18708 36964 18717
rect 43260 18844 43312 18896
rect 42708 18819 42760 18828
rect 42708 18785 42717 18819
rect 42717 18785 42751 18819
rect 42751 18785 42760 18819
rect 42708 18776 42760 18785
rect 44180 18819 44232 18828
rect 44180 18785 44189 18819
rect 44189 18785 44223 18819
rect 44223 18785 44232 18819
rect 44180 18776 44232 18785
rect 43444 18640 43496 18692
rect 14740 18572 14792 18624
rect 16028 18615 16080 18624
rect 16028 18581 16037 18615
rect 16037 18581 16071 18615
rect 16071 18581 16080 18615
rect 16028 18572 16080 18581
rect 17592 18615 17644 18624
rect 17592 18581 17601 18615
rect 17601 18581 17635 18615
rect 17635 18581 17644 18615
rect 17592 18572 17644 18581
rect 18052 18615 18104 18624
rect 18052 18581 18061 18615
rect 18061 18581 18095 18615
rect 18095 18581 18104 18615
rect 18052 18572 18104 18581
rect 25136 18572 25188 18624
rect 27068 18572 27120 18624
rect 27804 18615 27856 18624
rect 27804 18581 27813 18615
rect 27813 18581 27847 18615
rect 27847 18581 27856 18615
rect 27804 18572 27856 18581
rect 32588 18615 32640 18624
rect 32588 18581 32597 18615
rect 32597 18581 32631 18615
rect 32631 18581 32640 18615
rect 32588 18572 32640 18581
rect 35716 18572 35768 18624
rect 37464 18572 37516 18624
rect 38384 18615 38436 18624
rect 38384 18581 38393 18615
rect 38393 18581 38427 18615
rect 38427 18581 38436 18615
rect 38384 18572 38436 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 6276 18368 6328 18420
rect 6828 18368 6880 18420
rect 43444 18411 43496 18420
rect 2044 18275 2096 18284
rect 2044 18241 2053 18275
rect 2053 18241 2087 18275
rect 2087 18241 2096 18275
rect 2044 18232 2096 18241
rect 16028 18300 16080 18352
rect 16764 18300 16816 18352
rect 17040 18343 17092 18352
rect 17040 18309 17049 18343
rect 17049 18309 17083 18343
rect 17083 18309 17092 18343
rect 17040 18300 17092 18309
rect 17592 18300 17644 18352
rect 19432 18300 19484 18352
rect 14464 18232 14516 18284
rect 14556 18232 14608 18284
rect 14740 18275 14792 18284
rect 14740 18241 14749 18275
rect 14749 18241 14783 18275
rect 14783 18241 14792 18275
rect 14740 18232 14792 18241
rect 16948 18232 17000 18284
rect 17684 18232 17736 18284
rect 18144 18232 18196 18284
rect 18696 18275 18748 18284
rect 18696 18241 18705 18275
rect 18705 18241 18739 18275
rect 18739 18241 18748 18275
rect 18696 18232 18748 18241
rect 2872 18164 2924 18216
rect 2964 18207 3016 18216
rect 2964 18173 2973 18207
rect 2973 18173 3007 18207
rect 3007 18173 3016 18207
rect 2964 18164 3016 18173
rect 16028 18164 16080 18216
rect 15292 18096 15344 18148
rect 17040 18096 17092 18148
rect 18328 18164 18380 18216
rect 21088 18275 21140 18284
rect 14464 18071 14516 18080
rect 14464 18037 14473 18071
rect 14473 18037 14507 18071
rect 14507 18037 14516 18071
rect 14464 18028 14516 18037
rect 16672 18071 16724 18080
rect 16672 18037 16681 18071
rect 16681 18037 16715 18071
rect 16715 18037 16724 18071
rect 16672 18028 16724 18037
rect 16856 18071 16908 18080
rect 16856 18037 16874 18071
rect 16874 18037 16908 18071
rect 17592 18071 17644 18080
rect 16856 18028 16908 18037
rect 17592 18037 17601 18071
rect 17601 18037 17635 18071
rect 17635 18037 17644 18071
rect 17592 18028 17644 18037
rect 19432 18164 19484 18216
rect 21088 18241 21097 18275
rect 21097 18241 21131 18275
rect 21131 18241 21140 18275
rect 21088 18232 21140 18241
rect 21548 18232 21600 18284
rect 23480 18300 23532 18352
rect 25136 18343 25188 18352
rect 25136 18309 25170 18343
rect 25170 18309 25188 18343
rect 25136 18300 25188 18309
rect 26240 18300 26292 18352
rect 27804 18300 27856 18352
rect 34428 18300 34480 18352
rect 34888 18343 34940 18352
rect 34888 18309 34897 18343
rect 34897 18309 34931 18343
rect 34931 18309 34940 18343
rect 34888 18300 34940 18309
rect 35716 18300 35768 18352
rect 38384 18343 38436 18352
rect 23112 18232 23164 18284
rect 23572 18232 23624 18284
rect 25688 18232 25740 18284
rect 26056 18232 26108 18284
rect 26424 18232 26476 18284
rect 30196 18275 30248 18284
rect 30196 18241 30205 18275
rect 30205 18241 30239 18275
rect 30239 18241 30248 18275
rect 30196 18232 30248 18241
rect 32588 18232 32640 18284
rect 26976 18207 27028 18216
rect 26976 18173 26985 18207
rect 26985 18173 27019 18207
rect 27019 18173 27028 18207
rect 26976 18164 27028 18173
rect 30472 18207 30524 18216
rect 26240 18139 26292 18148
rect 26240 18105 26249 18139
rect 26249 18105 26283 18139
rect 26283 18105 26292 18139
rect 26240 18096 26292 18105
rect 19432 18071 19484 18080
rect 19432 18037 19441 18071
rect 19441 18037 19475 18071
rect 19475 18037 19484 18071
rect 19432 18028 19484 18037
rect 23756 18028 23808 18080
rect 26424 18028 26476 18080
rect 27712 18028 27764 18080
rect 30472 18173 30481 18207
rect 30481 18173 30515 18207
rect 30515 18173 30524 18207
rect 30472 18164 30524 18173
rect 33140 18275 33192 18284
rect 33140 18241 33149 18275
rect 33149 18241 33183 18275
rect 33183 18241 33192 18275
rect 34520 18275 34572 18284
rect 33140 18232 33192 18241
rect 34520 18241 34529 18275
rect 34529 18241 34563 18275
rect 34563 18241 34572 18275
rect 34520 18232 34572 18241
rect 34704 18275 34756 18284
rect 34704 18241 34711 18275
rect 34711 18241 34756 18275
rect 34704 18232 34756 18241
rect 33232 18164 33284 18216
rect 34980 18275 35032 18284
rect 34980 18241 34994 18275
rect 34994 18241 35028 18275
rect 35028 18241 35032 18275
rect 34980 18232 35032 18241
rect 35808 18232 35860 18284
rect 35992 18275 36044 18284
rect 35992 18241 36001 18275
rect 36001 18241 36035 18275
rect 36035 18241 36044 18275
rect 35992 18232 36044 18241
rect 38384 18309 38393 18343
rect 38393 18309 38427 18343
rect 38427 18309 38436 18343
rect 38384 18300 38436 18309
rect 43444 18377 43453 18411
rect 43453 18377 43487 18411
rect 43487 18377 43496 18411
rect 43444 18368 43496 18377
rect 37464 18275 37516 18284
rect 37464 18241 37473 18275
rect 37473 18241 37507 18275
rect 37507 18241 37516 18275
rect 37464 18232 37516 18241
rect 43352 18275 43404 18284
rect 43352 18241 43361 18275
rect 43361 18241 43395 18275
rect 43395 18241 43404 18275
rect 43352 18232 43404 18241
rect 35256 18164 35308 18216
rect 38752 18164 38804 18216
rect 39948 18207 40000 18216
rect 39948 18173 39957 18207
rect 39957 18173 39991 18207
rect 39991 18173 40000 18207
rect 39948 18164 40000 18173
rect 28540 18028 28592 18080
rect 28632 18028 28684 18080
rect 30656 18028 30708 18080
rect 35348 18028 35400 18080
rect 37280 18028 37332 18080
rect 37464 18071 37516 18080
rect 37464 18037 37473 18071
rect 37473 18037 37507 18071
rect 37507 18037 37516 18071
rect 37464 18028 37516 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 2872 17867 2924 17876
rect 2872 17833 2881 17867
rect 2881 17833 2915 17867
rect 2915 17833 2924 17867
rect 2872 17824 2924 17833
rect 16948 17824 17000 17876
rect 23296 17824 23348 17876
rect 26424 17824 26476 17876
rect 17316 17756 17368 17808
rect 26700 17756 26752 17808
rect 15568 17688 15620 17740
rect 1768 17620 1820 17672
rect 11704 17620 11756 17672
rect 17132 17688 17184 17740
rect 17868 17688 17920 17740
rect 26240 17731 26292 17740
rect 26240 17697 26249 17731
rect 26249 17697 26283 17731
rect 26283 17697 26292 17731
rect 26240 17688 26292 17697
rect 26976 17688 27028 17740
rect 15200 17595 15252 17604
rect 15200 17561 15218 17595
rect 15218 17561 15252 17595
rect 15200 17552 15252 17561
rect 17040 17620 17092 17672
rect 17500 17620 17552 17672
rect 17408 17484 17460 17536
rect 19432 17620 19484 17672
rect 20352 17620 20404 17672
rect 23480 17620 23532 17672
rect 26056 17663 26108 17672
rect 26056 17629 26065 17663
rect 26065 17629 26099 17663
rect 26099 17629 26108 17663
rect 26056 17620 26108 17629
rect 24860 17552 24912 17604
rect 25964 17552 26016 17604
rect 30472 17824 30524 17876
rect 28540 17756 28592 17808
rect 29552 17731 29604 17740
rect 29552 17697 29561 17731
rect 29561 17697 29595 17731
rect 29595 17697 29604 17731
rect 29552 17688 29604 17697
rect 33140 17824 33192 17876
rect 34704 17824 34756 17876
rect 35716 17824 35768 17876
rect 35992 17824 36044 17876
rect 27712 17620 27764 17672
rect 28632 17620 28684 17672
rect 28080 17595 28132 17604
rect 19432 17484 19484 17536
rect 27252 17484 27304 17536
rect 28080 17561 28089 17595
rect 28089 17561 28123 17595
rect 28123 17561 28132 17595
rect 28080 17552 28132 17561
rect 29460 17552 29512 17604
rect 30564 17552 30616 17604
rect 28816 17484 28868 17536
rect 31024 17484 31076 17536
rect 33324 17756 33376 17808
rect 32588 17688 32640 17740
rect 34520 17688 34572 17740
rect 34796 17731 34848 17740
rect 34796 17697 34805 17731
rect 34805 17697 34839 17731
rect 34839 17697 34848 17731
rect 34796 17688 34848 17697
rect 33232 17663 33284 17672
rect 33232 17629 33241 17663
rect 33241 17629 33275 17663
rect 33275 17629 33284 17663
rect 33232 17620 33284 17629
rect 34612 17620 34664 17672
rect 34888 17663 34940 17672
rect 34888 17629 34897 17663
rect 34897 17629 34931 17663
rect 34931 17629 34940 17663
rect 34888 17620 34940 17629
rect 35348 17620 35400 17672
rect 33140 17595 33192 17604
rect 33140 17561 33149 17595
rect 33149 17561 33183 17595
rect 33183 17561 33192 17595
rect 33140 17552 33192 17561
rect 38108 17688 38160 17740
rect 43628 17824 43680 17876
rect 42616 17756 42668 17808
rect 42984 17688 43036 17740
rect 35808 17663 35860 17672
rect 35808 17629 35817 17663
rect 35817 17629 35851 17663
rect 35851 17629 35860 17663
rect 35808 17620 35860 17629
rect 37004 17663 37056 17672
rect 37004 17629 37013 17663
rect 37013 17629 37047 17663
rect 37047 17629 37056 17663
rect 37004 17620 37056 17629
rect 42984 17552 43036 17604
rect 43168 17552 43220 17604
rect 35348 17484 35400 17536
rect 35716 17484 35768 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 15200 17280 15252 17332
rect 1768 17187 1820 17196
rect 1768 17153 1777 17187
rect 1777 17153 1811 17187
rect 1811 17153 1820 17187
rect 1768 17144 1820 17153
rect 14464 17144 14516 17196
rect 15568 17187 15620 17196
rect 1952 17119 2004 17128
rect 1952 17085 1961 17119
rect 1961 17085 1995 17119
rect 1995 17085 2004 17119
rect 1952 17076 2004 17085
rect 2780 17119 2832 17128
rect 2780 17085 2789 17119
rect 2789 17085 2823 17119
rect 2823 17085 2832 17119
rect 2780 17076 2832 17085
rect 15568 17153 15577 17187
rect 15577 17153 15611 17187
rect 15611 17153 15620 17187
rect 15568 17144 15620 17153
rect 16212 17144 16264 17196
rect 16764 17144 16816 17196
rect 16948 17187 17000 17196
rect 16948 17153 16957 17187
rect 16957 17153 16991 17187
rect 16991 17153 17000 17187
rect 16948 17144 17000 17153
rect 17132 17144 17184 17196
rect 17408 17280 17460 17332
rect 20628 17280 20680 17332
rect 23296 17280 23348 17332
rect 24860 17323 24912 17332
rect 23756 17255 23808 17264
rect 17500 17144 17552 17196
rect 19432 17187 19484 17196
rect 15292 16940 15344 16992
rect 17868 17076 17920 17128
rect 19432 17153 19441 17187
rect 19441 17153 19475 17187
rect 19475 17153 19484 17187
rect 19432 17144 19484 17153
rect 19616 17187 19668 17196
rect 19616 17153 19625 17187
rect 19625 17153 19659 17187
rect 19659 17153 19668 17187
rect 19616 17144 19668 17153
rect 20076 17144 20128 17196
rect 23756 17221 23790 17255
rect 23790 17221 23808 17255
rect 23756 17212 23808 17221
rect 20536 17144 20588 17196
rect 21824 17187 21876 17196
rect 21824 17153 21833 17187
rect 21833 17153 21867 17187
rect 21867 17153 21876 17187
rect 21824 17144 21876 17153
rect 22744 17144 22796 17196
rect 19524 17076 19576 17128
rect 20352 17076 20404 17128
rect 23296 17076 23348 17128
rect 23480 17119 23532 17128
rect 23480 17085 23489 17119
rect 23489 17085 23523 17119
rect 23523 17085 23532 17119
rect 23480 17076 23532 17085
rect 24860 17289 24869 17323
rect 24869 17289 24903 17323
rect 24903 17289 24912 17323
rect 24860 17280 24912 17289
rect 29644 17280 29696 17332
rect 30196 17280 30248 17332
rect 30564 17323 30616 17332
rect 30564 17289 30573 17323
rect 30573 17289 30607 17323
rect 30607 17289 30616 17323
rect 30564 17280 30616 17289
rect 25320 17255 25372 17264
rect 25320 17221 25329 17255
rect 25329 17221 25363 17255
rect 25363 17221 25372 17255
rect 25320 17212 25372 17221
rect 27620 17212 27672 17264
rect 29460 17212 29512 17264
rect 34888 17212 34940 17264
rect 35716 17212 35768 17264
rect 24768 17144 24820 17196
rect 28080 17144 28132 17196
rect 28816 17187 28868 17196
rect 28816 17153 28850 17187
rect 28850 17153 28868 17187
rect 28816 17144 28868 17153
rect 29736 17144 29788 17196
rect 32864 17187 32916 17196
rect 32864 17153 32873 17187
rect 32873 17153 32907 17187
rect 32907 17153 32916 17187
rect 32864 17144 32916 17153
rect 33048 17187 33100 17196
rect 33048 17153 33057 17187
rect 33057 17153 33091 17187
rect 33091 17153 33100 17187
rect 33048 17144 33100 17153
rect 27068 17119 27120 17128
rect 27068 17085 27077 17119
rect 27077 17085 27111 17119
rect 27111 17085 27120 17119
rect 27068 17076 27120 17085
rect 28540 17119 28592 17128
rect 28540 17085 28549 17119
rect 28549 17085 28583 17119
rect 28583 17085 28592 17119
rect 28540 17076 28592 17085
rect 37004 17144 37056 17196
rect 37464 17187 37516 17196
rect 37464 17153 37473 17187
rect 37473 17153 37507 17187
rect 37507 17153 37516 17187
rect 37464 17144 37516 17153
rect 42984 17144 43036 17196
rect 21180 17008 21232 17060
rect 16948 16940 17000 16992
rect 20260 16940 20312 16992
rect 22008 16983 22060 16992
rect 22008 16949 22017 16983
rect 22017 16949 22051 16983
rect 22051 16949 22060 16983
rect 22008 16940 22060 16949
rect 26332 17008 26384 17060
rect 27620 17008 27672 17060
rect 35900 17008 35952 17060
rect 23848 16940 23900 16992
rect 33784 16940 33836 16992
rect 38936 16940 38988 16992
rect 43996 16940 44048 16992
rect 44180 16983 44232 16992
rect 44180 16949 44189 16983
rect 44189 16949 44223 16983
rect 44223 16949 44232 16983
rect 44180 16940 44232 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 1952 16736 2004 16788
rect 15752 16779 15804 16788
rect 15752 16745 15761 16779
rect 15761 16745 15795 16779
rect 15795 16745 15804 16779
rect 15752 16736 15804 16745
rect 16028 16736 16080 16788
rect 16672 16736 16724 16788
rect 17500 16736 17552 16788
rect 23112 16779 23164 16788
rect 23112 16745 23121 16779
rect 23121 16745 23155 16779
rect 23155 16745 23164 16779
rect 23112 16736 23164 16745
rect 1676 16532 1728 16584
rect 6184 16600 6236 16652
rect 15292 16643 15344 16652
rect 15292 16609 15301 16643
rect 15301 16609 15335 16643
rect 15335 16609 15344 16643
rect 15292 16600 15344 16609
rect 15844 16668 15896 16720
rect 20812 16711 20864 16720
rect 20812 16677 20821 16711
rect 20821 16677 20855 16711
rect 20855 16677 20864 16711
rect 20812 16668 20864 16677
rect 22744 16711 22796 16720
rect 22744 16677 22753 16711
rect 22753 16677 22787 16711
rect 22787 16677 22796 16711
rect 22744 16668 22796 16677
rect 23296 16668 23348 16720
rect 15936 16600 15988 16652
rect 17316 16643 17368 16652
rect 12900 16396 12952 16448
rect 16028 16532 16080 16584
rect 15752 16464 15804 16516
rect 16672 16532 16724 16584
rect 16948 16532 17000 16584
rect 17316 16609 17325 16643
rect 17325 16609 17359 16643
rect 17359 16609 17368 16643
rect 17316 16600 17368 16609
rect 19524 16643 19576 16652
rect 19524 16609 19533 16643
rect 19533 16609 19567 16643
rect 19567 16609 19576 16643
rect 19524 16600 19576 16609
rect 20996 16600 21048 16652
rect 23940 16600 23992 16652
rect 17408 16532 17460 16584
rect 19248 16575 19300 16584
rect 19248 16541 19257 16575
rect 19257 16541 19291 16575
rect 19291 16541 19300 16575
rect 19248 16532 19300 16541
rect 21640 16575 21692 16584
rect 21640 16541 21649 16575
rect 21649 16541 21683 16575
rect 21683 16541 21692 16575
rect 21640 16532 21692 16541
rect 17684 16464 17736 16516
rect 19616 16464 19668 16516
rect 22192 16464 22244 16516
rect 24768 16600 24820 16652
rect 33048 16668 33100 16720
rect 31024 16643 31076 16652
rect 31024 16609 31033 16643
rect 31033 16609 31067 16643
rect 31067 16609 31076 16643
rect 31024 16600 31076 16609
rect 33784 16643 33836 16652
rect 33784 16609 33793 16643
rect 33793 16609 33827 16643
rect 33827 16609 33836 16643
rect 33784 16600 33836 16609
rect 34060 16643 34112 16652
rect 34060 16609 34069 16643
rect 34069 16609 34103 16643
rect 34103 16609 34112 16643
rect 34060 16600 34112 16609
rect 35348 16600 35400 16652
rect 37464 16600 37516 16652
rect 43996 16643 44048 16652
rect 43996 16609 44005 16643
rect 44005 16609 44039 16643
rect 44039 16609 44048 16643
rect 43996 16600 44048 16609
rect 44180 16643 44232 16652
rect 44180 16609 44189 16643
rect 44189 16609 44223 16643
rect 44223 16609 44232 16643
rect 44180 16600 44232 16609
rect 24400 16575 24452 16584
rect 24400 16541 24409 16575
rect 24409 16541 24443 16575
rect 24443 16541 24452 16575
rect 24400 16532 24452 16541
rect 24952 16532 25004 16584
rect 30748 16532 30800 16584
rect 34888 16532 34940 16584
rect 37004 16532 37056 16584
rect 37924 16575 37976 16584
rect 37924 16541 37933 16575
rect 37933 16541 37967 16575
rect 37967 16541 37976 16575
rect 37924 16532 37976 16541
rect 42340 16575 42392 16584
rect 42340 16541 42349 16575
rect 42349 16541 42383 16575
rect 42383 16541 42392 16575
rect 42340 16532 42392 16541
rect 18052 16396 18104 16448
rect 18696 16439 18748 16448
rect 18696 16405 18705 16439
rect 18705 16405 18739 16439
rect 18739 16405 18748 16439
rect 18696 16396 18748 16405
rect 19248 16396 19300 16448
rect 21088 16396 21140 16448
rect 32956 16464 33008 16516
rect 35808 16507 35860 16516
rect 23480 16396 23532 16448
rect 33232 16396 33284 16448
rect 35808 16473 35817 16507
rect 35817 16473 35851 16507
rect 35851 16473 35860 16507
rect 35808 16464 35860 16473
rect 40132 16464 40184 16516
rect 37280 16396 37332 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 15660 16192 15712 16244
rect 17684 16192 17736 16244
rect 17868 16235 17920 16244
rect 17868 16201 17877 16235
rect 17877 16201 17911 16235
rect 17911 16201 17920 16235
rect 17868 16192 17920 16201
rect 16764 16124 16816 16176
rect 1676 16099 1728 16108
rect 1676 16065 1685 16099
rect 1685 16065 1719 16099
rect 1719 16065 1728 16099
rect 1676 16056 1728 16065
rect 12900 16099 12952 16108
rect 12900 16065 12909 16099
rect 12909 16065 12943 16099
rect 12943 16065 12952 16099
rect 12900 16056 12952 16065
rect 15292 16056 15344 16108
rect 16028 16056 16080 16108
rect 2228 15988 2280 16040
rect 2780 16031 2832 16040
rect 2780 15997 2789 16031
rect 2789 15997 2823 16031
rect 2823 15997 2832 16031
rect 2780 15988 2832 15997
rect 13176 15988 13228 16040
rect 14740 16031 14792 16040
rect 14740 15997 14749 16031
rect 14749 15997 14783 16031
rect 14783 15997 14792 16031
rect 14740 15988 14792 15997
rect 15660 16031 15712 16040
rect 15660 15997 15669 16031
rect 15669 15997 15703 16031
rect 15703 15997 15712 16031
rect 15660 15988 15712 15997
rect 15844 16031 15896 16040
rect 15844 15997 15853 16031
rect 15853 15997 15887 16031
rect 15887 15997 15896 16031
rect 15844 15988 15896 15997
rect 16672 15988 16724 16040
rect 17132 16102 17184 16108
rect 17132 16068 17141 16102
rect 17141 16068 17175 16102
rect 17175 16068 17184 16102
rect 17132 16056 17184 16068
rect 17408 16056 17460 16108
rect 17592 16056 17644 16108
rect 3424 15852 3476 15904
rect 12532 15852 12584 15904
rect 16948 15920 17000 15972
rect 16580 15852 16632 15904
rect 16764 15852 16816 15904
rect 18512 16056 18564 16108
rect 19340 15963 19392 15972
rect 19340 15929 19349 15963
rect 19349 15929 19383 15963
rect 19383 15929 19392 15963
rect 19340 15920 19392 15929
rect 20260 16099 20312 16108
rect 20260 16065 20269 16099
rect 20269 16065 20303 16099
rect 20303 16065 20312 16099
rect 20260 16056 20312 16065
rect 22376 16192 22428 16244
rect 32956 16192 33008 16244
rect 33232 16235 33284 16244
rect 33232 16201 33241 16235
rect 33241 16201 33275 16235
rect 33275 16201 33284 16235
rect 33232 16192 33284 16201
rect 34888 16192 34940 16244
rect 21548 16124 21600 16176
rect 20812 16056 20864 16108
rect 22008 16056 22060 16108
rect 26516 16124 26568 16176
rect 27620 16124 27672 16176
rect 32864 16167 32916 16176
rect 32864 16133 32873 16167
rect 32873 16133 32907 16167
rect 32907 16133 32916 16167
rect 32864 16124 32916 16133
rect 33048 16167 33100 16176
rect 33048 16133 33057 16167
rect 33057 16133 33091 16167
rect 33091 16133 33100 16167
rect 33048 16124 33100 16133
rect 23848 15988 23900 16040
rect 20996 15920 21048 15972
rect 21088 15920 21140 15972
rect 26240 15920 26292 15972
rect 27068 16056 27120 16108
rect 27252 16056 27304 16108
rect 28540 16099 28592 16108
rect 21640 15852 21692 15904
rect 22560 15852 22612 15904
rect 23480 15852 23532 15904
rect 27068 15852 27120 15904
rect 27620 15895 27672 15904
rect 27620 15861 27629 15895
rect 27629 15861 27663 15895
rect 27663 15861 27672 15895
rect 27620 15852 27672 15861
rect 28540 16065 28549 16099
rect 28549 16065 28583 16099
rect 28583 16065 28592 16099
rect 28540 16056 28592 16065
rect 37372 16124 37424 16176
rect 33784 16056 33836 16108
rect 35808 16056 35860 16108
rect 36268 15988 36320 16040
rect 38108 16099 38160 16108
rect 38108 16065 38117 16099
rect 38117 16065 38151 16099
rect 38151 16065 38160 16099
rect 38108 16056 38160 16065
rect 43260 16056 43312 16108
rect 29552 15852 29604 15904
rect 29920 15895 29972 15904
rect 29920 15861 29929 15895
rect 29929 15861 29963 15895
rect 29963 15861 29972 15895
rect 29920 15852 29972 15861
rect 37464 15852 37516 15904
rect 37924 15895 37976 15904
rect 37924 15861 37933 15895
rect 37933 15861 37967 15895
rect 37967 15861 37976 15895
rect 37924 15852 37976 15861
rect 42708 15895 42760 15904
rect 42708 15861 42717 15895
rect 42717 15861 42751 15895
rect 42751 15861 42760 15895
rect 42708 15852 42760 15861
rect 43444 15895 43496 15904
rect 43444 15861 43453 15895
rect 43453 15861 43487 15895
rect 43487 15861 43496 15895
rect 43444 15852 43496 15861
rect 44180 15895 44232 15904
rect 44180 15861 44189 15895
rect 44189 15861 44223 15895
rect 44223 15861 44232 15895
rect 44180 15852 44232 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 2228 15691 2280 15700
rect 2228 15657 2237 15691
rect 2237 15657 2271 15691
rect 2271 15657 2280 15691
rect 2228 15648 2280 15657
rect 13176 15691 13228 15700
rect 13176 15657 13185 15691
rect 13185 15657 13219 15691
rect 13219 15657 13228 15691
rect 13176 15648 13228 15657
rect 15660 15648 15712 15700
rect 15936 15648 15988 15700
rect 16672 15648 16724 15700
rect 19984 15648 20036 15700
rect 20812 15648 20864 15700
rect 21180 15691 21232 15700
rect 21180 15657 21189 15691
rect 21189 15657 21223 15691
rect 21223 15657 21232 15691
rect 21180 15648 21232 15657
rect 22192 15691 22244 15700
rect 22192 15657 22201 15691
rect 22201 15657 22235 15691
rect 22235 15657 22244 15691
rect 22192 15648 22244 15657
rect 22560 15691 22612 15700
rect 22560 15657 22569 15691
rect 22569 15657 22603 15691
rect 22603 15657 22612 15691
rect 22560 15648 22612 15657
rect 22744 15648 22796 15700
rect 26516 15691 26568 15700
rect 17316 15580 17368 15632
rect 21824 15580 21876 15632
rect 26516 15657 26525 15691
rect 26525 15657 26559 15691
rect 26559 15657 26568 15691
rect 26516 15648 26568 15657
rect 16672 15555 16724 15564
rect 16672 15521 16681 15555
rect 16681 15521 16715 15555
rect 16715 15521 16724 15555
rect 21088 15555 21140 15564
rect 16672 15512 16724 15521
rect 21088 15521 21097 15555
rect 21097 15521 21131 15555
rect 21131 15521 21140 15555
rect 21088 15512 21140 15521
rect 2412 15444 2464 15496
rect 3424 15444 3476 15496
rect 13544 15444 13596 15496
rect 16580 15444 16632 15496
rect 17592 15444 17644 15496
rect 19248 15444 19300 15496
rect 20536 15487 20588 15496
rect 20536 15453 20545 15487
rect 20545 15453 20579 15487
rect 20579 15453 20588 15487
rect 20536 15444 20588 15453
rect 21548 15512 21600 15564
rect 22928 15512 22980 15564
rect 22284 15487 22336 15496
rect 22284 15453 22293 15487
rect 22293 15453 22327 15487
rect 22327 15453 22336 15487
rect 36084 15623 36136 15632
rect 36084 15589 36093 15623
rect 36093 15589 36127 15623
rect 36127 15589 36136 15623
rect 36084 15580 36136 15589
rect 23296 15555 23348 15564
rect 23296 15521 23305 15555
rect 23305 15521 23339 15555
rect 23339 15521 23348 15555
rect 23296 15512 23348 15521
rect 22284 15444 22336 15453
rect 29644 15487 29696 15496
rect 29644 15453 29653 15487
rect 29653 15453 29687 15487
rect 29687 15453 29696 15487
rect 29644 15444 29696 15453
rect 31024 15444 31076 15496
rect 31208 15487 31260 15496
rect 31208 15453 31242 15487
rect 31242 15453 31260 15487
rect 31208 15444 31260 15453
rect 27528 15376 27580 15428
rect 27620 15419 27672 15428
rect 27620 15385 27638 15419
rect 27638 15385 27672 15419
rect 27620 15376 27672 15385
rect 32956 15487 33008 15496
rect 32956 15453 32965 15487
rect 32965 15453 32999 15487
rect 32999 15453 33008 15487
rect 32956 15444 33008 15453
rect 33232 15444 33284 15496
rect 35808 15444 35860 15496
rect 37372 15512 37424 15564
rect 42616 15555 42668 15564
rect 42616 15521 42625 15555
rect 42625 15521 42659 15555
rect 42659 15521 42668 15555
rect 42616 15512 42668 15521
rect 44180 15555 44232 15564
rect 44180 15521 44189 15555
rect 44189 15521 44223 15555
rect 44223 15521 44232 15555
rect 44180 15512 44232 15521
rect 37740 15444 37792 15496
rect 38936 15487 38988 15496
rect 38936 15453 38945 15487
rect 38945 15453 38979 15487
rect 38979 15453 38988 15487
rect 38936 15444 38988 15453
rect 19248 15308 19300 15360
rect 24400 15308 24452 15360
rect 25964 15308 26016 15360
rect 29736 15351 29788 15360
rect 29736 15317 29745 15351
rect 29745 15317 29779 15351
rect 29779 15317 29788 15351
rect 29736 15308 29788 15317
rect 32312 15351 32364 15360
rect 32312 15317 32321 15351
rect 32321 15317 32355 15351
rect 32355 15317 32364 15351
rect 32312 15308 32364 15317
rect 33140 15351 33192 15360
rect 33140 15317 33149 15351
rect 33149 15317 33183 15351
rect 33183 15317 33192 15351
rect 33140 15308 33192 15317
rect 33600 15308 33652 15360
rect 36820 15351 36872 15360
rect 36820 15317 36829 15351
rect 36829 15317 36863 15351
rect 36863 15317 36872 15351
rect 36820 15308 36872 15317
rect 37280 15376 37332 15428
rect 43996 15419 44048 15428
rect 43996 15385 44005 15419
rect 44005 15385 44039 15419
rect 44039 15385 44048 15419
rect 43996 15376 44048 15385
rect 37372 15308 37424 15360
rect 39028 15351 39080 15360
rect 39028 15317 39037 15351
rect 39037 15317 39071 15351
rect 39071 15317 39080 15351
rect 39028 15308 39080 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 15844 15104 15896 15156
rect 18144 15104 18196 15156
rect 23664 15104 23716 15156
rect 19064 15036 19116 15088
rect 13544 14968 13596 15020
rect 18512 15011 18564 15020
rect 18512 14977 18521 15011
rect 18521 14977 18555 15011
rect 18555 14977 18564 15011
rect 18512 14968 18564 14977
rect 19984 14968 20036 15020
rect 20904 14968 20956 15020
rect 21180 15036 21232 15088
rect 22744 15036 22796 15088
rect 22928 15036 22980 15088
rect 23940 15079 23992 15088
rect 23940 15045 23949 15079
rect 23949 15045 23983 15079
rect 23983 15045 23992 15079
rect 23940 15036 23992 15045
rect 25780 15036 25832 15088
rect 22192 14968 22244 15020
rect 24216 14968 24268 15020
rect 25964 15036 26016 15088
rect 29552 15104 29604 15156
rect 26240 15011 26292 15020
rect 26240 14977 26249 15011
rect 26249 14977 26283 15011
rect 26283 14977 26292 15011
rect 26240 14968 26292 14977
rect 26976 14968 27028 15020
rect 30840 15036 30892 15088
rect 27436 14968 27488 15020
rect 33232 15036 33284 15088
rect 18788 14900 18840 14952
rect 23296 14900 23348 14952
rect 27068 14943 27120 14952
rect 27068 14909 27077 14943
rect 27077 14909 27111 14943
rect 27111 14909 27120 14943
rect 27068 14900 27120 14909
rect 14280 14764 14332 14816
rect 18052 14764 18104 14816
rect 19248 14764 19300 14816
rect 19432 14764 19484 14816
rect 19708 14807 19760 14816
rect 19708 14773 19717 14807
rect 19717 14773 19751 14807
rect 19751 14773 19760 14807
rect 19708 14764 19760 14773
rect 21088 14764 21140 14816
rect 22836 14832 22888 14884
rect 23848 14832 23900 14884
rect 26424 14832 26476 14884
rect 28448 14900 28500 14952
rect 30196 14832 30248 14884
rect 33140 14968 33192 15020
rect 33600 15011 33652 15020
rect 33600 14977 33609 15011
rect 33609 14977 33643 15011
rect 33643 14977 33652 15011
rect 33600 14968 33652 14977
rect 34060 14968 34112 15020
rect 32220 14832 32272 14884
rect 32956 14832 33008 14884
rect 43996 15104 44048 15156
rect 36084 15036 36136 15088
rect 37280 15036 37332 15088
rect 35992 14968 36044 15020
rect 36268 15011 36320 15020
rect 36268 14977 36277 15011
rect 36277 14977 36311 15011
rect 36311 14977 36320 15011
rect 36268 14968 36320 14977
rect 35532 14943 35584 14952
rect 35532 14909 35541 14943
rect 35541 14909 35575 14943
rect 35575 14909 35584 14943
rect 35532 14900 35584 14909
rect 36452 15011 36504 15020
rect 36452 14977 36461 15011
rect 36461 14977 36495 15011
rect 36495 14977 36504 15011
rect 36452 14968 36504 14977
rect 36820 14968 36872 15020
rect 37464 14968 37516 15020
rect 38936 15011 38988 15020
rect 38936 14977 38946 15011
rect 38946 14977 38980 15011
rect 38980 14977 38988 15011
rect 38936 14968 38988 14977
rect 36544 14832 36596 14884
rect 37372 14900 37424 14952
rect 37464 14832 37516 14884
rect 37648 14832 37700 14884
rect 37924 14900 37976 14952
rect 38384 14900 38436 14952
rect 43904 14968 43956 15020
rect 26976 14764 27028 14816
rect 28356 14764 28408 14816
rect 30012 14764 30064 14816
rect 30656 14764 30708 14816
rect 32404 14807 32456 14816
rect 32404 14773 32413 14807
rect 32413 14773 32447 14807
rect 32447 14773 32456 14807
rect 32404 14764 32456 14773
rect 34428 14764 34480 14816
rect 35348 14764 35400 14816
rect 37280 14764 37332 14816
rect 38292 14764 38344 14816
rect 38936 14764 38988 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 18512 14560 18564 14612
rect 22008 14560 22060 14612
rect 22928 14560 22980 14612
rect 26240 14560 26292 14612
rect 27068 14603 27120 14612
rect 27068 14569 27077 14603
rect 27077 14569 27111 14603
rect 27111 14569 27120 14603
rect 27068 14560 27120 14569
rect 27436 14603 27488 14612
rect 27436 14569 27445 14603
rect 27445 14569 27479 14603
rect 27479 14569 27488 14603
rect 27436 14560 27488 14569
rect 30012 14603 30064 14612
rect 30012 14569 30021 14603
rect 30021 14569 30055 14603
rect 30055 14569 30064 14603
rect 30012 14560 30064 14569
rect 30196 14603 30248 14612
rect 30196 14569 30205 14603
rect 30205 14569 30239 14603
rect 30239 14569 30248 14603
rect 30196 14560 30248 14569
rect 35992 14560 36044 14612
rect 36544 14560 36596 14612
rect 43904 14560 43956 14612
rect 22192 14492 22244 14544
rect 26148 14535 26200 14544
rect 26148 14501 26157 14535
rect 26157 14501 26191 14535
rect 26191 14501 26200 14535
rect 26148 14492 26200 14501
rect 14280 14467 14332 14476
rect 14280 14433 14289 14467
rect 14289 14433 14323 14467
rect 14323 14433 14332 14467
rect 14280 14424 14332 14433
rect 2044 14356 2096 14408
rect 9220 14356 9272 14408
rect 14004 14356 14056 14408
rect 15936 14331 15988 14340
rect 15936 14297 15945 14331
rect 15945 14297 15979 14331
rect 15979 14297 15988 14331
rect 15936 14288 15988 14297
rect 18052 14399 18104 14408
rect 18052 14365 18061 14399
rect 18061 14365 18095 14399
rect 18095 14365 18104 14399
rect 18788 14424 18840 14476
rect 22008 14424 22060 14476
rect 25780 14467 25832 14476
rect 25780 14433 25789 14467
rect 25789 14433 25823 14467
rect 25823 14433 25832 14467
rect 25780 14424 25832 14433
rect 29920 14467 29972 14476
rect 29920 14433 29929 14467
rect 29929 14433 29963 14467
rect 29963 14433 29972 14467
rect 29920 14424 29972 14433
rect 30196 14424 30248 14476
rect 18328 14399 18380 14408
rect 18052 14356 18104 14365
rect 18328 14365 18337 14399
rect 18337 14365 18371 14399
rect 18371 14365 18380 14399
rect 18328 14356 18380 14365
rect 19340 14356 19392 14408
rect 19708 14356 19760 14408
rect 18144 14288 18196 14340
rect 21916 14288 21968 14340
rect 22100 14288 22152 14340
rect 22284 14288 22336 14340
rect 22652 14399 22704 14408
rect 22652 14365 22661 14399
rect 22661 14365 22695 14399
rect 22695 14365 22704 14399
rect 22652 14356 22704 14365
rect 25964 14399 26016 14408
rect 25964 14365 25973 14399
rect 25973 14365 26007 14399
rect 26007 14365 26016 14399
rect 25964 14356 26016 14365
rect 26976 14399 27028 14408
rect 26976 14365 26985 14399
rect 26985 14365 27019 14399
rect 27019 14365 27028 14399
rect 26976 14356 27028 14365
rect 30104 14356 30156 14408
rect 31576 14356 31628 14408
rect 32404 14356 32456 14408
rect 36452 14492 36504 14544
rect 35348 14399 35400 14408
rect 35348 14365 35357 14399
rect 35357 14365 35391 14399
rect 35391 14365 35400 14399
rect 35348 14356 35400 14365
rect 35532 14467 35584 14476
rect 35532 14433 35541 14467
rect 35541 14433 35575 14467
rect 35575 14433 35584 14467
rect 35532 14424 35584 14433
rect 38200 14492 38252 14544
rect 36820 14424 36872 14476
rect 37464 14424 37516 14476
rect 37740 14467 37792 14476
rect 37740 14433 37749 14467
rect 37749 14433 37783 14467
rect 37783 14433 37792 14467
rect 37740 14424 37792 14433
rect 39028 14424 39080 14476
rect 42708 14424 42760 14476
rect 44088 14467 44140 14476
rect 44088 14433 44097 14467
rect 44097 14433 44131 14467
rect 44131 14433 44140 14467
rect 44088 14424 44140 14433
rect 37280 14356 37332 14408
rect 38016 14356 38068 14408
rect 38568 14356 38620 14408
rect 25688 14331 25740 14340
rect 25688 14297 25697 14331
rect 25697 14297 25731 14331
rect 25731 14297 25740 14331
rect 25688 14288 25740 14297
rect 29644 14288 29696 14340
rect 38936 14288 38988 14340
rect 43444 14288 43496 14340
rect 2228 14220 2280 14272
rect 20720 14220 20772 14272
rect 21640 14263 21692 14272
rect 21640 14229 21649 14263
rect 21649 14229 21683 14263
rect 21683 14229 21692 14263
rect 21640 14220 21692 14229
rect 23296 14263 23348 14272
rect 23296 14229 23305 14263
rect 23305 14229 23339 14263
rect 23339 14229 23348 14263
rect 23296 14220 23348 14229
rect 33508 14263 33560 14272
rect 33508 14229 33517 14263
rect 33517 14229 33551 14263
rect 33551 14229 33560 14263
rect 33508 14220 33560 14229
rect 34336 14220 34388 14272
rect 36544 14263 36596 14272
rect 36544 14229 36553 14263
rect 36553 14229 36587 14263
rect 36587 14229 36596 14263
rect 36544 14220 36596 14229
rect 38568 14220 38620 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 14004 14059 14056 14068
rect 14004 14025 14013 14059
rect 14013 14025 14047 14059
rect 14047 14025 14056 14059
rect 14004 14016 14056 14025
rect 17960 14016 18012 14068
rect 21180 14059 21232 14068
rect 21180 14025 21189 14059
rect 21189 14025 21223 14059
rect 21223 14025 21232 14059
rect 21180 14016 21232 14025
rect 22652 14016 22704 14068
rect 25872 14016 25924 14068
rect 29644 14059 29696 14068
rect 29644 14025 29653 14059
rect 29653 14025 29687 14059
rect 29687 14025 29696 14059
rect 29644 14016 29696 14025
rect 30104 14059 30156 14068
rect 30104 14025 30113 14059
rect 30113 14025 30147 14059
rect 30147 14025 30156 14059
rect 30104 14016 30156 14025
rect 33232 14016 33284 14068
rect 34336 14059 34388 14068
rect 34336 14025 34345 14059
rect 34345 14025 34379 14059
rect 34379 14025 34388 14059
rect 34336 14016 34388 14025
rect 34428 14059 34480 14068
rect 34428 14025 34437 14059
rect 34437 14025 34471 14059
rect 34471 14025 34480 14059
rect 34428 14016 34480 14025
rect 36544 14016 36596 14068
rect 38200 14016 38252 14068
rect 38384 14016 38436 14068
rect 38568 14016 38620 14068
rect 2228 13991 2280 14000
rect 2228 13957 2237 13991
rect 2237 13957 2271 13991
rect 2271 13957 2280 13991
rect 2228 13948 2280 13957
rect 2044 13923 2096 13932
rect 2044 13889 2053 13923
rect 2053 13889 2087 13923
rect 2087 13889 2096 13923
rect 2044 13880 2096 13889
rect 18052 13948 18104 14000
rect 19064 13948 19116 14000
rect 16672 13923 16724 13932
rect 16672 13889 16681 13923
rect 16681 13889 16715 13923
rect 16715 13889 16724 13923
rect 16672 13880 16724 13889
rect 16948 13923 17000 13932
rect 16948 13889 16982 13923
rect 16982 13889 17000 13923
rect 16948 13880 17000 13889
rect 2780 13855 2832 13864
rect 2780 13821 2789 13855
rect 2789 13821 2823 13855
rect 2823 13821 2832 13855
rect 2780 13812 2832 13821
rect 18328 13812 18380 13864
rect 19064 13855 19116 13864
rect 19064 13821 19073 13855
rect 19073 13821 19107 13855
rect 19107 13821 19116 13855
rect 19432 13880 19484 13932
rect 21824 13948 21876 14000
rect 21272 13923 21324 13932
rect 21272 13889 21281 13923
rect 21281 13889 21315 13923
rect 21315 13889 21324 13923
rect 21272 13880 21324 13889
rect 22836 13948 22888 14000
rect 29736 13948 29788 14000
rect 37096 13948 37148 14000
rect 37740 13948 37792 14000
rect 38476 13948 38528 14000
rect 38844 13991 38896 14000
rect 22284 13880 22336 13932
rect 26424 13880 26476 13932
rect 27528 13880 27580 13932
rect 28356 13880 28408 13932
rect 30196 13880 30248 13932
rect 19064 13812 19116 13821
rect 22100 13812 22152 13864
rect 29276 13812 29328 13864
rect 32220 13923 32272 13932
rect 32220 13889 32229 13923
rect 32229 13889 32263 13923
rect 32263 13889 32272 13923
rect 32220 13880 32272 13889
rect 32312 13880 32364 13932
rect 35808 13880 35860 13932
rect 37372 13880 37424 13932
rect 38844 13957 38853 13991
rect 38853 13957 38887 13991
rect 38887 13957 38896 13991
rect 38844 13948 38896 13957
rect 31484 13855 31536 13864
rect 31484 13821 31493 13855
rect 31493 13821 31527 13855
rect 31527 13821 31536 13855
rect 31484 13812 31536 13821
rect 33508 13812 33560 13864
rect 34428 13812 34480 13864
rect 36452 13812 36504 13864
rect 37096 13812 37148 13864
rect 37556 13812 37608 13864
rect 43720 13880 43772 13932
rect 24584 13744 24636 13796
rect 25504 13744 25556 13796
rect 27528 13787 27580 13796
rect 27528 13753 27537 13787
rect 27537 13753 27571 13787
rect 27571 13753 27580 13787
rect 27528 13744 27580 13753
rect 19248 13676 19300 13728
rect 27804 13676 27856 13728
rect 33968 13719 34020 13728
rect 33968 13685 33977 13719
rect 33977 13685 34011 13719
rect 34011 13685 34020 13719
rect 33968 13676 34020 13685
rect 37280 13719 37332 13728
rect 37280 13685 37289 13719
rect 37289 13685 37323 13719
rect 37323 13685 37332 13719
rect 37280 13676 37332 13685
rect 37464 13719 37516 13728
rect 37464 13685 37473 13719
rect 37473 13685 37507 13719
rect 37507 13685 37516 13719
rect 37464 13676 37516 13685
rect 38292 13719 38344 13728
rect 38292 13685 38301 13719
rect 38301 13685 38335 13719
rect 38335 13685 38344 13719
rect 38292 13676 38344 13685
rect 39120 13744 39172 13796
rect 42800 13719 42852 13728
rect 42800 13685 42809 13719
rect 42809 13685 42843 13719
rect 42843 13685 42852 13719
rect 42800 13676 42852 13685
rect 43536 13719 43588 13728
rect 43536 13685 43545 13719
rect 43545 13685 43579 13719
rect 43579 13685 43588 13719
rect 43536 13676 43588 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 16948 13472 17000 13524
rect 18052 13515 18104 13524
rect 18052 13481 18061 13515
rect 18061 13481 18095 13515
rect 18095 13481 18104 13515
rect 18052 13472 18104 13481
rect 18788 13472 18840 13524
rect 22284 13472 22336 13524
rect 25688 13472 25740 13524
rect 38292 13472 38344 13524
rect 38936 13515 38988 13524
rect 38936 13481 38945 13515
rect 38945 13481 38979 13515
rect 38979 13481 38988 13515
rect 38936 13472 38988 13481
rect 17224 13404 17276 13456
rect 1676 13268 1728 13320
rect 17960 13268 18012 13320
rect 19064 13404 19116 13456
rect 21916 13404 21968 13456
rect 18420 13379 18472 13388
rect 18420 13345 18429 13379
rect 18429 13345 18463 13379
rect 18463 13345 18472 13379
rect 18420 13336 18472 13345
rect 19248 13268 19300 13320
rect 20904 13268 20956 13320
rect 20996 13268 21048 13320
rect 21916 13268 21968 13320
rect 38016 13336 38068 13388
rect 42800 13336 42852 13388
rect 44088 13379 44140 13388
rect 44088 13345 44097 13379
rect 44097 13345 44131 13379
rect 44131 13345 44140 13379
rect 44088 13336 44140 13345
rect 22652 13268 22704 13320
rect 24400 13311 24452 13320
rect 24400 13277 24409 13311
rect 24409 13277 24443 13311
rect 24443 13277 24452 13311
rect 24400 13268 24452 13277
rect 33968 13268 34020 13320
rect 18512 13243 18564 13252
rect 18512 13209 18521 13243
rect 18521 13209 18555 13243
rect 18555 13209 18564 13243
rect 18512 13200 18564 13209
rect 24676 13243 24728 13252
rect 24676 13209 24710 13243
rect 24710 13209 24728 13243
rect 37372 13268 37424 13320
rect 37648 13311 37700 13320
rect 37648 13277 37657 13311
rect 37657 13277 37691 13311
rect 37691 13277 37700 13311
rect 37648 13268 37700 13277
rect 37832 13311 37884 13320
rect 37832 13277 37841 13311
rect 37841 13277 37875 13311
rect 37875 13277 37884 13311
rect 37832 13268 37884 13277
rect 39120 13268 39172 13320
rect 24676 13200 24728 13209
rect 38200 13200 38252 13252
rect 38568 13243 38620 13252
rect 38568 13209 38577 13243
rect 38577 13209 38611 13243
rect 38611 13209 38620 13243
rect 38568 13200 38620 13209
rect 38660 13200 38712 13252
rect 43536 13200 43588 13252
rect 21732 13132 21784 13184
rect 32680 13175 32732 13184
rect 32680 13141 32689 13175
rect 32689 13141 32723 13175
rect 32723 13141 32732 13175
rect 32680 13132 32732 13141
rect 36084 13132 36136 13184
rect 38108 13175 38160 13184
rect 38108 13141 38117 13175
rect 38117 13141 38151 13175
rect 38151 13141 38160 13175
rect 38108 13132 38160 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 18144 12928 18196 12980
rect 19432 12928 19484 12980
rect 18696 12903 18748 12912
rect 18696 12869 18705 12903
rect 18705 12869 18739 12903
rect 18739 12869 18748 12903
rect 18696 12860 18748 12869
rect 1676 12835 1728 12844
rect 1676 12801 1685 12835
rect 1685 12801 1719 12835
rect 1719 12801 1728 12835
rect 1676 12792 1728 12801
rect 9220 12835 9272 12844
rect 9220 12801 9229 12835
rect 9229 12801 9263 12835
rect 9263 12801 9272 12835
rect 9220 12792 9272 12801
rect 12716 12792 12768 12844
rect 18512 12835 18564 12844
rect 18512 12801 18521 12835
rect 18521 12801 18555 12835
rect 18555 12801 18564 12835
rect 18512 12792 18564 12801
rect 20720 12860 20772 12912
rect 20904 12903 20956 12912
rect 20904 12869 20913 12903
rect 20913 12869 20947 12903
rect 20947 12869 20956 12903
rect 20904 12860 20956 12869
rect 21916 12860 21968 12912
rect 19892 12835 19944 12844
rect 19892 12801 19901 12835
rect 19901 12801 19935 12835
rect 19935 12801 19944 12835
rect 19892 12792 19944 12801
rect 21272 12792 21324 12844
rect 22008 12835 22060 12844
rect 22008 12801 22017 12835
rect 22017 12801 22051 12835
rect 22051 12801 22060 12835
rect 22008 12792 22060 12801
rect 24584 12928 24636 12980
rect 25780 12971 25832 12980
rect 25780 12937 25789 12971
rect 25789 12937 25823 12971
rect 25823 12937 25832 12971
rect 25780 12928 25832 12937
rect 27436 12928 27488 12980
rect 36084 12971 36136 12980
rect 36084 12937 36093 12971
rect 36093 12937 36127 12971
rect 36127 12937 36136 12971
rect 36084 12928 36136 12937
rect 37832 12928 37884 12980
rect 27528 12860 27580 12912
rect 31116 12860 31168 12912
rect 31484 12860 31536 12912
rect 38660 12860 38712 12912
rect 23664 12835 23716 12844
rect 1860 12767 1912 12776
rect 1860 12733 1869 12767
rect 1869 12733 1903 12767
rect 1903 12733 1912 12767
rect 1860 12724 1912 12733
rect 2780 12767 2832 12776
rect 2780 12733 2789 12767
rect 2789 12733 2823 12767
rect 2823 12733 2832 12767
rect 2780 12724 2832 12733
rect 18696 12724 18748 12776
rect 21824 12724 21876 12776
rect 23664 12801 23673 12835
rect 23673 12801 23707 12835
rect 23707 12801 23716 12835
rect 23664 12792 23716 12801
rect 23848 12792 23900 12844
rect 27804 12835 27856 12844
rect 27804 12801 27813 12835
rect 27813 12801 27847 12835
rect 27847 12801 27856 12835
rect 27804 12792 27856 12801
rect 27988 12835 28040 12844
rect 27988 12801 27997 12835
rect 27997 12801 28031 12835
rect 28031 12801 28040 12835
rect 27988 12792 28040 12801
rect 29828 12835 29880 12844
rect 29828 12801 29837 12835
rect 29837 12801 29871 12835
rect 29871 12801 29880 12835
rect 29828 12792 29880 12801
rect 32680 12792 32732 12844
rect 33508 12835 33560 12844
rect 33508 12801 33517 12835
rect 33517 12801 33551 12835
rect 33551 12801 33560 12835
rect 33508 12792 33560 12801
rect 36544 12792 36596 12844
rect 38016 12792 38068 12844
rect 38200 12792 38252 12844
rect 43720 12792 43772 12844
rect 24400 12767 24452 12776
rect 24400 12733 24409 12767
rect 24409 12733 24443 12767
rect 24443 12733 24452 12767
rect 24400 12724 24452 12733
rect 34428 12724 34480 12776
rect 35716 12767 35768 12776
rect 35716 12733 35725 12767
rect 35725 12733 35759 12767
rect 35759 12733 35768 12767
rect 35716 12724 35768 12733
rect 38568 12767 38620 12776
rect 38568 12733 38577 12767
rect 38577 12733 38611 12767
rect 38611 12733 38620 12767
rect 38568 12724 38620 12733
rect 41420 12724 41472 12776
rect 23296 12656 23348 12708
rect 9404 12588 9456 12640
rect 21088 12631 21140 12640
rect 21088 12597 21097 12631
rect 21097 12597 21131 12631
rect 21131 12597 21140 12631
rect 21088 12588 21140 12597
rect 22652 12588 22704 12640
rect 24768 12588 24820 12640
rect 28816 12631 28868 12640
rect 28816 12597 28825 12631
rect 28825 12597 28859 12631
rect 28859 12597 28868 12631
rect 28816 12588 28868 12597
rect 30472 12631 30524 12640
rect 30472 12597 30481 12631
rect 30481 12597 30515 12631
rect 30515 12597 30524 12631
rect 30472 12588 30524 12597
rect 32128 12631 32180 12640
rect 32128 12597 32137 12631
rect 32137 12597 32171 12631
rect 32171 12597 32180 12631
rect 32128 12588 32180 12597
rect 35440 12631 35492 12640
rect 35440 12597 35449 12631
rect 35449 12597 35483 12631
rect 35483 12597 35492 12631
rect 35440 12588 35492 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 1860 12384 1912 12436
rect 18420 12427 18472 12436
rect 18420 12393 18429 12427
rect 18429 12393 18463 12427
rect 18463 12393 18472 12427
rect 18420 12384 18472 12393
rect 22008 12384 22060 12436
rect 23848 12427 23900 12436
rect 23848 12393 23857 12427
rect 23857 12393 23891 12427
rect 23891 12393 23900 12427
rect 23848 12384 23900 12393
rect 19892 12291 19944 12300
rect 19892 12257 19901 12291
rect 19901 12257 19935 12291
rect 19935 12257 19944 12291
rect 19892 12248 19944 12257
rect 20812 12248 20864 12300
rect 24584 12291 24636 12300
rect 24584 12257 24593 12291
rect 24593 12257 24627 12291
rect 24627 12257 24636 12291
rect 24584 12248 24636 12257
rect 32128 12248 32180 12300
rect 32312 12291 32364 12300
rect 32312 12257 32321 12291
rect 32321 12257 32355 12291
rect 32355 12257 32364 12291
rect 35348 12291 35400 12300
rect 32312 12248 32364 12257
rect 35348 12257 35357 12291
rect 35357 12257 35391 12291
rect 35391 12257 35400 12291
rect 38936 12316 38988 12368
rect 35348 12248 35400 12257
rect 38292 12248 38344 12300
rect 42708 12291 42760 12300
rect 4896 12180 4948 12232
rect 17868 12180 17920 12232
rect 22652 12223 22704 12232
rect 22652 12189 22670 12223
rect 22670 12189 22704 12223
rect 22652 12180 22704 12189
rect 22836 12180 22888 12232
rect 23664 12223 23716 12232
rect 23664 12189 23673 12223
rect 23673 12189 23707 12223
rect 23707 12189 23716 12223
rect 23664 12180 23716 12189
rect 18328 12112 18380 12164
rect 21640 12112 21692 12164
rect 27344 12180 27396 12232
rect 25688 12155 25740 12164
rect 25688 12121 25722 12155
rect 25722 12121 25740 12155
rect 25688 12112 25740 12121
rect 18604 12044 18656 12096
rect 24768 12044 24820 12096
rect 25872 12044 25924 12096
rect 27988 12180 28040 12232
rect 28448 12180 28500 12232
rect 31116 12180 31168 12232
rect 33324 12223 33376 12232
rect 33324 12189 33333 12223
rect 33333 12189 33367 12223
rect 33367 12189 33376 12223
rect 33324 12180 33376 12189
rect 30472 12112 30524 12164
rect 31024 12087 31076 12096
rect 31024 12053 31033 12087
rect 31033 12053 31067 12087
rect 31067 12053 31076 12087
rect 31024 12044 31076 12053
rect 31208 12044 31260 12096
rect 32128 12087 32180 12096
rect 32128 12053 32137 12087
rect 32137 12053 32171 12087
rect 32171 12053 32180 12087
rect 32128 12044 32180 12053
rect 33140 12087 33192 12096
rect 33140 12053 33149 12087
rect 33149 12053 33183 12087
rect 33183 12053 33192 12087
rect 33140 12044 33192 12053
rect 33784 12087 33836 12096
rect 33784 12053 33793 12087
rect 33793 12053 33827 12087
rect 33827 12053 33836 12087
rect 33784 12044 33836 12053
rect 35440 12180 35492 12232
rect 37648 12180 37700 12232
rect 42708 12257 42717 12291
rect 42717 12257 42751 12291
rect 42751 12257 42760 12291
rect 42708 12248 42760 12257
rect 44180 12223 44232 12232
rect 44180 12189 44189 12223
rect 44189 12189 44223 12223
rect 44223 12189 44232 12223
rect 44180 12180 44232 12189
rect 38844 12112 38896 12164
rect 43444 12112 43496 12164
rect 35532 12044 35584 12096
rect 35900 12087 35952 12096
rect 35900 12053 35909 12087
rect 35909 12053 35943 12087
rect 35943 12053 35952 12087
rect 36268 12087 36320 12096
rect 35900 12044 35952 12053
rect 36268 12053 36277 12087
rect 36277 12053 36311 12087
rect 36311 12053 36320 12087
rect 36268 12044 36320 12053
rect 38292 12044 38344 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 24676 11840 24728 11892
rect 25688 11883 25740 11892
rect 25688 11849 25697 11883
rect 25697 11849 25731 11883
rect 25731 11849 25740 11883
rect 25688 11840 25740 11849
rect 29828 11883 29880 11892
rect 29828 11849 29837 11883
rect 29837 11849 29871 11883
rect 29871 11849 29880 11883
rect 29828 11840 29880 11849
rect 30748 11840 30800 11892
rect 31208 11883 31260 11892
rect 31208 11849 31217 11883
rect 31217 11849 31251 11883
rect 31251 11849 31260 11883
rect 31208 11840 31260 11849
rect 32128 11883 32180 11892
rect 32128 11849 32137 11883
rect 32137 11849 32171 11883
rect 32171 11849 32180 11883
rect 32128 11840 32180 11849
rect 33324 11840 33376 11892
rect 35532 11883 35584 11892
rect 35532 11849 35541 11883
rect 35541 11849 35575 11883
rect 35575 11849 35584 11883
rect 35532 11840 35584 11849
rect 35716 11883 35768 11892
rect 35716 11849 35725 11883
rect 35725 11849 35759 11883
rect 35759 11849 35768 11883
rect 35716 11840 35768 11849
rect 36544 11840 36596 11892
rect 43444 11883 43496 11892
rect 43444 11849 43453 11883
rect 43453 11849 43487 11883
rect 43487 11849 43496 11883
rect 43444 11840 43496 11849
rect 20260 11815 20312 11824
rect 20260 11781 20269 11815
rect 20269 11781 20303 11815
rect 20303 11781 20312 11815
rect 20260 11772 20312 11781
rect 28816 11772 28868 11824
rect 33140 11772 33192 11824
rect 35900 11772 35952 11824
rect 36636 11772 36688 11824
rect 37096 11772 37148 11824
rect 37556 11815 37608 11824
rect 37556 11781 37565 11815
rect 37565 11781 37599 11815
rect 37599 11781 37608 11815
rect 37556 11772 37608 11781
rect 38108 11772 38160 11824
rect 17500 11704 17552 11756
rect 20812 11704 20864 11756
rect 23756 11747 23808 11756
rect 23756 11713 23765 11747
rect 23765 11713 23799 11747
rect 23799 11713 23808 11747
rect 23756 11704 23808 11713
rect 24400 11747 24452 11756
rect 24400 11713 24409 11747
rect 24409 11713 24443 11747
rect 24443 11713 24452 11747
rect 24400 11704 24452 11713
rect 25044 11747 25096 11756
rect 25044 11713 25053 11747
rect 25053 11713 25087 11747
rect 25087 11713 25096 11747
rect 25044 11704 25096 11713
rect 25872 11747 25924 11756
rect 25872 11713 25881 11747
rect 25881 11713 25915 11747
rect 25915 11713 25924 11747
rect 25872 11704 25924 11713
rect 28448 11747 28500 11756
rect 28448 11713 28457 11747
rect 28457 11713 28491 11747
rect 28491 11713 28500 11747
rect 28448 11704 28500 11713
rect 31024 11704 31076 11756
rect 33508 11747 33560 11756
rect 16672 11636 16724 11688
rect 19064 11679 19116 11688
rect 18512 11568 18564 11620
rect 19064 11645 19073 11679
rect 19073 11645 19107 11679
rect 19107 11645 19116 11679
rect 19064 11636 19116 11645
rect 31300 11679 31352 11688
rect 31300 11645 31309 11679
rect 31309 11645 31343 11679
rect 31343 11645 31352 11679
rect 31300 11636 31352 11645
rect 33508 11713 33517 11747
rect 33517 11713 33551 11747
rect 33551 11713 33560 11747
rect 33508 11704 33560 11713
rect 34704 11747 34756 11756
rect 34704 11713 34713 11747
rect 34713 11713 34747 11747
rect 34747 11713 34756 11747
rect 34704 11704 34756 11713
rect 37188 11704 37240 11756
rect 38200 11747 38252 11756
rect 38200 11713 38209 11747
rect 38209 11713 38243 11747
rect 38243 11713 38252 11747
rect 38200 11704 38252 11713
rect 38292 11747 38344 11756
rect 38292 11713 38301 11747
rect 38301 11713 38335 11747
rect 38335 11713 38344 11747
rect 38292 11704 38344 11713
rect 42892 11704 42944 11756
rect 44180 11747 44232 11756
rect 44180 11713 44189 11747
rect 44189 11713 44223 11747
rect 44223 11713 44232 11747
rect 44180 11704 44232 11713
rect 36176 11679 36228 11688
rect 36176 11645 36185 11679
rect 36185 11645 36219 11679
rect 36219 11645 36228 11679
rect 36176 11636 36228 11645
rect 37372 11636 37424 11688
rect 35716 11568 35768 11620
rect 36268 11568 36320 11620
rect 17684 11500 17736 11552
rect 19616 11500 19668 11552
rect 20720 11500 20772 11552
rect 24216 11500 24268 11552
rect 25412 11500 25464 11552
rect 37832 11500 37884 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 18512 11339 18564 11348
rect 18512 11305 18521 11339
rect 18521 11305 18555 11339
rect 18555 11305 18564 11339
rect 18512 11296 18564 11305
rect 18696 11339 18748 11348
rect 18696 11305 18705 11339
rect 18705 11305 18739 11339
rect 18739 11305 18748 11339
rect 18696 11296 18748 11305
rect 21640 11339 21692 11348
rect 21640 11305 21649 11339
rect 21649 11305 21683 11339
rect 21683 11305 21692 11339
rect 21640 11296 21692 11305
rect 24400 11296 24452 11348
rect 25044 11296 25096 11348
rect 26792 11296 26844 11348
rect 27344 11339 27396 11348
rect 27344 11305 27353 11339
rect 27353 11305 27387 11339
rect 27387 11305 27396 11339
rect 27344 11296 27396 11305
rect 31300 11296 31352 11348
rect 34704 11296 34756 11348
rect 17132 11160 17184 11212
rect 18236 11228 18288 11280
rect 19432 11228 19484 11280
rect 17684 11160 17736 11212
rect 19340 11160 19392 11212
rect 3240 11092 3292 11144
rect 17776 11135 17828 11144
rect 17776 11101 17785 11135
rect 17785 11101 17819 11135
rect 17819 11101 17828 11135
rect 17776 11092 17828 11101
rect 17868 11135 17920 11144
rect 17868 11101 17877 11135
rect 17877 11101 17911 11135
rect 17911 11101 17920 11135
rect 17868 11092 17920 11101
rect 19064 11092 19116 11144
rect 19616 11135 19668 11144
rect 19616 11101 19625 11135
rect 19625 11101 19659 11135
rect 19659 11101 19668 11135
rect 19616 11092 19668 11101
rect 23480 11135 23532 11144
rect 23480 11101 23489 11135
rect 23489 11101 23523 11135
rect 23523 11101 23532 11135
rect 23480 11092 23532 11101
rect 24216 11092 24268 11144
rect 18328 11067 18380 11076
rect 18328 11033 18337 11067
rect 18337 11033 18371 11067
rect 18371 11033 18380 11067
rect 18328 11024 18380 11033
rect 17592 10999 17644 11008
rect 17592 10965 17601 10999
rect 17601 10965 17635 10999
rect 17635 10965 17644 10999
rect 17592 10956 17644 10965
rect 17776 10956 17828 11008
rect 20812 11024 20864 11076
rect 24768 11092 24820 11144
rect 25412 11092 25464 11144
rect 27988 11160 28040 11212
rect 30196 11135 30248 11144
rect 30196 11101 30205 11135
rect 30205 11101 30239 11135
rect 30239 11101 30248 11135
rect 30196 11092 30248 11101
rect 33508 11092 33560 11144
rect 35348 11092 35400 11144
rect 36176 11160 36228 11212
rect 43720 11203 43772 11212
rect 43720 11169 43729 11203
rect 43729 11169 43763 11203
rect 43763 11169 43772 11203
rect 43720 11160 43772 11169
rect 37372 11092 37424 11144
rect 44180 11135 44232 11144
rect 44180 11101 44189 11135
rect 44189 11101 44223 11135
rect 44223 11101 44232 11135
rect 44180 11092 44232 11101
rect 27620 11067 27672 11076
rect 27620 11033 27629 11067
rect 27629 11033 27663 11067
rect 27663 11033 27672 11067
rect 27620 11024 27672 11033
rect 27804 11024 27856 11076
rect 32312 11067 32364 11076
rect 32312 11033 32321 11067
rect 32321 11033 32355 11067
rect 32355 11033 32364 11067
rect 32312 11024 32364 11033
rect 33784 11024 33836 11076
rect 36636 11024 36688 11076
rect 37648 11024 37700 11076
rect 43996 11067 44048 11076
rect 43996 11033 44005 11067
rect 44005 11033 44039 11067
rect 44039 11033 44048 11067
rect 43996 11024 44048 11033
rect 28172 10956 28224 11008
rect 30840 10999 30892 11008
rect 30840 10965 30849 10999
rect 30849 10965 30883 10999
rect 30883 10965 30892 10999
rect 30840 10956 30892 10965
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 17868 10752 17920 10804
rect 20260 10752 20312 10804
rect 23664 10795 23716 10804
rect 23664 10761 23673 10795
rect 23673 10761 23707 10795
rect 23707 10761 23716 10795
rect 23664 10752 23716 10761
rect 27344 10752 27396 10804
rect 30196 10795 30248 10804
rect 17592 10684 17644 10736
rect 19064 10684 19116 10736
rect 30196 10761 30205 10795
rect 30205 10761 30239 10795
rect 30239 10761 30248 10795
rect 30196 10752 30248 10761
rect 43996 10752 44048 10804
rect 2596 10659 2648 10668
rect 2596 10625 2605 10659
rect 2605 10625 2639 10659
rect 2639 10625 2648 10659
rect 2596 10616 2648 10625
rect 4988 10616 5040 10668
rect 17776 10659 17828 10668
rect 17776 10625 17785 10659
rect 17785 10625 17819 10659
rect 17819 10625 17828 10659
rect 17776 10616 17828 10625
rect 18420 10616 18472 10668
rect 18696 10591 18748 10600
rect 18696 10557 18705 10591
rect 18705 10557 18739 10591
rect 18739 10557 18748 10591
rect 18696 10548 18748 10557
rect 17500 10523 17552 10532
rect 17500 10489 17509 10523
rect 17509 10489 17543 10523
rect 17543 10489 17552 10523
rect 17500 10480 17552 10489
rect 1860 10412 1912 10464
rect 2136 10412 2188 10464
rect 23112 10616 23164 10668
rect 24216 10659 24268 10668
rect 24216 10625 24225 10659
rect 24225 10625 24259 10659
rect 24259 10625 24268 10659
rect 24216 10616 24268 10625
rect 24952 10616 25004 10668
rect 28172 10659 28224 10668
rect 28172 10625 28181 10659
rect 28181 10625 28215 10659
rect 28215 10625 28224 10659
rect 28172 10616 28224 10625
rect 28448 10616 28500 10668
rect 43352 10659 43404 10668
rect 43352 10625 43361 10659
rect 43361 10625 43395 10659
rect 43395 10625 43404 10659
rect 43352 10616 43404 10625
rect 44180 10659 44232 10668
rect 44180 10625 44189 10659
rect 44189 10625 44223 10659
rect 44223 10625 44232 10659
rect 44180 10616 44232 10625
rect 20812 10591 20864 10600
rect 20812 10557 20821 10591
rect 20821 10557 20855 10591
rect 20855 10557 20864 10591
rect 20812 10548 20864 10557
rect 21640 10548 21692 10600
rect 24860 10548 24912 10600
rect 21916 10480 21968 10532
rect 20812 10412 20864 10464
rect 25412 10412 25464 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 1400 10115 1452 10124
rect 1400 10081 1409 10115
rect 1409 10081 1443 10115
rect 1443 10081 1452 10115
rect 1400 10072 1452 10081
rect 3240 10115 3292 10124
rect 3240 10081 3249 10115
rect 3249 10081 3283 10115
rect 3283 10081 3292 10115
rect 3240 10072 3292 10081
rect 17684 10208 17736 10260
rect 18696 10251 18748 10260
rect 18696 10217 18705 10251
rect 18705 10217 18739 10251
rect 18739 10217 18748 10251
rect 18696 10208 18748 10217
rect 20720 10208 20772 10260
rect 21916 10183 21968 10192
rect 21916 10149 21925 10183
rect 21925 10149 21959 10183
rect 21959 10149 21968 10183
rect 23112 10251 23164 10260
rect 23112 10217 23121 10251
rect 23121 10217 23155 10251
rect 23155 10217 23164 10251
rect 23112 10208 23164 10217
rect 32312 10208 32364 10260
rect 21916 10140 21968 10149
rect 23664 10140 23716 10192
rect 19432 10072 19484 10124
rect 24216 10072 24268 10124
rect 28448 10072 28500 10124
rect 3976 10047 4028 10056
rect 3976 10013 3985 10047
rect 3985 10013 4019 10047
rect 4019 10013 4028 10047
rect 3976 10004 4028 10013
rect 17684 9936 17736 9988
rect 20352 10004 20404 10056
rect 22928 10004 22980 10056
rect 20536 9979 20588 9988
rect 20536 9945 20545 9979
rect 20545 9945 20579 9979
rect 20579 9945 20588 9979
rect 20536 9936 20588 9945
rect 24860 10004 24912 10056
rect 30840 10004 30892 10056
rect 25596 9936 25648 9988
rect 19432 9868 19484 9920
rect 20996 9911 21048 9920
rect 20996 9877 21005 9911
rect 21005 9877 21039 9911
rect 21039 9877 21048 9911
rect 20996 9868 21048 9877
rect 22284 9911 22336 9920
rect 22284 9877 22293 9911
rect 22293 9877 22327 9911
rect 22327 9877 22336 9911
rect 22284 9868 22336 9877
rect 23112 9911 23164 9920
rect 23112 9877 23139 9911
rect 23139 9877 23164 9911
rect 23112 9868 23164 9877
rect 24676 9868 24728 9920
rect 27620 9936 27672 9988
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 17684 9707 17736 9716
rect 17684 9673 17693 9707
rect 17693 9673 17727 9707
rect 17727 9673 17736 9707
rect 17684 9664 17736 9673
rect 24952 9707 25004 9716
rect 24952 9673 24961 9707
rect 24961 9673 24995 9707
rect 24995 9673 25004 9707
rect 24952 9664 25004 9673
rect 25596 9707 25648 9716
rect 25596 9673 25605 9707
rect 25605 9673 25639 9707
rect 25639 9673 25648 9707
rect 25596 9664 25648 9673
rect 3976 9596 4028 9648
rect 17776 9571 17828 9580
rect 1952 9503 2004 9512
rect 1952 9469 1961 9503
rect 1961 9469 1995 9503
rect 1995 9469 2004 9503
rect 1952 9460 2004 9469
rect 2504 9460 2556 9512
rect 2780 9503 2832 9512
rect 2780 9469 2789 9503
rect 2789 9469 2823 9503
rect 2823 9469 2832 9503
rect 2780 9460 2832 9469
rect 17776 9537 17785 9571
rect 17785 9537 17819 9571
rect 17819 9537 17828 9571
rect 17776 9528 17828 9537
rect 18420 9571 18472 9580
rect 18420 9537 18429 9571
rect 18429 9537 18463 9571
rect 18463 9537 18472 9571
rect 18420 9528 18472 9537
rect 18696 9528 18748 9580
rect 19340 9571 19392 9580
rect 19340 9537 19349 9571
rect 19349 9537 19383 9571
rect 19383 9537 19392 9571
rect 19340 9528 19392 9537
rect 19616 9571 19668 9580
rect 19616 9537 19650 9571
rect 19650 9537 19668 9571
rect 19616 9528 19668 9537
rect 22376 9571 22428 9580
rect 22376 9537 22385 9571
rect 22385 9537 22419 9571
rect 22419 9537 22428 9571
rect 22376 9528 22428 9537
rect 23112 9528 23164 9580
rect 23664 9571 23716 9580
rect 23664 9537 23673 9571
rect 23673 9537 23707 9571
rect 23707 9537 23716 9571
rect 23664 9528 23716 9537
rect 24676 9528 24728 9580
rect 25412 9571 25464 9580
rect 25412 9537 25421 9571
rect 25421 9537 25455 9571
rect 25455 9537 25464 9571
rect 25412 9528 25464 9537
rect 18236 9503 18288 9512
rect 18236 9469 18245 9503
rect 18245 9469 18279 9503
rect 18279 9469 18288 9503
rect 18236 9460 18288 9469
rect 20536 9460 20588 9512
rect 23480 9460 23532 9512
rect 20352 9392 20404 9444
rect 23020 9392 23072 9444
rect 23848 9367 23900 9376
rect 23848 9333 23857 9367
rect 23857 9333 23891 9367
rect 23891 9333 23900 9367
rect 23848 9324 23900 9333
rect 42524 9324 42576 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 1952 9163 2004 9172
rect 1952 9129 1961 9163
rect 1961 9129 1995 9163
rect 1995 9129 2004 9163
rect 1952 9120 2004 9129
rect 2504 9163 2556 9172
rect 2504 9129 2513 9163
rect 2513 9129 2547 9163
rect 2547 9129 2556 9163
rect 2504 9120 2556 9129
rect 19616 9163 19668 9172
rect 19616 9129 19625 9163
rect 19625 9129 19659 9163
rect 19659 9129 19668 9163
rect 19616 9120 19668 9129
rect 22284 9120 22336 9172
rect 42524 9027 42576 9036
rect 42524 8993 42533 9027
rect 42533 8993 42567 9027
rect 42567 8993 42576 9027
rect 42524 8984 42576 8993
rect 2596 8959 2648 8968
rect 2596 8925 2605 8959
rect 2605 8925 2639 8959
rect 2639 8925 2648 8959
rect 2596 8916 2648 8925
rect 19432 8916 19484 8968
rect 20536 8916 20588 8968
rect 22836 8916 22888 8968
rect 22928 8959 22980 8968
rect 22928 8925 22937 8959
rect 22937 8925 22971 8959
rect 22971 8925 22980 8959
rect 22928 8916 22980 8925
rect 23480 8916 23532 8968
rect 42340 8959 42392 8968
rect 42340 8925 42349 8959
rect 42349 8925 42383 8959
rect 42383 8925 42392 8959
rect 42340 8916 42392 8925
rect 20352 8848 20404 8900
rect 21180 8891 21232 8900
rect 21180 8857 21214 8891
rect 21214 8857 21232 8891
rect 21180 8848 21232 8857
rect 23020 8848 23072 8900
rect 45100 8848 45152 8900
rect 22376 8780 22428 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 21180 8619 21232 8628
rect 21180 8585 21189 8619
rect 21189 8585 21223 8619
rect 21223 8585 21232 8619
rect 21180 8576 21232 8585
rect 22928 8576 22980 8628
rect 2136 8551 2188 8560
rect 2136 8517 2145 8551
rect 2145 8517 2179 8551
rect 2179 8517 2188 8551
rect 2136 8508 2188 8517
rect 23848 8551 23900 8560
rect 23848 8517 23866 8551
rect 23866 8517 23900 8551
rect 23848 8508 23900 8517
rect 1860 8440 1912 8492
rect 20996 8483 21048 8492
rect 20996 8449 21005 8483
rect 21005 8449 21039 8483
rect 21039 8449 21048 8483
rect 20996 8440 21048 8449
rect 24768 8440 24820 8492
rect 42340 8440 42392 8492
rect 2872 8415 2924 8424
rect 2872 8381 2881 8415
rect 2881 8381 2915 8415
rect 2915 8381 2924 8415
rect 2872 8372 2924 8381
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 44180 7871 44232 7880
rect 44180 7837 44189 7871
rect 44189 7837 44223 7871
rect 44223 7837 44232 7871
rect 44180 7828 44232 7837
rect 26332 7692 26384 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 3424 7395 3476 7404
rect 3424 7361 3433 7395
rect 3433 7361 3467 7395
rect 3467 7361 3476 7395
rect 3424 7352 3476 7361
rect 43628 7352 43680 7404
rect 3516 7191 3568 7200
rect 3516 7157 3525 7191
rect 3525 7157 3559 7191
rect 3559 7157 3568 7191
rect 3516 7148 3568 7157
rect 4068 7191 4120 7200
rect 4068 7157 4077 7191
rect 4077 7157 4111 7191
rect 4111 7157 4120 7191
rect 4068 7148 4120 7157
rect 43996 7148 44048 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 4068 6808 4120 6860
rect 4712 6851 4764 6860
rect 4712 6817 4721 6851
rect 4721 6817 4755 6851
rect 4755 6817 4764 6851
rect 4712 6808 4764 6817
rect 1676 6740 1728 6792
rect 3516 6672 3568 6724
rect 4068 6672 4120 6724
rect 14740 6808 14792 6860
rect 42708 6851 42760 6860
rect 42708 6817 42717 6851
rect 42717 6817 42751 6851
rect 42751 6817 42760 6851
rect 42708 6808 42760 6817
rect 43996 6851 44048 6860
rect 43996 6817 44005 6851
rect 44005 6817 44039 6851
rect 44039 6817 44048 6851
rect 43996 6808 44048 6817
rect 44180 6783 44232 6792
rect 44180 6749 44189 6783
rect 44189 6749 44223 6783
rect 44223 6749 44232 6783
rect 44180 6740 44232 6749
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 1676 6307 1728 6316
rect 1676 6273 1685 6307
rect 1685 6273 1719 6307
rect 1719 6273 1728 6307
rect 1676 6264 1728 6273
rect 44180 6264 44232 6316
rect 2136 6196 2188 6248
rect 2780 6239 2832 6248
rect 2780 6205 2789 6239
rect 2789 6205 2823 6239
rect 2823 6205 2832 6239
rect 2780 6196 2832 6205
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 2136 5899 2188 5908
rect 2136 5865 2145 5899
rect 2145 5865 2179 5899
rect 2179 5865 2188 5899
rect 2136 5856 2188 5865
rect 1584 5695 1636 5704
rect 1584 5661 1593 5695
rect 1593 5661 1627 5695
rect 1627 5661 1636 5695
rect 1584 5652 1636 5661
rect 2044 5652 2096 5704
rect 5908 5788 5960 5840
rect 6276 5720 6328 5772
rect 42708 5763 42760 5772
rect 42708 5729 42717 5763
rect 42717 5729 42751 5763
rect 42751 5729 42760 5763
rect 42708 5720 42760 5729
rect 3792 5695 3844 5704
rect 3792 5661 3801 5695
rect 3801 5661 3835 5695
rect 3835 5661 3844 5695
rect 3792 5652 3844 5661
rect 4160 5652 4212 5704
rect 44180 5695 44232 5704
rect 44180 5661 44189 5695
rect 44189 5661 44223 5695
rect 44223 5661 44232 5695
rect 44180 5652 44232 5661
rect 43996 5627 44048 5636
rect 43996 5593 44005 5627
rect 44005 5593 44039 5627
rect 44039 5593 44048 5627
rect 43996 5584 44048 5593
rect 2872 5559 2924 5568
rect 2872 5525 2881 5559
rect 2881 5525 2915 5559
rect 2915 5525 2924 5559
rect 2872 5516 2924 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 2872 5244 2924 5296
rect 1584 5176 1636 5228
rect 4620 5176 4672 5228
rect 42800 5219 42852 5228
rect 42800 5185 42809 5219
rect 42809 5185 42843 5219
rect 42843 5185 42852 5219
rect 42800 5176 42852 5185
rect 2780 5151 2832 5160
rect 2780 5117 2789 5151
rect 2789 5117 2823 5151
rect 2823 5117 2832 5151
rect 2780 5108 2832 5117
rect 4620 4972 4672 5024
rect 4896 5015 4948 5024
rect 4896 4981 4905 5015
rect 4905 4981 4939 5015
rect 4939 4981 4948 5015
rect 4896 4972 4948 4981
rect 42524 4972 42576 5024
rect 43628 5015 43680 5024
rect 43628 4981 43637 5015
rect 43637 4981 43671 5015
rect 43671 4981 43680 5015
rect 43628 4972 43680 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 4804 4768 4856 4820
rect 2964 4632 3016 4684
rect 3148 4564 3200 4616
rect 11796 4700 11848 4752
rect 4068 4675 4120 4684
rect 4068 4641 4077 4675
rect 4077 4641 4111 4675
rect 4111 4641 4120 4675
rect 4068 4632 4120 4641
rect 4620 4632 4672 4684
rect 4804 4675 4856 4684
rect 4804 4641 4813 4675
rect 4813 4641 4847 4675
rect 4847 4641 4856 4675
rect 4804 4632 4856 4641
rect 38016 4675 38068 4684
rect 38016 4641 38025 4675
rect 38025 4641 38059 4675
rect 38059 4641 38068 4675
rect 38016 4632 38068 4641
rect 43628 4700 43680 4752
rect 42524 4675 42576 4684
rect 42524 4641 42533 4675
rect 42533 4641 42567 4675
rect 42567 4641 42576 4675
rect 42524 4632 42576 4641
rect 44088 4675 44140 4684
rect 44088 4641 44097 4675
rect 44097 4641 44131 4675
rect 44131 4641 44140 4675
rect 44088 4632 44140 4641
rect 6276 4564 6328 4616
rect 37372 4607 37424 4616
rect 37372 4573 37381 4607
rect 37381 4573 37415 4607
rect 37415 4573 37424 4607
rect 37372 4564 37424 4573
rect 37556 4539 37608 4548
rect 37556 4505 37565 4539
rect 37565 4505 37599 4539
rect 37599 4505 37608 4539
rect 37556 4496 37608 4505
rect 4160 4428 4212 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 2044 4131 2096 4140
rect 2044 4097 2053 4131
rect 2053 4097 2087 4131
rect 2087 4097 2096 4131
rect 2044 4088 2096 4097
rect 4896 4088 4948 4140
rect 11796 4131 11848 4140
rect 2780 4063 2832 4072
rect 2780 4029 2789 4063
rect 2789 4029 2823 4063
rect 2823 4029 2832 4063
rect 4160 4063 4212 4072
rect 2780 4020 2832 4029
rect 4160 4029 4169 4063
rect 4169 4029 4203 4063
rect 4203 4029 4212 4063
rect 4160 4020 4212 4029
rect 11796 4097 11805 4131
rect 11805 4097 11839 4131
rect 11839 4097 11848 4131
rect 11796 4088 11848 4097
rect 18696 4088 18748 4140
rect 36544 4131 36596 4140
rect 36544 4097 36553 4131
rect 36553 4097 36587 4131
rect 36587 4097 36596 4131
rect 36544 4088 36596 4097
rect 37372 4088 37424 4140
rect 42984 4088 43036 4140
rect 43352 4131 43404 4140
rect 43352 4097 43361 4131
rect 43361 4097 43395 4131
rect 43395 4097 43404 4131
rect 43352 4088 43404 4097
rect 2320 3952 2372 4004
rect 6184 3952 6236 4004
rect 9496 3952 9548 4004
rect 38200 4020 38252 4072
rect 38844 4063 38896 4072
rect 38844 4029 38853 4063
rect 38853 4029 38887 4063
rect 38887 4029 38896 4063
rect 38844 4020 38896 4029
rect 36452 3952 36504 4004
rect 37464 3952 37516 4004
rect 38292 3952 38344 4004
rect 41328 4020 41380 4072
rect 1584 3884 1636 3936
rect 3884 3884 3936 3936
rect 4712 3884 4764 3936
rect 5540 3884 5592 3936
rect 6368 3927 6420 3936
rect 6368 3893 6377 3927
rect 6377 3893 6411 3927
rect 6411 3893 6420 3927
rect 6368 3884 6420 3893
rect 7288 3884 7340 3936
rect 9220 3884 9272 3936
rect 11888 3927 11940 3936
rect 11888 3893 11897 3927
rect 11897 3893 11931 3927
rect 11931 3893 11940 3927
rect 11888 3884 11940 3893
rect 12440 3927 12492 3936
rect 12440 3893 12449 3927
rect 12449 3893 12483 3927
rect 12483 3893 12492 3927
rect 12440 3884 12492 3893
rect 15476 3884 15528 3936
rect 20812 3884 20864 3936
rect 24216 3927 24268 3936
rect 24216 3893 24225 3927
rect 24225 3893 24259 3927
rect 24259 3893 24268 3927
rect 24216 3884 24268 3893
rect 37280 3927 37332 3936
rect 37280 3893 37289 3927
rect 37289 3893 37323 3927
rect 37323 3893 37332 3927
rect 37280 3884 37332 3893
rect 41880 3884 41932 3936
rect 42432 3927 42484 3936
rect 42432 3893 42441 3927
rect 42441 3893 42475 3927
rect 42475 3893 42484 3927
rect 42432 3884 42484 3893
rect 43444 3927 43496 3936
rect 43444 3893 43453 3927
rect 43453 3893 43487 3927
rect 43487 3893 43496 3927
rect 43444 3884 43496 3893
rect 43536 3884 43588 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 2964 3544 3016 3596
rect 6368 3612 6420 3664
rect 5540 3587 5592 3596
rect 5540 3553 5549 3587
rect 5549 3553 5583 3587
rect 5583 3553 5592 3587
rect 5540 3544 5592 3553
rect 5816 3587 5868 3596
rect 5816 3553 5825 3587
rect 5825 3553 5859 3587
rect 5859 3553 5868 3587
rect 5816 3544 5868 3553
rect 1400 3519 1452 3528
rect 1400 3485 1409 3519
rect 1409 3485 1443 3519
rect 1443 3485 1452 3519
rect 1400 3476 1452 3485
rect 4528 3519 4580 3528
rect 4528 3485 4537 3519
rect 4537 3485 4571 3519
rect 4571 3485 4580 3519
rect 4528 3476 4580 3485
rect 12808 3680 12860 3732
rect 13268 3680 13320 3732
rect 38292 3723 38344 3732
rect 38292 3689 38301 3723
rect 38301 3689 38335 3723
rect 38335 3689 38344 3723
rect 38292 3680 38344 3689
rect 38844 3723 38896 3732
rect 38844 3689 38853 3723
rect 38853 3689 38887 3723
rect 38887 3689 38896 3723
rect 38844 3680 38896 3689
rect 9496 3612 9548 3664
rect 9220 3587 9272 3596
rect 9220 3553 9229 3587
rect 9229 3553 9263 3587
rect 9263 3553 9272 3587
rect 9404 3587 9456 3596
rect 9220 3544 9272 3553
rect 9404 3553 9413 3587
rect 9413 3553 9447 3587
rect 9447 3553 9456 3587
rect 9404 3544 9456 3553
rect 9680 3587 9732 3596
rect 9680 3553 9689 3587
rect 9689 3553 9723 3587
rect 9723 3553 9732 3587
rect 9680 3544 9732 3553
rect 12992 3544 13044 3596
rect 15476 3587 15528 3596
rect 15476 3553 15485 3587
rect 15485 3553 15519 3587
rect 15519 3553 15528 3587
rect 15476 3544 15528 3553
rect 16120 3587 16172 3596
rect 16120 3553 16129 3587
rect 16129 3553 16163 3587
rect 16163 3553 16172 3587
rect 16120 3544 16172 3553
rect 13360 3476 13412 3528
rect 16856 3476 16908 3528
rect 18788 3476 18840 3528
rect 36544 3612 36596 3664
rect 20812 3587 20864 3596
rect 20812 3553 20821 3587
rect 20821 3553 20855 3587
rect 20855 3553 20864 3587
rect 20812 3544 20864 3553
rect 21272 3587 21324 3596
rect 21272 3553 21281 3587
rect 21281 3553 21315 3587
rect 21315 3553 21324 3587
rect 21272 3544 21324 3553
rect 22100 3476 22152 3528
rect 24768 3519 24820 3528
rect 2228 3408 2280 3460
rect 3700 3408 3752 3460
rect 13084 3408 13136 3460
rect 15752 3408 15804 3460
rect 24768 3485 24777 3519
rect 24777 3485 24811 3519
rect 24811 3485 24820 3519
rect 24768 3476 24820 3485
rect 4620 3340 4672 3392
rect 7472 3340 7524 3392
rect 13176 3340 13228 3392
rect 13268 3340 13320 3392
rect 24400 3408 24452 3460
rect 29184 3476 29236 3528
rect 35532 3544 35584 3596
rect 36084 3587 36136 3596
rect 36084 3553 36093 3587
rect 36093 3553 36127 3587
rect 36127 3553 36136 3587
rect 36084 3544 36136 3553
rect 36452 3544 36504 3596
rect 42800 3680 42852 3732
rect 43996 3680 44048 3732
rect 42432 3612 42484 3664
rect 35624 3519 35676 3528
rect 35624 3485 35633 3519
rect 35633 3485 35667 3519
rect 35667 3485 35676 3519
rect 35624 3476 35676 3485
rect 38200 3519 38252 3528
rect 38200 3485 38209 3519
rect 38209 3485 38243 3519
rect 38243 3485 38252 3519
rect 38200 3476 38252 3485
rect 40040 3519 40092 3528
rect 40040 3485 40049 3519
rect 40049 3485 40083 3519
rect 40083 3485 40092 3519
rect 40040 3476 40092 3485
rect 41880 3587 41932 3596
rect 41880 3553 41889 3587
rect 41889 3553 41923 3587
rect 41923 3553 41932 3587
rect 41880 3544 41932 3553
rect 42524 3587 42576 3596
rect 42524 3553 42533 3587
rect 42533 3553 42567 3587
rect 42567 3553 42576 3587
rect 42524 3544 42576 3553
rect 43904 3476 43956 3528
rect 37372 3408 37424 3460
rect 39948 3408 40000 3460
rect 18972 3340 19024 3392
rect 23756 3383 23808 3392
rect 23756 3349 23765 3383
rect 23765 3349 23799 3383
rect 23799 3349 23808 3383
rect 23756 3340 23808 3349
rect 24584 3340 24636 3392
rect 29368 3340 29420 3392
rect 36544 3340 36596 3392
rect 42892 3408 42944 3460
rect 40224 3340 40276 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 2228 3179 2280 3188
rect 2228 3145 2237 3179
rect 2237 3145 2271 3179
rect 2271 3145 2280 3179
rect 2228 3136 2280 3145
rect 4528 3136 4580 3188
rect 2320 3043 2372 3052
rect 2320 3009 2329 3043
rect 2329 3009 2363 3043
rect 2363 3009 2372 3043
rect 2320 3000 2372 3009
rect 3148 3000 3200 3052
rect 9588 3136 9640 3188
rect 15752 3179 15804 3188
rect 7472 3111 7524 3120
rect 7472 3077 7481 3111
rect 7481 3077 7515 3111
rect 7515 3077 7524 3111
rect 7472 3068 7524 3077
rect 13176 3111 13228 3120
rect 7288 3043 7340 3052
rect 7288 3009 7297 3043
rect 7297 3009 7331 3043
rect 7331 3009 7340 3043
rect 7288 3000 7340 3009
rect 3700 2932 3752 2984
rect 3976 2975 4028 2984
rect 3976 2941 3985 2975
rect 3985 2941 4019 2975
rect 4019 2941 4028 2975
rect 3976 2932 4028 2941
rect 7104 2932 7156 2984
rect 664 2864 716 2916
rect 4712 2864 4764 2916
rect 5172 2864 5224 2916
rect 13176 3077 13185 3111
rect 13185 3077 13219 3111
rect 13219 3077 13228 3111
rect 13176 3068 13228 3077
rect 13360 3043 13412 3052
rect 13360 3009 13369 3043
rect 13369 3009 13403 3043
rect 13403 3009 13412 3043
rect 15752 3145 15761 3179
rect 15761 3145 15795 3179
rect 15795 3145 15804 3179
rect 15752 3136 15804 3145
rect 37556 3136 37608 3188
rect 13360 3000 13412 3009
rect 18696 3068 18748 3120
rect 18972 3111 19024 3120
rect 18972 3077 18981 3111
rect 18981 3077 19015 3111
rect 19015 3077 19024 3111
rect 18972 3068 19024 3077
rect 24584 3111 24636 3120
rect 24584 3077 24593 3111
rect 24593 3077 24627 3111
rect 24627 3077 24636 3111
rect 24584 3068 24636 3077
rect 29368 3111 29420 3120
rect 29368 3077 29377 3111
rect 29377 3077 29411 3111
rect 29411 3077 29420 3111
rect 29368 3068 29420 3077
rect 18788 3043 18840 3052
rect 11612 2975 11664 2984
rect 11612 2941 11621 2975
rect 11621 2941 11655 2975
rect 11655 2941 11664 2975
rect 11612 2932 11664 2941
rect 11704 2932 11756 2984
rect 18788 3009 18797 3043
rect 18797 3009 18831 3043
rect 18831 3009 18840 3043
rect 18788 3000 18840 3009
rect 22100 3043 22152 3052
rect 22100 3009 22109 3043
rect 22109 3009 22143 3043
rect 22143 3009 22152 3043
rect 22100 3000 22152 3009
rect 24400 3043 24452 3052
rect 24400 3009 24409 3043
rect 24409 3009 24443 3043
rect 24443 3009 24452 3043
rect 24400 3000 24452 3009
rect 29184 3043 29236 3052
rect 29184 3009 29193 3043
rect 29193 3009 29227 3043
rect 29227 3009 29236 3043
rect 29184 3000 29236 3009
rect 35624 3000 35676 3052
rect 36544 3043 36596 3052
rect 36544 3009 36553 3043
rect 36553 3009 36587 3043
rect 36587 3009 36596 3043
rect 36544 3000 36596 3009
rect 42984 3136 43036 3188
rect 40040 3043 40092 3052
rect 40040 3009 40049 3043
rect 40049 3009 40083 3043
rect 40083 3009 40092 3043
rect 40040 3000 40092 3009
rect 42892 3000 42944 3052
rect 44180 3000 44232 3052
rect 19340 2975 19392 2984
rect 19340 2941 19349 2975
rect 19349 2941 19383 2975
rect 19383 2941 19392 2975
rect 19340 2932 19392 2941
rect 22284 2975 22336 2984
rect 22284 2941 22293 2975
rect 22293 2941 22327 2975
rect 22327 2941 22336 2975
rect 22284 2932 22336 2941
rect 23204 2975 23256 2984
rect 23204 2941 23213 2975
rect 23213 2941 23247 2975
rect 23247 2941 23256 2975
rect 23204 2932 23256 2941
rect 25136 2975 25188 2984
rect 25136 2941 25145 2975
rect 25145 2941 25179 2975
rect 25179 2941 25188 2975
rect 25136 2932 25188 2941
rect 29644 2975 29696 2984
rect 29644 2941 29653 2975
rect 29653 2941 29687 2975
rect 29687 2941 29696 2975
rect 29644 2932 29696 2941
rect 40224 2975 40276 2984
rect 23020 2864 23072 2916
rect 1400 2796 1452 2848
rect 3240 2796 3292 2848
rect 3976 2796 4028 2848
rect 6552 2796 6604 2848
rect 17040 2839 17092 2848
rect 17040 2805 17049 2839
rect 17049 2805 17083 2839
rect 17083 2805 17092 2839
rect 17040 2796 17092 2805
rect 40224 2941 40233 2975
rect 40233 2941 40267 2975
rect 40267 2941 40276 2975
rect 40224 2932 40276 2941
rect 41236 2975 41288 2984
rect 41236 2941 41245 2975
rect 41245 2941 41279 2975
rect 41279 2941 41288 2975
rect 41236 2932 41288 2941
rect 43812 2796 43864 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 3424 2592 3476 2644
rect 15936 2592 15988 2644
rect 22284 2592 22336 2644
rect 42984 2635 43036 2644
rect 42984 2601 42993 2635
rect 42993 2601 43027 2635
rect 43027 2601 43036 2635
rect 42984 2592 43036 2601
rect 1400 2499 1452 2508
rect 1400 2465 1409 2499
rect 1409 2465 1443 2499
rect 1443 2465 1452 2499
rect 1400 2456 1452 2465
rect 1584 2499 1636 2508
rect 1584 2465 1593 2499
rect 1593 2465 1627 2499
rect 1627 2465 1636 2499
rect 1584 2456 1636 2465
rect 2780 2499 2832 2508
rect 2780 2465 2789 2499
rect 2789 2465 2823 2499
rect 2823 2465 2832 2499
rect 2780 2456 2832 2465
rect 3792 2499 3844 2508
rect 3792 2465 3801 2499
rect 3801 2465 3835 2499
rect 3835 2465 3844 2499
rect 3792 2456 3844 2465
rect 4620 2456 4672 2508
rect 4712 2499 4764 2508
rect 4712 2465 4721 2499
rect 4721 2465 4755 2499
rect 4755 2465 4764 2499
rect 6368 2499 6420 2508
rect 4712 2456 4764 2465
rect 6368 2465 6377 2499
rect 6377 2465 6411 2499
rect 6411 2465 6420 2499
rect 6368 2456 6420 2465
rect 6552 2499 6604 2508
rect 6552 2465 6561 2499
rect 6561 2465 6595 2499
rect 6595 2465 6604 2499
rect 6552 2456 6604 2465
rect 6644 2456 6696 2508
rect 12440 2524 12492 2576
rect 23020 2524 23072 2576
rect 43352 2524 43404 2576
rect 11888 2499 11940 2508
rect 11888 2465 11897 2499
rect 11897 2465 11931 2499
rect 11931 2465 11940 2499
rect 11888 2456 11940 2465
rect 12256 2499 12308 2508
rect 12256 2465 12265 2499
rect 12265 2465 12299 2499
rect 12299 2465 12308 2499
rect 12256 2456 12308 2465
rect 16856 2499 16908 2508
rect 16856 2465 16865 2499
rect 16865 2465 16899 2499
rect 16899 2465 16908 2499
rect 16856 2456 16908 2465
rect 17040 2499 17092 2508
rect 17040 2465 17049 2499
rect 17049 2465 17083 2499
rect 17083 2465 17092 2499
rect 17040 2456 17092 2465
rect 17408 2499 17460 2508
rect 17408 2465 17417 2499
rect 17417 2465 17451 2499
rect 17451 2465 17460 2499
rect 17408 2456 17460 2465
rect 24216 2456 24268 2508
rect 24584 2456 24636 2508
rect 37280 2499 37332 2508
rect 37280 2465 37289 2499
rect 37289 2465 37323 2499
rect 37323 2465 37332 2499
rect 37280 2456 37332 2465
rect 37464 2499 37516 2508
rect 37464 2465 37473 2499
rect 37473 2465 37507 2499
rect 37507 2465 37516 2499
rect 37464 2456 37516 2465
rect 38660 2499 38712 2508
rect 38660 2465 38669 2499
rect 38669 2465 38703 2499
rect 38703 2465 38712 2499
rect 38660 2456 38712 2465
rect 41328 2499 41380 2508
rect 41328 2465 41337 2499
rect 41337 2465 41371 2499
rect 41371 2465 41380 2499
rect 41328 2456 41380 2465
rect 43444 2456 43496 2508
rect 43536 2388 43588 2440
rect 23756 2320 23808 2372
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect -10 45200 102 46000
rect 634 45200 746 46000
rect 1922 45200 2034 46000
rect 2566 45200 2678 46000
rect 3210 45200 3322 46000
rect 4498 45200 4610 46000
rect 5142 45200 5254 46000
rect 5786 45200 5898 46000
rect 7074 45200 7186 46000
rect 7718 45200 7830 46000
rect 8362 45200 8474 46000
rect 9650 45200 9762 46000
rect 10294 45200 10406 46000
rect 10938 45200 11050 46000
rect 12226 45200 12338 46000
rect 12870 45200 12982 46000
rect 13514 45200 13626 46000
rect 14802 45200 14914 46000
rect 15446 45200 15558 46000
rect 16090 45200 16202 46000
rect 17378 45200 17490 46000
rect 18022 45200 18134 46000
rect 18666 45200 18778 46000
rect 19954 45200 20066 46000
rect 20598 45200 20710 46000
rect 21242 45200 21354 46000
rect 22530 45200 22642 46000
rect 23174 45200 23286 46000
rect 23818 45200 23930 46000
rect 24462 45200 24574 46000
rect 25750 45200 25862 46000
rect 26394 45200 26506 46000
rect 27038 45200 27150 46000
rect 28326 45200 28438 46000
rect 28970 45200 29082 46000
rect 29614 45200 29726 46000
rect 30902 45200 31014 46000
rect 31546 45200 31658 46000
rect 32190 45200 32302 46000
rect 33478 45200 33590 46000
rect 34122 45200 34234 46000
rect 34766 45200 34878 46000
rect 36054 45200 36166 46000
rect 36698 45200 36810 46000
rect 37342 45200 37454 46000
rect 38630 45200 38742 46000
rect 39274 45200 39386 46000
rect 39918 45200 40030 46000
rect 41206 45200 41318 46000
rect 41850 45200 41962 46000
rect 42494 45200 42606 46000
rect 43782 45200 43894 46000
rect 44426 45200 44538 46000
rect 45070 45200 45182 46000
rect 45714 45200 45826 46000
rect 1860 43308 1912 43314
rect 1860 43250 1912 43256
rect 1872 42945 1900 43250
rect 1964 43194 1992 45200
rect 1964 43178 2084 43194
rect 1964 43172 2096 43178
rect 1964 43166 2044 43172
rect 2044 43114 2096 43120
rect 1858 42936 1914 42945
rect 1858 42871 1914 42880
rect 2608 42362 2636 45200
rect 2870 44976 2926 44985
rect 2870 44911 2926 44920
rect 2780 43104 2832 43110
rect 2780 43046 2832 43052
rect 2596 42356 2648 42362
rect 2596 42298 2648 42304
rect 2792 42294 2820 43046
rect 2884 42770 2912 44911
rect 4540 43874 4568 45200
rect 4540 43846 4660 43874
rect 2962 43616 3018 43625
rect 2962 43551 3018 43560
rect 2872 42764 2924 42770
rect 2872 42706 2924 42712
rect 2780 42288 2832 42294
rect 2780 42230 2832 42236
rect 2870 42256 2926 42265
rect 2870 42191 2926 42200
rect 2884 42158 2912 42191
rect 1860 42152 1912 42158
rect 1860 42094 1912 42100
rect 2872 42152 2924 42158
rect 2872 42094 2924 42100
rect 1872 41138 1900 42094
rect 2976 41750 3004 43551
rect 3332 43308 3384 43314
rect 3332 43250 3384 43256
rect 3240 42696 3292 42702
rect 3240 42638 3292 42644
rect 3148 42560 3200 42566
rect 3148 42502 3200 42508
rect 2964 41744 3016 41750
rect 2964 41686 3016 41692
rect 2872 41676 2924 41682
rect 2872 41618 2924 41624
rect 1860 41132 1912 41138
rect 1860 41074 1912 41080
rect 2320 41064 2372 41070
rect 2320 41006 2372 41012
rect 2332 40662 2360 41006
rect 2884 40730 2912 41618
rect 3056 41540 3108 41546
rect 3056 41482 3108 41488
rect 3068 41274 3096 41482
rect 3056 41268 3108 41274
rect 3056 41210 3108 41216
rect 3160 41206 3188 42502
rect 3148 41200 3200 41206
rect 3148 41142 3200 41148
rect 3252 41138 3280 42638
rect 3240 41132 3292 41138
rect 3240 41074 3292 41080
rect 3344 41018 3372 43250
rect 3608 43240 3660 43246
rect 3608 43182 3660 43188
rect 3792 43240 3844 43246
rect 3792 43182 3844 43188
rect 3976 43240 4028 43246
rect 3976 43182 4028 43188
rect 3160 40990 3372 41018
rect 2872 40724 2924 40730
rect 2872 40666 2924 40672
rect 2320 40656 2372 40662
rect 2320 40598 2372 40604
rect 1952 40520 2004 40526
rect 1952 40462 2004 40468
rect 1964 40050 1992 40462
rect 1952 40044 2004 40050
rect 1952 39986 2004 39992
rect 1398 37496 1454 37505
rect 1398 37431 1454 37440
rect 1412 37262 1440 37431
rect 1400 37256 1452 37262
rect 1400 37198 1452 37204
rect 1768 30728 1820 30734
rect 1768 30670 1820 30676
rect 1780 30258 1808 30670
rect 1768 30252 1820 30258
rect 1768 30194 1820 30200
rect 2228 30184 2280 30190
rect 2228 30126 2280 30132
rect 2240 29850 2268 30126
rect 2228 29844 2280 29850
rect 2228 29786 2280 29792
rect 2136 23724 2188 23730
rect 2136 23666 2188 23672
rect 1398 23216 1454 23225
rect 1398 23151 1400 23160
rect 1452 23151 1454 23160
rect 1400 23122 1452 23128
rect 1952 22568 2004 22574
rect 1952 22510 2004 22516
rect 1964 22234 1992 22510
rect 1952 22228 2004 22234
rect 1952 22170 2004 22176
rect 1676 20936 1728 20942
rect 1676 20878 1728 20884
rect 1688 20466 1716 20878
rect 1676 20460 1728 20466
rect 1676 20402 1728 20408
rect 2044 20392 2096 20398
rect 2044 20334 2096 20340
rect 2056 20058 2084 20334
rect 2044 20052 2096 20058
rect 2044 19994 2096 20000
rect 2148 19854 2176 23666
rect 2136 19848 2188 19854
rect 2136 19790 2188 19796
rect 2044 18760 2096 18766
rect 2044 18702 2096 18708
rect 2056 18290 2084 18702
rect 2044 18284 2096 18290
rect 2044 18226 2096 18232
rect 1768 17672 1820 17678
rect 1768 17614 1820 17620
rect 1780 17202 1808 17614
rect 1768 17196 1820 17202
rect 1768 17138 1820 17144
rect 1952 17128 2004 17134
rect 1952 17070 2004 17076
rect 1964 16794 1992 17070
rect 1952 16788 2004 16794
rect 1952 16730 2004 16736
rect 1676 16584 1728 16590
rect 1676 16526 1728 16532
rect 1688 16114 1716 16526
rect 1676 16108 1728 16114
rect 1676 16050 1728 16056
rect 2228 16040 2280 16046
rect 2228 15982 2280 15988
rect 2240 15706 2268 15982
rect 2228 15700 2280 15706
rect 2228 15642 2280 15648
rect 2044 14408 2096 14414
rect 2044 14350 2096 14356
rect 2056 13938 2084 14350
rect 2228 14272 2280 14278
rect 2228 14214 2280 14220
rect 2240 14006 2268 14214
rect 2228 14000 2280 14006
rect 2228 13942 2280 13948
rect 2044 13932 2096 13938
rect 2044 13874 2096 13880
rect 1676 13320 1728 13326
rect 1676 13262 1728 13268
rect 1688 12850 1716 13262
rect 1676 12844 1728 12850
rect 1676 12786 1728 12792
rect 1860 12776 1912 12782
rect 1860 12718 1912 12724
rect 1872 12442 1900 12718
rect 1860 12436 1912 12442
rect 1860 12378 1912 12384
rect 1860 10464 1912 10470
rect 1860 10406 1912 10412
rect 2136 10464 2188 10470
rect 2136 10406 2188 10412
rect 1398 10296 1454 10305
rect 1398 10231 1454 10240
rect 1412 10130 1440 10231
rect 1400 10124 1452 10130
rect 1400 10066 1452 10072
rect 1872 8498 1900 10406
rect 1952 9512 2004 9518
rect 1952 9454 2004 9460
rect 1964 9178 1992 9454
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 2148 8566 2176 10406
rect 2136 8560 2188 8566
rect 2136 8502 2188 8508
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 1676 6792 1728 6798
rect 1676 6734 1728 6740
rect 1688 6322 1716 6734
rect 1676 6316 1728 6322
rect 1676 6258 1728 6264
rect 2136 6248 2188 6254
rect 2136 6190 2188 6196
rect 2148 5914 2176 6190
rect 2136 5908 2188 5914
rect 2136 5850 2188 5856
rect 1584 5704 1636 5710
rect 1584 5646 1636 5652
rect 2044 5704 2096 5710
rect 2044 5646 2096 5652
rect 1596 5234 1624 5646
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 2056 4146 2084 5646
rect 2044 4140 2096 4146
rect 2044 4082 2096 4088
rect 2332 4010 2360 40598
rect 2778 40216 2834 40225
rect 2778 40151 2834 40160
rect 2792 39982 2820 40151
rect 2872 40112 2924 40118
rect 2872 40054 2924 40060
rect 2780 39976 2832 39982
rect 2780 39918 2832 39924
rect 2884 39642 2912 40054
rect 2872 39636 2924 39642
rect 2872 39578 2924 39584
rect 2688 37188 2740 37194
rect 2688 37130 2740 37136
rect 2700 36922 2728 37130
rect 2688 36916 2740 36922
rect 2688 36858 2740 36864
rect 2780 30184 2832 30190
rect 2780 30126 2832 30132
rect 2792 30025 2820 30126
rect 2778 30016 2834 30025
rect 2778 29951 2834 29960
rect 2412 29640 2464 29646
rect 2412 29582 2464 29588
rect 2424 15502 2452 29582
rect 3056 23588 3108 23594
rect 3056 23530 3108 23536
rect 2780 23520 2832 23526
rect 2780 23462 2832 23468
rect 2792 23186 2820 23462
rect 2780 23180 2832 23186
rect 2780 23122 2832 23128
rect 3068 23050 3096 23530
rect 3056 23044 3108 23050
rect 3056 22986 3108 22992
rect 2872 22568 2924 22574
rect 2964 22568 3016 22574
rect 2872 22510 2924 22516
rect 2962 22536 2964 22545
rect 3016 22536 3018 22545
rect 2884 22098 2912 22510
rect 2962 22471 3018 22480
rect 3160 22098 3188 40990
rect 3620 40526 3648 43182
rect 3608 40520 3660 40526
rect 3608 40462 3660 40468
rect 3804 39642 3832 43182
rect 3988 41818 4016 43182
rect 4214 43004 4522 43024
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42928 4522 42948
rect 4632 42702 4660 43846
rect 4620 42696 4672 42702
rect 4620 42638 4672 42644
rect 4988 42220 5040 42226
rect 4988 42162 5040 42168
rect 4214 41916 4522 41936
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41840 4522 41860
rect 5000 41818 5028 42162
rect 3976 41812 4028 41818
rect 3976 41754 4028 41760
rect 4988 41812 5040 41818
rect 4988 41754 5040 41760
rect 4620 41608 4672 41614
rect 4620 41550 4672 41556
rect 4214 40828 4522 40848
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40752 4522 40772
rect 3884 40520 3936 40526
rect 3884 40462 3936 40468
rect 3792 39636 3844 39642
rect 3792 39578 3844 39584
rect 3330 38176 3386 38185
rect 3330 38111 3386 38120
rect 3240 37664 3292 37670
rect 3240 37606 3292 37612
rect 3252 37262 3280 37606
rect 3240 37256 3292 37262
rect 3240 37198 3292 37204
rect 3344 25974 3372 38111
rect 3332 25968 3384 25974
rect 3332 25910 3384 25916
rect 2872 22092 2924 22098
rect 2872 22034 2924 22040
rect 3148 22092 3200 22098
rect 3148 22034 3200 22040
rect 3896 20942 3924 40462
rect 4632 40186 4660 41550
rect 4712 41064 4764 41070
rect 4712 41006 4764 41012
rect 4620 40180 4672 40186
rect 4620 40122 4672 40128
rect 4632 39982 4660 40122
rect 4620 39976 4672 39982
rect 4620 39918 4672 39924
rect 4214 39740 4522 39760
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39664 4522 39684
rect 4214 38652 4522 38672
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38576 4522 38596
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 3976 25832 4028 25838
rect 3976 25774 4028 25780
rect 3988 25498 4016 25774
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 3976 25492 4028 25498
rect 3976 25434 4028 25440
rect 3976 25288 4028 25294
rect 3976 25230 4028 25236
rect 3988 22030 4016 25230
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 3976 22024 4028 22030
rect 3976 21966 4028 21972
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 3884 20936 3936 20942
rect 3884 20878 3936 20884
rect 2778 20496 2834 20505
rect 2778 20431 2834 20440
rect 2792 20398 2820 20431
rect 2780 20392 2832 20398
rect 2780 20334 2832 20340
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 3976 19848 4028 19854
rect 3976 19790 4028 19796
rect 2962 18456 3018 18465
rect 2962 18391 3018 18400
rect 2976 18222 3004 18391
rect 2872 18216 2924 18222
rect 2872 18158 2924 18164
rect 2964 18216 3016 18222
rect 2964 18158 3016 18164
rect 2884 17882 2912 18158
rect 2872 17876 2924 17882
rect 2872 17818 2924 17824
rect 2780 17128 2832 17134
rect 2778 17096 2780 17105
rect 2832 17096 2834 17105
rect 2778 17031 2834 17040
rect 2780 16040 2832 16046
rect 2780 15982 2832 15988
rect 2792 15745 2820 15982
rect 3424 15904 3476 15910
rect 3424 15846 3476 15852
rect 2778 15736 2834 15745
rect 2778 15671 2834 15680
rect 3436 15502 3464 15846
rect 2412 15496 2464 15502
rect 2412 15438 2464 15444
rect 3424 15496 3476 15502
rect 3424 15438 3476 15444
rect 2778 14376 2834 14385
rect 2778 14311 2834 14320
rect 2792 13870 2820 14311
rect 2780 13864 2832 13870
rect 2780 13806 2832 13812
rect 2778 13016 2834 13025
rect 2778 12951 2834 12960
rect 2792 12782 2820 12951
rect 2780 12776 2832 12782
rect 2780 12718 2832 12724
rect 3240 11144 3292 11150
rect 3240 11086 3292 11092
rect 2596 10668 2648 10674
rect 2596 10610 2648 10616
rect 2504 9512 2556 9518
rect 2504 9454 2556 9460
rect 2516 9178 2544 9454
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 2608 8974 2636 10610
rect 3252 10130 3280 11086
rect 3240 10124 3292 10130
rect 3240 10066 3292 10072
rect 2870 9616 2926 9625
rect 2870 9551 2926 9560
rect 2780 9512 2832 9518
rect 2780 9454 2832 9460
rect 2596 8968 2648 8974
rect 2792 8945 2820 9454
rect 2596 8910 2648 8916
rect 2778 8936 2834 8945
rect 2778 8871 2834 8880
rect 2884 8430 2912 9551
rect 2872 8424 2924 8430
rect 2872 8366 2924 8372
rect 3436 7410 3464 15438
rect 3988 10062 4016 19790
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 3976 10056 4028 10062
rect 3976 9998 4028 10004
rect 3988 9654 4016 9998
rect 3976 9648 4028 9654
rect 3976 9590 4028 9596
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 3424 7404 3476 7410
rect 3424 7346 3476 7352
rect 3516 7200 3568 7206
rect 3516 7142 3568 7148
rect 4068 7200 4120 7206
rect 4068 7142 4120 7148
rect 3528 6730 3556 7142
rect 3974 6896 4030 6905
rect 4080 6866 4108 7142
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 3974 6831 4030 6840
rect 4068 6860 4120 6866
rect 3988 6746 4016 6831
rect 4068 6802 4120 6808
rect 3988 6730 4108 6746
rect 3516 6724 3568 6730
rect 3988 6724 4120 6730
rect 3988 6718 4068 6724
rect 3516 6666 3568 6672
rect 4068 6666 4120 6672
rect 2780 6248 2832 6254
rect 2778 6216 2780 6225
rect 2832 6216 2834 6225
rect 2778 6151 2834 6160
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 2872 5568 2924 5574
rect 2872 5510 2924 5516
rect 2884 5302 2912 5510
rect 2872 5296 2924 5302
rect 2872 5238 2924 5244
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 2792 4865 2820 5102
rect 2778 4856 2834 4865
rect 2778 4791 2834 4800
rect 2964 4684 3016 4690
rect 2964 4626 3016 4632
rect 2778 4176 2834 4185
rect 2778 4111 2834 4120
rect 2792 4078 2820 4111
rect 2780 4072 2832 4078
rect 2780 4014 2832 4020
rect 2320 4004 2372 4010
rect 2320 3946 2372 3952
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 1400 3528 1452 3534
rect 1398 3496 1400 3505
rect 1452 3496 1454 3505
rect 1398 3431 1454 3440
rect 664 2916 716 2922
rect 664 2858 716 2864
rect 676 800 704 2858
rect 1400 2848 1452 2854
rect 1400 2790 1452 2796
rect 1412 2514 1440 2790
rect 1596 2514 1624 3878
rect 2228 3460 2280 3466
rect 2228 3402 2280 3408
rect 2240 3194 2268 3402
rect 2228 3188 2280 3194
rect 2228 3130 2280 3136
rect 2332 3058 2360 3946
rect 2976 3602 3004 4626
rect 3148 4616 3200 4622
rect 3148 4558 3200 4564
rect 2964 3596 3016 3602
rect 2964 3538 3016 3544
rect 3160 3058 3188 4558
rect 3700 3460 3752 3466
rect 3700 3402 3752 3408
rect 2320 3052 2372 3058
rect 2320 2994 2372 3000
rect 3148 3052 3200 3058
rect 3148 2994 3200 3000
rect 3712 2990 3740 3402
rect 3700 2984 3752 2990
rect 3700 2926 3752 2932
rect 3240 2848 3292 2854
rect 3240 2790 3292 2796
rect 1400 2508 1452 2514
rect 1400 2450 1452 2456
rect 1584 2508 1636 2514
rect 1584 2450 1636 2456
rect 2780 2508 2832 2514
rect 2780 2450 2832 2456
rect 2792 1465 2820 2450
rect 2778 1456 2834 1465
rect 2778 1391 2834 1400
rect 3252 800 3280 2790
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 3436 2145 3464 2586
rect 3804 2514 3832 5646
rect 4172 5114 4200 5646
rect 4632 5234 4660 39918
rect 4724 16574 4752 41006
rect 4804 40996 4856 41002
rect 4804 40938 4856 40944
rect 4816 39438 4844 40938
rect 4804 39432 4856 39438
rect 4804 39374 4856 39380
rect 4816 37942 4844 39374
rect 4804 37936 4856 37942
rect 4804 37878 4856 37884
rect 4816 35894 4844 37878
rect 4816 35866 4936 35894
rect 4724 16546 4844 16574
rect 4712 6860 4764 6866
rect 4712 6802 4764 6808
rect 4620 5228 4672 5234
rect 4620 5170 4672 5176
rect 4080 5086 4200 5114
rect 4080 4690 4108 5086
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 4632 4690 4660 4966
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 4620 4684 4672 4690
rect 4620 4626 4672 4632
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 4172 4078 4200 4422
rect 4160 4072 4212 4078
rect 4160 4014 4212 4020
rect 4724 3942 4752 6802
rect 4816 4826 4844 16546
rect 4908 12238 4936 35866
rect 4896 12232 4948 12238
rect 4896 12174 4948 12180
rect 5000 10674 5028 41754
rect 5184 41682 5212 45200
rect 7760 43314 7788 45200
rect 7748 43308 7800 43314
rect 7748 43250 7800 43256
rect 6552 43104 6604 43110
rect 6552 43046 6604 43052
rect 8024 43104 8076 43110
rect 8024 43046 8076 43052
rect 6460 42628 6512 42634
rect 6460 42570 6512 42576
rect 6368 42016 6420 42022
rect 6368 41958 6420 41964
rect 6380 41682 6408 41958
rect 5172 41676 5224 41682
rect 5172 41618 5224 41624
rect 6368 41676 6420 41682
rect 6368 41618 6420 41624
rect 6472 41274 6500 42570
rect 6564 41682 6592 43046
rect 7104 42696 7156 42702
rect 7104 42638 7156 42644
rect 7116 42158 7144 42638
rect 7104 42152 7156 42158
rect 7104 42094 7156 42100
rect 7472 42084 7524 42090
rect 7472 42026 7524 42032
rect 6552 41676 6604 41682
rect 6552 41618 6604 41624
rect 6460 41268 6512 41274
rect 6460 41210 6512 41216
rect 5632 41132 5684 41138
rect 5632 41074 5684 41080
rect 5644 40526 5672 41074
rect 6644 41064 6696 41070
rect 6644 41006 6696 41012
rect 5632 40520 5684 40526
rect 5632 40462 5684 40468
rect 5906 40488 5962 40497
rect 5644 40118 5672 40462
rect 5906 40423 5962 40432
rect 5920 40390 5948 40423
rect 5908 40384 5960 40390
rect 5908 40326 5960 40332
rect 5632 40112 5684 40118
rect 5632 40054 5684 40060
rect 5644 39438 5672 40054
rect 5632 39432 5684 39438
rect 5632 39374 5684 39380
rect 5172 26240 5224 26246
rect 5172 26182 5224 26188
rect 5184 25906 5212 26182
rect 5172 25900 5224 25906
rect 5172 25842 5224 25848
rect 5540 21548 5592 21554
rect 5540 21490 5592 21496
rect 5172 21480 5224 21486
rect 5172 21422 5224 21428
rect 4988 10668 5040 10674
rect 4988 10610 5040 10616
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 4804 4684 4856 4690
rect 4804 4626 4856 4632
rect 3884 3936 3936 3942
rect 3884 3878 3936 3884
rect 4712 3936 4764 3942
rect 4712 3878 4764 3884
rect 3792 2508 3844 2514
rect 3792 2450 3844 2456
rect 3422 2136 3478 2145
rect 3422 2071 3478 2080
rect 3896 800 3924 3878
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 4528 3528 4580 3534
rect 4528 3470 4580 3476
rect 4540 3194 4568 3470
rect 4620 3392 4672 3398
rect 4620 3334 4672 3340
rect 4528 3188 4580 3194
rect 4528 3130 4580 3136
rect 3976 2984 4028 2990
rect 3976 2926 4028 2932
rect 3988 2854 4016 2926
rect 3976 2848 4028 2854
rect 3976 2790 4028 2796
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 4632 2514 4660 3334
rect 4712 2916 4764 2922
rect 4712 2858 4764 2864
rect 4724 2514 4752 2858
rect 4620 2508 4672 2514
rect 4620 2450 4672 2456
rect 4712 2508 4764 2514
rect 4712 2450 4764 2456
rect 4816 2258 4844 4626
rect 4908 4146 4936 4966
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 5184 2922 5212 21422
rect 5552 21146 5580 21490
rect 5540 21140 5592 21146
rect 5540 21082 5592 21088
rect 5552 20942 5580 21082
rect 5540 20936 5592 20942
rect 5540 20878 5592 20884
rect 5920 5846 5948 40326
rect 6656 26234 6684 41006
rect 7484 40458 7512 42026
rect 7472 40452 7524 40458
rect 7472 40394 7524 40400
rect 7932 36780 7984 36786
rect 7932 36722 7984 36728
rect 6564 26206 6684 26234
rect 6368 22636 6420 22642
rect 6368 22578 6420 22584
rect 6184 22568 6236 22574
rect 6184 22510 6236 22516
rect 6196 22234 6224 22510
rect 6184 22228 6236 22234
rect 6184 22170 6236 22176
rect 6092 22092 6144 22098
rect 6092 22034 6144 22040
rect 6104 20346 6132 22034
rect 6196 22030 6224 22170
rect 6380 22030 6408 22578
rect 6184 22024 6236 22030
rect 6184 21966 6236 21972
rect 6368 22024 6420 22030
rect 6368 21966 6420 21972
rect 6380 21622 6408 21966
rect 6368 21616 6420 21622
rect 6368 21558 6420 21564
rect 6564 21486 6592 26206
rect 7944 21690 7972 36722
rect 8036 30666 8064 43046
rect 10336 42770 10364 45200
rect 11520 43104 11572 43110
rect 11520 43046 11572 43052
rect 11612 43104 11664 43110
rect 11612 43046 11664 43052
rect 10324 42764 10376 42770
rect 10324 42706 10376 42712
rect 9312 42696 9364 42702
rect 9312 42638 9364 42644
rect 9324 42226 9352 42638
rect 10048 42628 10100 42634
rect 10048 42570 10100 42576
rect 9312 42220 9364 42226
rect 9312 42162 9364 42168
rect 10060 41818 10088 42570
rect 11532 42226 11560 43046
rect 11624 42770 11652 43046
rect 12268 42770 12296 45200
rect 12532 43308 12584 43314
rect 12532 43250 12584 43256
rect 12440 43104 12492 43110
rect 12440 43046 12492 43052
rect 11612 42764 11664 42770
rect 11612 42706 11664 42712
rect 12256 42764 12308 42770
rect 12256 42706 12308 42712
rect 11796 42628 11848 42634
rect 11796 42570 11848 42576
rect 11808 42362 11836 42570
rect 11796 42356 11848 42362
rect 11796 42298 11848 42304
rect 12452 42294 12480 43046
rect 12544 42566 12572 43250
rect 12532 42560 12584 42566
rect 12532 42502 12584 42508
rect 12440 42288 12492 42294
rect 12440 42230 12492 42236
rect 11520 42220 11572 42226
rect 11520 42162 11572 42168
rect 10048 41812 10100 41818
rect 10048 41754 10100 41760
rect 12164 41744 12216 41750
rect 12164 41686 12216 41692
rect 12072 41608 12124 41614
rect 12072 41550 12124 41556
rect 10968 41540 11020 41546
rect 10968 41482 11020 41488
rect 9312 41200 9364 41206
rect 9312 41142 9364 41148
rect 9324 40526 9352 41142
rect 10692 41132 10744 41138
rect 10692 41074 10744 41080
rect 9588 41064 9640 41070
rect 9588 41006 9640 41012
rect 9600 40934 9628 41006
rect 9588 40928 9640 40934
rect 9588 40870 9640 40876
rect 8852 40520 8904 40526
rect 8852 40462 8904 40468
rect 9312 40520 9364 40526
rect 9312 40462 9364 40468
rect 8024 30660 8076 30666
rect 8024 30602 8076 30608
rect 7932 21684 7984 21690
rect 7932 21626 7984 21632
rect 8208 21684 8260 21690
rect 8208 21626 8260 21632
rect 6552 21480 6604 21486
rect 6552 21422 6604 21428
rect 6828 21004 6880 21010
rect 6828 20946 6880 20952
rect 6104 20318 6224 20346
rect 6196 16658 6224 20318
rect 6840 18426 6868 20946
rect 8220 20262 8248 21626
rect 8208 20256 8260 20262
rect 8208 20198 8260 20204
rect 6276 18420 6328 18426
rect 6276 18362 6328 18368
rect 6828 18420 6880 18426
rect 6828 18362 6880 18368
rect 6184 16652 6236 16658
rect 6184 16594 6236 16600
rect 5908 5840 5960 5846
rect 5908 5782 5960 5788
rect 6196 4010 6224 16594
rect 6288 5778 6316 18362
rect 6276 5772 6328 5778
rect 6276 5714 6328 5720
rect 6276 4616 6328 4622
rect 6276 4558 6328 4564
rect 6184 4004 6236 4010
rect 6184 3946 6236 3952
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5552 3602 5580 3878
rect 5540 3596 5592 3602
rect 5540 3538 5592 3544
rect 5816 3596 5868 3602
rect 5816 3538 5868 3544
rect 5172 2916 5224 2922
rect 5172 2858 5224 2864
rect 4540 2230 4844 2258
rect 4540 800 4568 2230
rect 5828 800 5856 3538
rect 6288 2774 6316 4558
rect 6368 3936 6420 3942
rect 6368 3878 6420 3884
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 6380 3670 6408 3878
rect 6368 3664 6420 3670
rect 6368 3606 6420 3612
rect 7300 3058 7328 3878
rect 8220 3641 8248 20198
rect 8864 19922 8892 40462
rect 8852 19916 8904 19922
rect 8852 19858 8904 19864
rect 9220 14408 9272 14414
rect 9220 14350 9272 14356
rect 9232 12850 9260 14350
rect 9220 12844 9272 12850
rect 9220 12786 9272 12792
rect 9404 12640 9456 12646
rect 9404 12582 9456 12588
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 8206 3632 8262 3641
rect 9232 3602 9260 3878
rect 9416 3602 9444 12582
rect 9496 4004 9548 4010
rect 9496 3946 9548 3952
rect 9508 3670 9536 3946
rect 9496 3664 9548 3670
rect 9496 3606 9548 3612
rect 8206 3567 8262 3576
rect 9220 3596 9272 3602
rect 9220 3538 9272 3544
rect 9404 3596 9456 3602
rect 9404 3538 9456 3544
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 7484 3126 7512 3334
rect 9600 3194 9628 40870
rect 10704 40594 10732 41074
rect 10692 40588 10744 40594
rect 10692 40530 10744 40536
rect 10140 40452 10192 40458
rect 10140 40394 10192 40400
rect 10152 39506 10180 40394
rect 10140 39500 10192 39506
rect 10140 39442 10192 39448
rect 10980 23730 11008 41482
rect 12084 41138 12112 41550
rect 11060 41132 11112 41138
rect 11060 41074 11112 41080
rect 12072 41132 12124 41138
rect 12072 41074 12124 41080
rect 11072 41002 11100 41074
rect 11060 40996 11112 41002
rect 11060 40938 11112 40944
rect 12084 40526 12112 41074
rect 12072 40520 12124 40526
rect 12072 40462 12124 40468
rect 12084 40118 12112 40462
rect 12072 40112 12124 40118
rect 12072 40054 12124 40060
rect 12176 39982 12204 41686
rect 12544 41274 12572 42502
rect 12912 42158 12940 45200
rect 13084 43308 13136 43314
rect 13084 43250 13136 43256
rect 13096 42906 13124 43250
rect 13556 43178 13584 45200
rect 14096 43240 14148 43246
rect 14096 43182 14148 43188
rect 13544 43172 13596 43178
rect 13544 43114 13596 43120
rect 13084 42900 13136 42906
rect 13084 42842 13136 42848
rect 12900 42152 12952 42158
rect 12900 42094 12952 42100
rect 12992 41540 13044 41546
rect 12992 41482 13044 41488
rect 12532 41268 12584 41274
rect 12532 41210 12584 41216
rect 12164 39976 12216 39982
rect 12164 39918 12216 39924
rect 12176 33862 12204 39918
rect 12164 33856 12216 33862
rect 12164 33798 12216 33804
rect 10968 23724 11020 23730
rect 10968 23666 11020 23672
rect 11520 20800 11572 20806
rect 11520 20742 11572 20748
rect 11532 20466 11560 20742
rect 11520 20460 11572 20466
rect 11520 20402 11572 20408
rect 12256 20460 12308 20466
rect 12256 20402 12308 20408
rect 12268 19854 12296 20402
rect 12532 20392 12584 20398
rect 12532 20334 12584 20340
rect 12256 19848 12308 19854
rect 12256 19790 12308 19796
rect 12268 19378 12296 19790
rect 12256 19372 12308 19378
rect 12256 19314 12308 19320
rect 11704 18692 11756 18698
rect 11704 18634 11756 18640
rect 11716 17678 11744 18634
rect 11704 17672 11756 17678
rect 11704 17614 11756 17620
rect 9680 3596 9732 3602
rect 9680 3538 9732 3544
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 7472 3120 7524 3126
rect 7472 3062 7524 3068
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 7104 2984 7156 2990
rect 7104 2926 7156 2932
rect 6552 2848 6604 2854
rect 6552 2790 6604 2796
rect 6288 2746 6408 2774
rect 6380 2514 6408 2746
rect 6564 2514 6592 2790
rect 6368 2508 6420 2514
rect 6368 2450 6420 2456
rect 6552 2508 6604 2514
rect 6552 2450 6604 2456
rect 6644 2508 6696 2514
rect 6644 2450 6696 2456
rect 6656 1306 6684 2450
rect 6472 1278 6684 1306
rect 6472 800 6500 1278
rect 7116 800 7144 2926
rect 9692 800 9720 3538
rect 11716 2990 11744 17614
rect 12544 15910 12572 20334
rect 12808 19780 12860 19786
rect 12808 19722 12860 19728
rect 12716 19440 12768 19446
rect 12716 19382 12768 19388
rect 12624 19372 12676 19378
rect 12624 19314 12676 19320
rect 12636 18766 12664 19314
rect 12624 18760 12676 18766
rect 12624 18702 12676 18708
rect 12532 15904 12584 15910
rect 12532 15846 12584 15852
rect 12728 12850 12756 19382
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 11796 4752 11848 4758
rect 11796 4694 11848 4700
rect 11808 4146 11836 4694
rect 11796 4140 11848 4146
rect 11796 4082 11848 4088
rect 11888 3936 11940 3942
rect 11888 3878 11940 3884
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 11612 2984 11664 2990
rect 11612 2926 11664 2932
rect 11704 2984 11756 2990
rect 11704 2926 11756 2932
rect 11624 800 11652 2926
rect 11900 2514 11928 3878
rect 12452 2582 12480 3878
rect 12820 3738 12848 19722
rect 12900 16448 12952 16454
rect 12900 16390 12952 16396
rect 12912 16114 12940 16390
rect 12900 16108 12952 16114
rect 12900 16050 12952 16056
rect 12808 3732 12860 3738
rect 12808 3674 12860 3680
rect 13004 3602 13032 41482
rect 13096 40186 13124 42842
rect 14004 42084 14056 42090
rect 14004 42026 14056 42032
rect 14016 41138 14044 42026
rect 14004 41132 14056 41138
rect 14004 41074 14056 41080
rect 13268 40928 13320 40934
rect 13268 40870 13320 40876
rect 13084 40180 13136 40186
rect 13084 40122 13136 40128
rect 13176 16040 13228 16046
rect 13176 15982 13228 15988
rect 13188 15706 13216 15982
rect 13176 15700 13228 15706
rect 13176 15642 13228 15648
rect 13280 6914 13308 40870
rect 13912 33040 13964 33046
rect 13912 32982 13964 32988
rect 13924 31822 13952 32982
rect 13912 31816 13964 31822
rect 13912 31758 13964 31764
rect 13924 31278 13952 31758
rect 14016 31754 14044 41074
rect 14108 40730 14136 43182
rect 14844 42770 14872 45200
rect 19574 43548 19882 43568
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43472 19882 43492
rect 20812 43104 20864 43110
rect 20812 43046 20864 43052
rect 20824 42770 20852 43046
rect 21284 42770 21312 45200
rect 22652 43104 22704 43110
rect 22652 43046 22704 43052
rect 22560 42900 22612 42906
rect 22560 42842 22612 42848
rect 14832 42764 14884 42770
rect 14832 42706 14884 42712
rect 20812 42764 20864 42770
rect 20812 42706 20864 42712
rect 21272 42764 21324 42770
rect 21272 42706 21324 42712
rect 14372 42696 14424 42702
rect 14372 42638 14424 42644
rect 15752 42696 15804 42702
rect 15752 42638 15804 42644
rect 14384 41750 14412 42638
rect 14556 42628 14608 42634
rect 14556 42570 14608 42576
rect 14464 42152 14516 42158
rect 14464 42094 14516 42100
rect 14372 41744 14424 41750
rect 14372 41686 14424 41692
rect 14476 41274 14504 42094
rect 14568 41818 14596 42570
rect 15764 42294 15792 42638
rect 20996 42628 21048 42634
rect 20996 42570 21048 42576
rect 19574 42460 19882 42480
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42384 19882 42404
rect 21008 42362 21036 42570
rect 20996 42356 21048 42362
rect 20996 42298 21048 42304
rect 15752 42288 15804 42294
rect 15752 42230 15804 42236
rect 20812 42220 20864 42226
rect 20812 42162 20864 42168
rect 20824 42090 20852 42162
rect 20812 42084 20864 42090
rect 20812 42026 20864 42032
rect 14556 41812 14608 41818
rect 14556 41754 14608 41760
rect 14648 41608 14700 41614
rect 14648 41550 14700 41556
rect 14464 41268 14516 41274
rect 14464 41210 14516 41216
rect 14660 41138 14688 41550
rect 19574 41372 19882 41392
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41296 19882 41316
rect 14648 41132 14700 41138
rect 14648 41074 14700 41080
rect 14096 40724 14148 40730
rect 14096 40666 14148 40672
rect 14660 40458 14688 41074
rect 14648 40452 14700 40458
rect 14648 40394 14700 40400
rect 20824 40390 20852 42026
rect 22572 41614 22600 42842
rect 22664 42226 22692 43046
rect 22652 42220 22704 42226
rect 22652 42162 22704 42168
rect 23216 42158 23244 45200
rect 23860 44130 23888 45200
rect 23848 44124 23900 44130
rect 23848 44066 23900 44072
rect 23480 43376 23532 43382
rect 23480 43318 23532 43324
rect 22836 42152 22888 42158
rect 22836 42094 22888 42100
rect 23204 42152 23256 42158
rect 23204 42094 23256 42100
rect 22848 41818 22876 42094
rect 23492 41818 23520 43318
rect 24504 42838 24532 45200
rect 24860 44124 24912 44130
rect 24860 44066 24912 44072
rect 24872 43246 24900 44066
rect 25792 43382 25820 45200
rect 25780 43376 25832 43382
rect 25780 43318 25832 43324
rect 24860 43240 24912 43246
rect 24860 43182 24912 43188
rect 24492 42832 24544 42838
rect 24492 42774 24544 42780
rect 27080 42770 27108 45200
rect 27160 43104 27212 43110
rect 27160 43046 27212 43052
rect 27804 43104 27856 43110
rect 27804 43046 27856 43052
rect 27068 42764 27120 42770
rect 27068 42706 27120 42712
rect 26424 42696 26476 42702
rect 26424 42638 26476 42644
rect 24584 42628 24636 42634
rect 24584 42570 24636 42576
rect 24596 41818 24624 42570
rect 26436 42226 26464 42638
rect 27068 42628 27120 42634
rect 27068 42570 27120 42576
rect 27080 42362 27108 42570
rect 27068 42356 27120 42362
rect 27068 42298 27120 42304
rect 26424 42220 26476 42226
rect 26424 42162 26476 42168
rect 27068 42084 27120 42090
rect 27068 42026 27120 42032
rect 22836 41812 22888 41818
rect 22836 41754 22888 41760
rect 23480 41812 23532 41818
rect 23480 41754 23532 41760
rect 24584 41812 24636 41818
rect 24584 41754 24636 41760
rect 27080 41682 27108 42026
rect 27068 41676 27120 41682
rect 27068 41618 27120 41624
rect 22560 41608 22612 41614
rect 22560 41550 22612 41556
rect 22836 41608 22888 41614
rect 22836 41550 22888 41556
rect 24400 41608 24452 41614
rect 24400 41550 24452 41556
rect 20812 40384 20864 40390
rect 20812 40326 20864 40332
rect 19574 40284 19882 40304
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40208 19882 40228
rect 19248 40044 19300 40050
rect 19248 39986 19300 39992
rect 20536 40044 20588 40050
rect 20536 39986 20588 39992
rect 16396 39976 16448 39982
rect 16396 39918 16448 39924
rect 18696 39976 18748 39982
rect 18696 39918 18748 39924
rect 16408 38350 16436 39918
rect 18708 39506 18736 39918
rect 19260 39642 19288 39986
rect 19984 39840 20036 39846
rect 19984 39782 20036 39788
rect 19248 39636 19300 39642
rect 19248 39578 19300 39584
rect 18696 39500 18748 39506
rect 18696 39442 18748 39448
rect 19996 39438 20024 39782
rect 19984 39432 20036 39438
rect 19984 39374 20036 39380
rect 19574 39196 19882 39216
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39120 19882 39140
rect 16948 38956 17000 38962
rect 16948 38898 17000 38904
rect 18420 38956 18472 38962
rect 18420 38898 18472 38904
rect 16764 38888 16816 38894
rect 16764 38830 16816 38836
rect 15844 38344 15896 38350
rect 15844 38286 15896 38292
rect 16396 38344 16448 38350
rect 16396 38286 16448 38292
rect 15856 36174 15884 38286
rect 16672 36576 16724 36582
rect 16672 36518 16724 36524
rect 16684 36174 16712 36518
rect 15844 36168 15896 36174
rect 15844 36110 15896 36116
rect 16672 36168 16724 36174
rect 16672 36110 16724 36116
rect 15856 34542 15884 36110
rect 15384 34536 15436 34542
rect 15384 34478 15436 34484
rect 15844 34536 15896 34542
rect 15844 34478 15896 34484
rect 15396 34066 15424 34478
rect 15384 34060 15436 34066
rect 15384 34002 15436 34008
rect 16212 33924 16264 33930
rect 16212 33866 16264 33872
rect 16224 33114 16252 33866
rect 16488 33380 16540 33386
rect 16488 33322 16540 33328
rect 16212 33108 16264 33114
rect 16212 33050 16264 33056
rect 16396 32972 16448 32978
rect 16396 32914 16448 32920
rect 15752 32904 15804 32910
rect 15752 32846 15804 32852
rect 15568 32428 15620 32434
rect 15568 32370 15620 32376
rect 14372 32224 14424 32230
rect 14372 32166 14424 32172
rect 14384 31754 14412 32166
rect 15580 31958 15608 32370
rect 15568 31952 15620 31958
rect 15568 31894 15620 31900
rect 14016 31726 14136 31754
rect 13912 31272 13964 31278
rect 13912 31214 13964 31220
rect 13924 29306 13952 31214
rect 13912 29300 13964 29306
rect 13912 29242 13964 29248
rect 14108 20466 14136 31726
rect 14372 31748 14424 31754
rect 14372 31690 14424 31696
rect 15580 31482 15608 31894
rect 15568 31476 15620 31482
rect 15568 31418 15620 31424
rect 15476 31340 15528 31346
rect 15476 31282 15528 31288
rect 15488 30938 15516 31282
rect 15476 30932 15528 30938
rect 15476 30874 15528 30880
rect 15580 29714 15608 31418
rect 15764 31346 15792 32846
rect 16408 32722 16436 32914
rect 16500 32910 16528 33322
rect 16672 33312 16724 33318
rect 16672 33254 16724 33260
rect 16684 32910 16712 33254
rect 16488 32904 16540 32910
rect 16488 32846 16540 32852
rect 16672 32904 16724 32910
rect 16672 32846 16724 32852
rect 16408 32694 16528 32722
rect 16396 32496 16448 32502
rect 16396 32438 16448 32444
rect 15936 32428 15988 32434
rect 16212 32428 16264 32434
rect 15936 32370 15988 32376
rect 16132 32388 16212 32416
rect 15948 31754 15976 32370
rect 16028 32360 16080 32366
rect 16028 32302 16080 32308
rect 15856 31726 15976 31754
rect 15752 31340 15804 31346
rect 15752 31282 15804 31288
rect 15856 31210 15884 31726
rect 15936 31680 15988 31686
rect 15936 31622 15988 31628
rect 15844 31204 15896 31210
rect 15844 31146 15896 31152
rect 15856 30870 15884 31146
rect 15844 30864 15896 30870
rect 15844 30806 15896 30812
rect 15948 30734 15976 31622
rect 16040 30802 16068 32302
rect 16132 31890 16160 32388
rect 16212 32370 16264 32376
rect 16408 32366 16436 32438
rect 16500 32366 16528 32694
rect 16776 32570 16804 38830
rect 16856 38752 16908 38758
rect 16856 38694 16908 38700
rect 16868 38350 16896 38694
rect 16856 38344 16908 38350
rect 16856 38286 16908 38292
rect 16960 38010 16988 38898
rect 17316 38208 17368 38214
rect 17316 38150 17368 38156
rect 16948 38004 17000 38010
rect 16948 37946 17000 37952
rect 17328 37806 17356 38150
rect 18432 38010 18460 38898
rect 19996 38842 20024 39374
rect 20444 39364 20496 39370
rect 20444 39306 20496 39312
rect 20076 39296 20128 39302
rect 20076 39238 20128 39244
rect 20088 38962 20116 39238
rect 20076 38956 20128 38962
rect 20076 38898 20128 38904
rect 19996 38814 20116 38842
rect 19340 38752 19392 38758
rect 19340 38694 19392 38700
rect 19352 38554 19380 38694
rect 19340 38548 19392 38554
rect 19340 38490 19392 38496
rect 20088 38350 20116 38814
rect 20260 38412 20312 38418
rect 20260 38354 20312 38360
rect 20076 38344 20128 38350
rect 20076 38286 20128 38292
rect 19432 38276 19484 38282
rect 19432 38218 19484 38224
rect 18420 38004 18472 38010
rect 18420 37946 18472 37952
rect 19340 38004 19392 38010
rect 19340 37946 19392 37952
rect 19352 37913 19380 37946
rect 19338 37904 19394 37913
rect 17592 37868 17644 37874
rect 17592 37810 17644 37816
rect 18604 37868 18656 37874
rect 18604 37810 18656 37816
rect 18880 37868 18932 37874
rect 19338 37839 19394 37848
rect 18880 37810 18932 37816
rect 17316 37800 17368 37806
rect 17316 37742 17368 37748
rect 17132 37664 17184 37670
rect 17132 37606 17184 37612
rect 17144 36650 17172 37606
rect 17328 37262 17356 37742
rect 17316 37256 17368 37262
rect 17316 37198 17368 37204
rect 17604 37194 17632 37810
rect 18616 37262 18644 37810
rect 18892 37466 18920 37810
rect 19340 37800 19392 37806
rect 19340 37742 19392 37748
rect 18880 37460 18932 37466
rect 18880 37402 18932 37408
rect 17776 37256 17828 37262
rect 17776 37198 17828 37204
rect 18604 37256 18656 37262
rect 18604 37198 18656 37204
rect 17592 37188 17644 37194
rect 17592 37130 17644 37136
rect 17604 36718 17632 37130
rect 17592 36712 17644 36718
rect 17592 36654 17644 36660
rect 16856 36644 16908 36650
rect 16856 36586 16908 36592
rect 17132 36644 17184 36650
rect 17132 36586 17184 36592
rect 16764 32564 16816 32570
rect 16764 32506 16816 32512
rect 16396 32360 16448 32366
rect 16396 32302 16448 32308
rect 16488 32360 16540 32366
rect 16488 32302 16540 32308
rect 16212 32224 16264 32230
rect 16212 32166 16264 32172
rect 16120 31884 16172 31890
rect 16120 31826 16172 31832
rect 16132 31346 16160 31826
rect 16120 31340 16172 31346
rect 16120 31282 16172 31288
rect 16028 30796 16080 30802
rect 16028 30738 16080 30744
rect 15936 30728 15988 30734
rect 15936 30670 15988 30676
rect 15844 30184 15896 30190
rect 15844 30126 15896 30132
rect 15856 29850 15884 30126
rect 15844 29844 15896 29850
rect 15844 29786 15896 29792
rect 15568 29708 15620 29714
rect 15568 29650 15620 29656
rect 14464 29640 14516 29646
rect 14464 29582 14516 29588
rect 14188 29504 14240 29510
rect 14188 29446 14240 29452
rect 14200 29170 14228 29446
rect 14280 29232 14332 29238
rect 14280 29174 14332 29180
rect 14188 29164 14240 29170
rect 14188 29106 14240 29112
rect 14292 28558 14320 29174
rect 14280 28552 14332 28558
rect 14280 28494 14332 28500
rect 14292 26994 14320 28494
rect 14476 28218 14504 29582
rect 15200 29028 15252 29034
rect 15200 28970 15252 28976
rect 15212 28762 15240 28970
rect 16224 28778 16252 32166
rect 16500 31940 16528 32302
rect 16776 32230 16804 32506
rect 16764 32224 16816 32230
rect 16764 32166 16816 32172
rect 16672 32020 16724 32026
rect 16672 31962 16724 31968
rect 16500 31912 16620 31940
rect 16488 31816 16540 31822
rect 16488 31758 16540 31764
rect 16396 31272 16448 31278
rect 16396 31214 16448 31220
rect 16408 30870 16436 31214
rect 16500 31142 16528 31758
rect 16592 31754 16620 31912
rect 16684 31754 16712 31962
rect 16580 31748 16632 31754
rect 16580 31690 16632 31696
rect 16672 31748 16724 31754
rect 16672 31690 16724 31696
rect 16684 31346 16712 31690
rect 16672 31340 16724 31346
rect 16672 31282 16724 31288
rect 16488 31136 16540 31142
rect 16488 31078 16540 31084
rect 16396 30864 16448 30870
rect 16396 30806 16448 30812
rect 16500 30734 16528 31078
rect 16672 30932 16724 30938
rect 16672 30874 16724 30880
rect 16488 30728 16540 30734
rect 16488 30670 16540 30676
rect 16684 30326 16712 30874
rect 16868 30802 16896 36586
rect 17604 36106 17632 36654
rect 17788 36174 17816 37198
rect 18420 36780 18472 36786
rect 18420 36722 18472 36728
rect 18432 36582 18460 36722
rect 18420 36576 18472 36582
rect 18420 36518 18472 36524
rect 18432 36174 18460 36518
rect 18616 36378 18644 37198
rect 18892 36854 18920 37402
rect 19352 36854 19380 37742
rect 19444 37738 19472 38218
rect 19574 38108 19882 38128
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38032 19882 38052
rect 19522 37904 19578 37913
rect 19522 37839 19524 37848
rect 19576 37839 19578 37848
rect 19524 37810 19576 37816
rect 19432 37732 19484 37738
rect 19432 37674 19484 37680
rect 19524 37664 19576 37670
rect 19524 37606 19576 37612
rect 19536 37330 19564 37606
rect 19524 37324 19576 37330
rect 19524 37266 19576 37272
rect 19536 37210 19564 37266
rect 19444 37182 19564 37210
rect 18880 36848 18932 36854
rect 18880 36790 18932 36796
rect 19340 36848 19392 36854
rect 19340 36790 19392 36796
rect 19444 36650 19472 37182
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 19432 36644 19484 36650
rect 19432 36586 19484 36592
rect 19892 36644 19944 36650
rect 19892 36586 19944 36592
rect 18604 36372 18656 36378
rect 18604 36314 18656 36320
rect 18696 36236 18748 36242
rect 18696 36178 18748 36184
rect 17776 36168 17828 36174
rect 17776 36110 17828 36116
rect 18420 36168 18472 36174
rect 18420 36110 18472 36116
rect 17592 36100 17644 36106
rect 17592 36042 17644 36048
rect 18604 36100 18656 36106
rect 18604 36042 18656 36048
rect 18616 35630 18644 36042
rect 18604 35624 18656 35630
rect 18604 35566 18656 35572
rect 18708 35442 18736 36178
rect 19904 36174 19932 36586
rect 20088 36310 20116 38286
rect 20272 38214 20300 38354
rect 20352 38276 20404 38282
rect 20352 38218 20404 38224
rect 20260 38208 20312 38214
rect 20260 38150 20312 38156
rect 20272 37806 20300 38150
rect 20260 37800 20312 37806
rect 20180 37748 20260 37754
rect 20180 37742 20312 37748
rect 20180 37726 20300 37742
rect 20180 37262 20208 37726
rect 20260 37664 20312 37670
rect 20260 37606 20312 37612
rect 20168 37256 20220 37262
rect 20168 37198 20220 37204
rect 20272 36922 20300 37606
rect 20364 36922 20392 38218
rect 20456 38010 20484 39306
rect 20548 39098 20576 39986
rect 20720 39840 20772 39846
rect 20720 39782 20772 39788
rect 20732 39370 20760 39782
rect 21640 39432 21692 39438
rect 21640 39374 21692 39380
rect 20720 39364 20772 39370
rect 20720 39306 20772 39312
rect 20812 39296 20864 39302
rect 20812 39238 20864 39244
rect 20536 39092 20588 39098
rect 20536 39034 20588 39040
rect 20824 38894 20852 39238
rect 21652 38894 21680 39374
rect 22192 38956 22244 38962
rect 22192 38898 22244 38904
rect 20812 38888 20864 38894
rect 20812 38830 20864 38836
rect 21640 38888 21692 38894
rect 21640 38830 21692 38836
rect 20444 38004 20496 38010
rect 20444 37946 20496 37952
rect 20536 37256 20588 37262
rect 20536 37198 20588 37204
rect 20260 36916 20312 36922
rect 20260 36858 20312 36864
rect 20352 36916 20404 36922
rect 20352 36858 20404 36864
rect 20364 36802 20392 36858
rect 20272 36786 20392 36802
rect 20260 36780 20392 36786
rect 20312 36774 20392 36780
rect 20444 36780 20496 36786
rect 20260 36722 20312 36728
rect 20444 36722 20496 36728
rect 20076 36304 20128 36310
rect 20076 36246 20128 36252
rect 19892 36168 19944 36174
rect 19892 36110 19944 36116
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 20088 35630 20116 36246
rect 20456 35834 20484 36722
rect 20548 36378 20576 37198
rect 20628 36780 20680 36786
rect 20628 36722 20680 36728
rect 20720 36780 20772 36786
rect 20720 36722 20772 36728
rect 20536 36372 20588 36378
rect 20536 36314 20588 36320
rect 20640 36038 20668 36722
rect 20732 36106 20760 36722
rect 20824 36718 20852 38830
rect 21652 38418 21680 38830
rect 22204 38554 22232 38898
rect 22192 38548 22244 38554
rect 22192 38490 22244 38496
rect 21640 38412 21692 38418
rect 21640 38354 21692 38360
rect 21548 38344 21600 38350
rect 21468 38292 21548 38298
rect 21468 38286 21600 38292
rect 21272 38276 21324 38282
rect 21272 38218 21324 38224
rect 21468 38270 21588 38286
rect 21284 38010 21312 38218
rect 21272 38004 21324 38010
rect 21272 37946 21324 37952
rect 21468 37806 21496 38270
rect 21652 37874 21680 38354
rect 21640 37868 21692 37874
rect 21640 37810 21692 37816
rect 21456 37800 21508 37806
rect 21456 37742 21508 37748
rect 21180 37120 21232 37126
rect 21180 37062 21232 37068
rect 21192 36854 21220 37062
rect 21180 36848 21232 36854
rect 21180 36790 21232 36796
rect 20812 36712 20864 36718
rect 20812 36654 20864 36660
rect 20812 36576 20864 36582
rect 20812 36518 20864 36524
rect 20824 36242 20852 36518
rect 20812 36236 20864 36242
rect 20812 36178 20864 36184
rect 21192 36174 21220 36790
rect 20996 36168 21048 36174
rect 20996 36110 21048 36116
rect 21180 36168 21232 36174
rect 21180 36110 21232 36116
rect 20720 36100 20772 36106
rect 20720 36042 20772 36048
rect 20628 36032 20680 36038
rect 20628 35974 20680 35980
rect 20444 35828 20496 35834
rect 20444 35770 20496 35776
rect 20076 35624 20128 35630
rect 20076 35566 20128 35572
rect 18616 35414 18736 35442
rect 17224 35012 17276 35018
rect 17224 34954 17276 34960
rect 17408 35012 17460 35018
rect 17408 34954 17460 34960
rect 17236 34202 17264 34954
rect 17420 34746 17448 34954
rect 17592 34944 17644 34950
rect 17592 34886 17644 34892
rect 17408 34740 17460 34746
rect 17408 34682 17460 34688
rect 16948 34196 17000 34202
rect 16948 34138 17000 34144
rect 17224 34196 17276 34202
rect 17224 34138 17276 34144
rect 16960 33522 16988 34138
rect 17420 34066 17448 34682
rect 17408 34060 17460 34066
rect 17408 34002 17460 34008
rect 17604 33522 17632 34886
rect 17868 33992 17920 33998
rect 17868 33934 17920 33940
rect 16948 33516 17000 33522
rect 16948 33458 17000 33464
rect 17592 33516 17644 33522
rect 17592 33458 17644 33464
rect 17776 33516 17828 33522
rect 17776 33458 17828 33464
rect 17788 31822 17816 33458
rect 17880 33454 17908 33934
rect 18616 33658 18644 35414
rect 19984 35080 20036 35086
rect 19984 35022 20036 35028
rect 19432 34944 19484 34950
rect 19432 34886 19484 34892
rect 18696 34604 18748 34610
rect 18696 34546 18748 34552
rect 18708 33658 18736 34546
rect 18880 33856 18932 33862
rect 18880 33798 18932 33804
rect 18892 33658 18920 33798
rect 18604 33652 18656 33658
rect 18604 33594 18656 33600
rect 18696 33652 18748 33658
rect 18696 33594 18748 33600
rect 18880 33652 18932 33658
rect 18880 33594 18932 33600
rect 17868 33448 17920 33454
rect 17868 33390 17920 33396
rect 17880 32978 17908 33390
rect 17960 33380 18012 33386
rect 17960 33322 18012 33328
rect 17972 32978 18000 33322
rect 18616 33318 18644 33594
rect 19444 33590 19472 34886
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 19996 34746 20024 35022
rect 19984 34740 20036 34746
rect 19984 34682 20036 34688
rect 20732 34678 20760 36042
rect 20812 35692 20864 35698
rect 20812 35634 20864 35640
rect 20720 34672 20772 34678
rect 20720 34614 20772 34620
rect 19708 34604 19760 34610
rect 19708 34546 19760 34552
rect 19720 34202 19748 34546
rect 19708 34196 19760 34202
rect 19708 34138 19760 34144
rect 20732 34066 20760 34614
rect 20824 34134 20852 35634
rect 21008 35630 21036 36110
rect 20996 35624 21048 35630
rect 20996 35566 21048 35572
rect 21272 35556 21324 35562
rect 21272 35498 21324 35504
rect 21284 34678 21312 35498
rect 21272 34672 21324 34678
rect 21272 34614 21324 34620
rect 20996 34400 21048 34406
rect 20996 34342 21048 34348
rect 20812 34128 20864 34134
rect 20812 34070 20864 34076
rect 20720 34060 20772 34066
rect 20720 34002 20772 34008
rect 19984 33992 20036 33998
rect 19984 33934 20036 33940
rect 20260 33992 20312 33998
rect 20260 33934 20312 33940
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 19996 33590 20024 33934
rect 19340 33584 19392 33590
rect 19340 33526 19392 33532
rect 19432 33584 19484 33590
rect 19432 33526 19484 33532
rect 19984 33584 20036 33590
rect 19984 33526 20036 33532
rect 19248 33448 19300 33454
rect 19248 33390 19300 33396
rect 18604 33312 18656 33318
rect 18604 33254 18656 33260
rect 19260 33046 19288 33390
rect 19352 33114 19380 33526
rect 20272 33522 20300 33934
rect 20732 33522 20760 34002
rect 20260 33516 20312 33522
rect 20260 33458 20312 33464
rect 20720 33516 20772 33522
rect 20720 33458 20772 33464
rect 20732 33386 20760 33458
rect 20824 33454 20852 34070
rect 21008 33930 21036 34342
rect 20996 33924 21048 33930
rect 20996 33866 21048 33872
rect 21284 33522 21312 34614
rect 21272 33516 21324 33522
rect 21272 33458 21324 33464
rect 20812 33448 20864 33454
rect 20812 33390 20864 33396
rect 20720 33380 20772 33386
rect 20720 33322 20772 33328
rect 19340 33108 19392 33114
rect 19340 33050 19392 33056
rect 19248 33040 19300 33046
rect 19248 32982 19300 32988
rect 17868 32972 17920 32978
rect 17868 32914 17920 32920
rect 17960 32972 18012 32978
rect 17960 32914 18012 32920
rect 18512 32972 18564 32978
rect 18512 32914 18564 32920
rect 17880 32026 17908 32914
rect 18420 32904 18472 32910
rect 18420 32846 18472 32852
rect 18432 32434 18460 32846
rect 18144 32428 18196 32434
rect 18144 32370 18196 32376
rect 18420 32428 18472 32434
rect 18420 32370 18472 32376
rect 17868 32020 17920 32026
rect 17868 31962 17920 31968
rect 17776 31816 17828 31822
rect 17776 31758 17828 31764
rect 17500 31680 17552 31686
rect 17500 31622 17552 31628
rect 16856 30796 16908 30802
rect 16856 30738 16908 30744
rect 17316 30728 17368 30734
rect 17316 30670 17368 30676
rect 16672 30320 16724 30326
rect 16672 30262 16724 30268
rect 16764 30252 16816 30258
rect 16764 30194 16816 30200
rect 16776 29850 16804 30194
rect 17328 30122 17356 30670
rect 17316 30116 17368 30122
rect 17316 30058 17368 30064
rect 16764 29844 16816 29850
rect 16764 29786 16816 29792
rect 16488 29708 16540 29714
rect 16488 29650 16540 29656
rect 16396 29572 16448 29578
rect 16396 29514 16448 29520
rect 15200 28756 15252 28762
rect 15200 28698 15252 28704
rect 15948 28750 16252 28778
rect 14464 28212 14516 28218
rect 14464 28154 14516 28160
rect 15212 28014 15240 28698
rect 15200 28008 15252 28014
rect 15200 27950 15252 27956
rect 14280 26988 14332 26994
rect 14280 26930 14332 26936
rect 15476 26988 15528 26994
rect 15476 26930 15528 26936
rect 15488 26586 15516 26930
rect 15476 26580 15528 26586
rect 15476 26522 15528 26528
rect 15568 25968 15620 25974
rect 15568 25910 15620 25916
rect 15580 25362 15608 25910
rect 15844 25900 15896 25906
rect 15948 25888 15976 28750
rect 16408 28694 16436 29514
rect 16500 28762 16528 29650
rect 17408 29504 17460 29510
rect 17408 29446 17460 29452
rect 17040 29164 17092 29170
rect 17040 29106 17092 29112
rect 16672 29028 16724 29034
rect 16672 28970 16724 28976
rect 16488 28756 16540 28762
rect 16488 28698 16540 28704
rect 16396 28688 16448 28694
rect 16396 28630 16448 28636
rect 16580 28552 16632 28558
rect 16580 28494 16632 28500
rect 16120 28416 16172 28422
rect 16120 28358 16172 28364
rect 16028 28076 16080 28082
rect 16132 28064 16160 28358
rect 16080 28036 16160 28064
rect 16028 28018 16080 28024
rect 16132 27674 16160 28036
rect 16592 27674 16620 28494
rect 16120 27668 16172 27674
rect 16120 27610 16172 27616
rect 16580 27668 16632 27674
rect 16580 27610 16632 27616
rect 16684 27606 16712 28970
rect 16856 28620 16908 28626
rect 16856 28562 16908 28568
rect 16868 28082 16896 28562
rect 17052 28150 17080 29106
rect 17316 29096 17368 29102
rect 17316 29038 17368 29044
rect 17224 28960 17276 28966
rect 17224 28902 17276 28908
rect 17236 28626 17264 28902
rect 17328 28694 17356 29038
rect 17316 28688 17368 28694
rect 17316 28630 17368 28636
rect 17224 28620 17276 28626
rect 17224 28562 17276 28568
rect 17040 28144 17092 28150
rect 17040 28086 17092 28092
rect 16856 28076 16908 28082
rect 16856 28018 16908 28024
rect 16764 27872 16816 27878
rect 16764 27814 16816 27820
rect 16672 27600 16724 27606
rect 16672 27542 16724 27548
rect 16672 27464 16724 27470
rect 16776 27418 16804 27814
rect 16868 27470 16896 28018
rect 16724 27412 16804 27418
rect 16672 27406 16804 27412
rect 16856 27464 16908 27470
rect 16856 27406 16908 27412
rect 16684 27390 16804 27406
rect 16684 27062 16712 27390
rect 16868 27130 16896 27406
rect 16856 27124 16908 27130
rect 16856 27066 16908 27072
rect 17420 27062 17448 29446
rect 17512 28558 17540 31622
rect 17592 30320 17644 30326
rect 17592 30262 17644 30268
rect 17604 29646 17632 30262
rect 17684 30048 17736 30054
rect 17684 29990 17736 29996
rect 17696 29714 17724 29990
rect 17684 29708 17736 29714
rect 17684 29650 17736 29656
rect 17880 29646 17908 31962
rect 18156 30938 18184 32370
rect 18328 32360 18380 32366
rect 18328 32302 18380 32308
rect 18340 31958 18368 32302
rect 18328 31952 18380 31958
rect 18328 31894 18380 31900
rect 18524 31686 18552 32914
rect 19156 32836 19208 32842
rect 19156 32778 19208 32784
rect 19168 32298 19196 32778
rect 19156 32292 19208 32298
rect 19156 32234 19208 32240
rect 18972 32224 19024 32230
rect 18972 32166 19024 32172
rect 18984 31754 19012 32166
rect 19260 31822 19288 32982
rect 21180 32904 21232 32910
rect 21180 32846 21232 32852
rect 19432 32768 19484 32774
rect 19432 32710 19484 32716
rect 19444 32502 19472 32710
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 19432 32496 19484 32502
rect 19432 32438 19484 32444
rect 20628 32496 20680 32502
rect 20628 32438 20680 32444
rect 20352 32224 20404 32230
rect 20352 32166 20404 32172
rect 19248 31816 19300 31822
rect 19248 31758 19300 31764
rect 18972 31748 19024 31754
rect 18972 31690 19024 31696
rect 18512 31680 18564 31686
rect 18512 31622 18564 31628
rect 18144 30932 18196 30938
rect 18144 30874 18196 30880
rect 17960 30796 18012 30802
rect 17960 30738 18012 30744
rect 18144 30796 18196 30802
rect 18144 30738 18196 30744
rect 17592 29640 17644 29646
rect 17592 29582 17644 29588
rect 17868 29640 17920 29646
rect 17868 29582 17920 29588
rect 17972 29306 18000 30738
rect 18052 30728 18104 30734
rect 18052 30670 18104 30676
rect 18064 29850 18092 30670
rect 18052 29844 18104 29850
rect 18052 29786 18104 29792
rect 18156 29306 18184 30738
rect 18524 30734 18552 31622
rect 18604 31476 18656 31482
rect 18604 31418 18656 31424
rect 18616 30870 18644 31418
rect 18984 31278 19012 31690
rect 19156 31680 19208 31686
rect 19156 31622 19208 31628
rect 19168 31278 19196 31622
rect 19260 31414 19288 31758
rect 20364 31754 20392 32166
rect 20352 31748 20404 31754
rect 20352 31690 20404 31696
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 19248 31408 19300 31414
rect 19248 31350 19300 31356
rect 20168 31340 20220 31346
rect 20168 31282 20220 31288
rect 18972 31272 19024 31278
rect 18972 31214 19024 31220
rect 19156 31272 19208 31278
rect 19156 31214 19208 31220
rect 18604 30864 18656 30870
rect 18604 30806 18656 30812
rect 18512 30728 18564 30734
rect 18512 30670 18564 30676
rect 18236 30252 18288 30258
rect 18236 30194 18288 30200
rect 17960 29300 18012 29306
rect 17960 29242 18012 29248
rect 18144 29300 18196 29306
rect 18144 29242 18196 29248
rect 18248 29102 18276 30194
rect 18328 29640 18380 29646
rect 18328 29582 18380 29588
rect 18236 29096 18288 29102
rect 18236 29038 18288 29044
rect 18340 29034 18368 29582
rect 18420 29572 18472 29578
rect 18420 29514 18472 29520
rect 18432 29170 18460 29514
rect 18420 29164 18472 29170
rect 18420 29106 18472 29112
rect 17868 29028 17920 29034
rect 17868 28970 17920 28976
rect 18328 29028 18380 29034
rect 18328 28970 18380 28976
rect 17500 28552 17552 28558
rect 17500 28494 17552 28500
rect 17880 28218 17908 28970
rect 18328 28552 18380 28558
rect 18328 28494 18380 28500
rect 18052 28416 18104 28422
rect 18052 28358 18104 28364
rect 17868 28212 17920 28218
rect 17868 28154 17920 28160
rect 17684 28076 17736 28082
rect 17684 28018 17736 28024
rect 17696 27470 17724 28018
rect 17880 27538 17908 28154
rect 18064 28082 18092 28358
rect 18052 28076 18104 28082
rect 18052 28018 18104 28024
rect 17960 27940 18012 27946
rect 17960 27882 18012 27888
rect 17972 27674 18000 27882
rect 18340 27878 18368 28494
rect 18328 27872 18380 27878
rect 18328 27814 18380 27820
rect 17960 27668 18012 27674
rect 17960 27610 18012 27616
rect 17868 27532 17920 27538
rect 17868 27474 17920 27480
rect 17684 27464 17736 27470
rect 17684 27406 17736 27412
rect 17592 27328 17644 27334
rect 17592 27270 17644 27276
rect 16672 27056 16724 27062
rect 16672 26998 16724 27004
rect 17408 27056 17460 27062
rect 17408 26998 17460 27004
rect 16212 26784 16264 26790
rect 16212 26726 16264 26732
rect 16120 26512 16172 26518
rect 16120 26454 16172 26460
rect 15896 25860 15976 25888
rect 15844 25842 15896 25848
rect 15844 25696 15896 25702
rect 15844 25638 15896 25644
rect 15568 25356 15620 25362
rect 15568 25298 15620 25304
rect 15580 24274 15608 25298
rect 15856 25294 15884 25638
rect 15844 25288 15896 25294
rect 15844 25230 15896 25236
rect 15568 24268 15620 24274
rect 15568 24210 15620 24216
rect 15580 23202 15608 24210
rect 15752 23724 15804 23730
rect 15752 23666 15804 23672
rect 16028 23724 16080 23730
rect 16028 23666 16080 23672
rect 15488 23174 15608 23202
rect 15488 23118 15516 23174
rect 15476 23112 15528 23118
rect 15476 23054 15528 23060
rect 15488 22778 15516 23054
rect 15660 23044 15712 23050
rect 15660 22986 15712 22992
rect 15476 22772 15528 22778
rect 15476 22714 15528 22720
rect 15488 22094 15516 22714
rect 15672 22574 15700 22986
rect 15764 22642 15792 23666
rect 15936 23520 15988 23526
rect 15936 23462 15988 23468
rect 15948 22642 15976 23462
rect 15752 22636 15804 22642
rect 15752 22578 15804 22584
rect 15936 22636 15988 22642
rect 15936 22578 15988 22584
rect 15660 22568 15712 22574
rect 15660 22510 15712 22516
rect 15488 22066 15608 22094
rect 15292 22024 15344 22030
rect 15292 21966 15344 21972
rect 14740 21888 14792 21894
rect 14740 21830 14792 21836
rect 14752 20942 14780 21830
rect 14556 20936 14608 20942
rect 14556 20878 14608 20884
rect 14740 20936 14792 20942
rect 14740 20878 14792 20884
rect 14096 20460 14148 20466
rect 14096 20402 14148 20408
rect 14568 20058 14596 20878
rect 15200 20800 15252 20806
rect 15200 20742 15252 20748
rect 15212 20466 15240 20742
rect 15200 20460 15252 20466
rect 15200 20402 15252 20408
rect 14556 20052 14608 20058
rect 14556 19994 14608 20000
rect 13544 19372 13596 19378
rect 13544 19314 13596 19320
rect 13556 18970 13584 19314
rect 13544 18964 13596 18970
rect 13544 18906 13596 18912
rect 13556 15502 13584 18906
rect 14568 18698 14596 19994
rect 15304 19786 15332 21966
rect 15476 21344 15528 21350
rect 15580 21332 15608 22066
rect 15752 21956 15804 21962
rect 15752 21898 15804 21904
rect 15528 21304 15608 21332
rect 15476 21286 15528 21292
rect 15488 20534 15516 21286
rect 15764 21026 15792 21898
rect 15764 20998 15976 21026
rect 15948 20942 15976 20998
rect 15936 20936 15988 20942
rect 15936 20878 15988 20884
rect 15568 20868 15620 20874
rect 15568 20810 15620 20816
rect 15660 20868 15712 20874
rect 15660 20810 15712 20816
rect 15476 20528 15528 20534
rect 15476 20470 15528 20476
rect 15384 20460 15436 20466
rect 15384 20402 15436 20408
rect 15292 19780 15344 19786
rect 15292 19722 15344 19728
rect 15292 19440 15344 19446
rect 15396 19428 15424 20402
rect 15344 19400 15424 19428
rect 15292 19382 15344 19388
rect 15108 19372 15160 19378
rect 15160 19320 15240 19334
rect 15108 19314 15240 19320
rect 15120 19306 15240 19314
rect 15212 18766 15240 19306
rect 15292 19236 15344 19242
rect 15292 19178 15344 19184
rect 15200 18760 15252 18766
rect 15200 18702 15252 18708
rect 14556 18692 14608 18698
rect 14556 18634 14608 18640
rect 14568 18290 14596 18634
rect 14740 18624 14792 18630
rect 14740 18566 14792 18572
rect 14752 18290 14780 18566
rect 14464 18284 14516 18290
rect 14464 18226 14516 18232
rect 14556 18284 14608 18290
rect 14556 18226 14608 18232
rect 14740 18284 14792 18290
rect 14740 18226 14792 18232
rect 14476 18086 14504 18226
rect 15304 18154 15332 19178
rect 15488 18834 15516 20470
rect 15580 19990 15608 20810
rect 15568 19984 15620 19990
rect 15568 19926 15620 19932
rect 15580 19310 15608 19926
rect 15672 19446 15700 20810
rect 15844 20256 15896 20262
rect 15844 20198 15896 20204
rect 15856 19922 15884 20198
rect 15844 19916 15896 19922
rect 15844 19858 15896 19864
rect 15948 19786 15976 20878
rect 15936 19780 15988 19786
rect 15936 19722 15988 19728
rect 15660 19440 15712 19446
rect 15660 19382 15712 19388
rect 16040 19334 16068 23666
rect 16132 22642 16160 26454
rect 16224 26382 16252 26726
rect 16212 26376 16264 26382
rect 16212 26318 16264 26324
rect 16580 26240 16632 26246
rect 16580 26182 16632 26188
rect 16592 26042 16620 26182
rect 16580 26036 16632 26042
rect 16580 25978 16632 25984
rect 16684 25906 16712 26998
rect 17420 26586 17448 26998
rect 17604 26994 17632 27270
rect 17592 26988 17644 26994
rect 17592 26930 17644 26936
rect 17696 26586 17724 27406
rect 17880 27146 17908 27474
rect 17972 27470 18000 27610
rect 18340 27606 18368 27814
rect 18328 27600 18380 27606
rect 18328 27542 18380 27548
rect 17960 27464 18012 27470
rect 17960 27406 18012 27412
rect 17788 27118 17908 27146
rect 17788 26926 17816 27118
rect 17868 26988 17920 26994
rect 17868 26930 17920 26936
rect 17776 26920 17828 26926
rect 17776 26862 17828 26868
rect 17408 26580 17460 26586
rect 17408 26522 17460 26528
rect 17684 26580 17736 26586
rect 17684 26522 17736 26528
rect 17880 26450 17908 26930
rect 17868 26444 17920 26450
rect 17868 26386 17920 26392
rect 16764 26376 16816 26382
rect 16764 26318 16816 26324
rect 16672 25900 16724 25906
rect 16672 25842 16724 25848
rect 16776 25838 16804 26318
rect 17040 26308 17092 26314
rect 17040 26250 17092 26256
rect 17052 25906 17080 26250
rect 17040 25900 17092 25906
rect 17040 25842 17092 25848
rect 16764 25832 16816 25838
rect 16764 25774 16816 25780
rect 16776 25498 16804 25774
rect 16764 25492 16816 25498
rect 16764 25434 16816 25440
rect 17880 25294 17908 26386
rect 17972 26382 18000 27406
rect 18340 26382 18368 27542
rect 17960 26376 18012 26382
rect 17960 26318 18012 26324
rect 18328 26376 18380 26382
rect 18328 26318 18380 26324
rect 17972 25906 18000 26318
rect 18052 26240 18104 26246
rect 18052 26182 18104 26188
rect 17960 25900 18012 25906
rect 17960 25842 18012 25848
rect 17972 25498 18000 25842
rect 17960 25492 18012 25498
rect 17960 25434 18012 25440
rect 18064 25362 18092 26182
rect 18144 25900 18196 25906
rect 18144 25842 18196 25848
rect 18156 25498 18184 25842
rect 18144 25492 18196 25498
rect 18144 25434 18196 25440
rect 18052 25356 18104 25362
rect 18052 25298 18104 25304
rect 18616 25294 18644 30806
rect 18984 29578 19012 31214
rect 20180 30938 20208 31282
rect 20168 30932 20220 30938
rect 20168 30874 20220 30880
rect 19340 30592 19392 30598
rect 19340 30534 19392 30540
rect 20640 30546 20668 32438
rect 20720 32224 20772 32230
rect 20720 32166 20772 32172
rect 20732 30734 20760 32166
rect 21192 31822 21220 32846
rect 21284 32570 21312 33458
rect 21364 33312 21416 33318
rect 21364 33254 21416 33260
rect 21376 32774 21404 33254
rect 21364 32768 21416 32774
rect 21364 32710 21416 32716
rect 21272 32564 21324 32570
rect 21272 32506 21324 32512
rect 21180 31816 21232 31822
rect 21180 31758 21232 31764
rect 21192 31278 21220 31758
rect 21180 31272 21232 31278
rect 21180 31214 21232 31220
rect 21284 31142 21312 32506
rect 21376 32434 21404 32710
rect 21364 32428 21416 32434
rect 21364 32370 21416 32376
rect 21272 31136 21324 31142
rect 21272 31078 21324 31084
rect 21284 30870 21312 31078
rect 21272 30864 21324 30870
rect 21272 30806 21324 30812
rect 20720 30728 20772 30734
rect 20720 30670 20772 30676
rect 20904 30728 20956 30734
rect 20904 30670 20956 30676
rect 20916 30546 20944 30670
rect 19352 30326 19380 30534
rect 20640 30518 20944 30546
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19340 30320 19392 30326
rect 19340 30262 19392 30268
rect 19248 30252 19300 30258
rect 19248 30194 19300 30200
rect 19064 30184 19116 30190
rect 19064 30126 19116 30132
rect 18972 29572 19024 29578
rect 18972 29514 19024 29520
rect 18972 29300 19024 29306
rect 18972 29242 19024 29248
rect 18984 29186 19012 29242
rect 18892 29170 19012 29186
rect 19076 29170 19104 30126
rect 19260 29850 19288 30194
rect 19248 29844 19300 29850
rect 19248 29786 19300 29792
rect 19352 29238 19380 30262
rect 20444 30252 20496 30258
rect 20444 30194 20496 30200
rect 19984 29844 20036 29850
rect 19984 29786 20036 29792
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 19432 29300 19484 29306
rect 19432 29242 19484 29248
rect 19340 29232 19392 29238
rect 19340 29174 19392 29180
rect 18880 29164 19012 29170
rect 18932 29158 19012 29164
rect 19064 29164 19116 29170
rect 18880 29106 18932 29112
rect 19064 29106 19116 29112
rect 19076 28626 19104 29106
rect 19248 29096 19300 29102
rect 19248 29038 19300 29044
rect 19064 28620 19116 28626
rect 19064 28562 19116 28568
rect 19260 26382 19288 29038
rect 19444 28082 19472 29242
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 19432 28076 19484 28082
rect 19432 28018 19484 28024
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 19996 26518 20024 29786
rect 20456 29646 20484 30194
rect 20444 29640 20496 29646
rect 20444 29582 20496 29588
rect 20456 29170 20484 29582
rect 20444 29164 20496 29170
rect 20444 29106 20496 29112
rect 20168 27396 20220 27402
rect 20168 27338 20220 27344
rect 19984 26512 20036 26518
rect 19984 26454 20036 26460
rect 19248 26376 19300 26382
rect 19248 26318 19300 26324
rect 19260 25770 19288 26318
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19984 25900 20036 25906
rect 19984 25842 20036 25848
rect 19248 25764 19300 25770
rect 19248 25706 19300 25712
rect 17868 25288 17920 25294
rect 17868 25230 17920 25236
rect 18604 25288 18656 25294
rect 18604 25230 18656 25236
rect 19064 25288 19116 25294
rect 19064 25230 19116 25236
rect 18144 24268 18196 24274
rect 18144 24210 18196 24216
rect 16396 24200 16448 24206
rect 16396 24142 16448 24148
rect 16408 23662 16436 24142
rect 17960 24132 18012 24138
rect 17960 24074 18012 24080
rect 16948 24064 17000 24070
rect 16948 24006 17000 24012
rect 16396 23656 16448 23662
rect 16396 23598 16448 23604
rect 16960 23186 16988 24006
rect 17972 23866 18000 24074
rect 17960 23860 18012 23866
rect 17960 23802 18012 23808
rect 18156 23730 18184 24210
rect 18604 24200 18656 24206
rect 18604 24142 18656 24148
rect 17224 23724 17276 23730
rect 17224 23666 17276 23672
rect 18144 23724 18196 23730
rect 18144 23666 18196 23672
rect 18236 23724 18288 23730
rect 18236 23666 18288 23672
rect 17236 23322 17264 23666
rect 17224 23316 17276 23322
rect 17224 23258 17276 23264
rect 16948 23180 17000 23186
rect 16948 23122 17000 23128
rect 16120 22636 16172 22642
rect 16120 22578 16172 22584
rect 16132 22094 16160 22578
rect 16304 22568 16356 22574
rect 16304 22510 16356 22516
rect 16316 22098 16344 22510
rect 16960 22438 16988 23122
rect 17236 22642 17264 23258
rect 18052 23180 18104 23186
rect 18052 23122 18104 23128
rect 17224 22636 17276 22642
rect 17224 22578 17276 22584
rect 17776 22636 17828 22642
rect 17776 22578 17828 22584
rect 16672 22432 16724 22438
rect 16672 22374 16724 22380
rect 16948 22432 17000 22438
rect 16948 22374 17000 22380
rect 16132 22066 16252 22094
rect 15568 19304 15620 19310
rect 15568 19246 15620 19252
rect 15856 19306 16068 19334
rect 15476 18828 15528 18834
rect 15476 18770 15528 18776
rect 15292 18148 15344 18154
rect 15292 18090 15344 18096
rect 14464 18080 14516 18086
rect 14464 18022 14516 18028
rect 14476 17202 14504 18022
rect 15568 17740 15620 17746
rect 15568 17682 15620 17688
rect 15200 17604 15252 17610
rect 15200 17546 15252 17552
rect 15212 17338 15240 17546
rect 15200 17332 15252 17338
rect 15200 17274 15252 17280
rect 15580 17202 15608 17682
rect 14464 17196 14516 17202
rect 14464 17138 14516 17144
rect 15568 17196 15620 17202
rect 15568 17138 15620 17144
rect 15292 16992 15344 16998
rect 15292 16934 15344 16940
rect 15304 16658 15332 16934
rect 15752 16788 15804 16794
rect 15752 16730 15804 16736
rect 15292 16652 15344 16658
rect 15292 16594 15344 16600
rect 15304 16114 15332 16594
rect 15764 16522 15792 16730
rect 15856 16726 15884 19306
rect 16120 19304 16172 19310
rect 16120 19246 16172 19252
rect 16132 18766 16160 19246
rect 16120 18760 16172 18766
rect 16120 18702 16172 18708
rect 16028 18624 16080 18630
rect 16028 18566 16080 18572
rect 16040 18358 16068 18566
rect 16028 18352 16080 18358
rect 16028 18294 16080 18300
rect 16028 18216 16080 18222
rect 16132 18170 16160 18702
rect 16080 18164 16160 18170
rect 16028 18158 16160 18164
rect 16040 18142 16160 18158
rect 16224 17202 16252 22066
rect 16304 22092 16356 22098
rect 16304 22034 16356 22040
rect 16316 21010 16344 22034
rect 16684 22030 16712 22374
rect 16672 22024 16724 22030
rect 16672 21966 16724 21972
rect 16396 21888 16448 21894
rect 16396 21830 16448 21836
rect 16304 21004 16356 21010
rect 16304 20946 16356 20952
rect 16316 20602 16344 20946
rect 16408 20602 16436 21830
rect 16684 20942 16712 21966
rect 17788 21690 17816 22578
rect 18064 22506 18092 23122
rect 18248 23050 18276 23666
rect 18616 23662 18644 24142
rect 18604 23656 18656 23662
rect 18604 23598 18656 23604
rect 18616 23186 18644 23598
rect 18604 23180 18656 23186
rect 18604 23122 18656 23128
rect 18236 23044 18288 23050
rect 18236 22986 18288 22992
rect 18052 22500 18104 22506
rect 18052 22442 18104 22448
rect 18144 22094 18196 22098
rect 18248 22094 18276 22986
rect 18604 22432 18656 22438
rect 18604 22374 18656 22380
rect 18144 22092 18276 22094
rect 18196 22066 18276 22092
rect 18144 22034 18196 22040
rect 17776 21684 17828 21690
rect 17776 21626 17828 21632
rect 17500 21344 17552 21350
rect 17500 21286 17552 21292
rect 17512 21010 17540 21286
rect 17788 21010 17816 21626
rect 18156 21622 18184 22034
rect 18328 21956 18380 21962
rect 18328 21898 18380 21904
rect 18144 21616 18196 21622
rect 18144 21558 18196 21564
rect 18236 21548 18288 21554
rect 18236 21490 18288 21496
rect 18248 21350 18276 21490
rect 18236 21344 18288 21350
rect 18236 21286 18288 21292
rect 17500 21004 17552 21010
rect 17500 20946 17552 20952
rect 17776 21004 17828 21010
rect 17776 20946 17828 20952
rect 16672 20936 16724 20942
rect 16672 20878 16724 20884
rect 17408 20868 17460 20874
rect 17408 20810 17460 20816
rect 16304 20596 16356 20602
rect 16304 20538 16356 20544
rect 16396 20596 16448 20602
rect 16396 20538 16448 20544
rect 16408 20058 16436 20538
rect 17420 20466 17448 20810
rect 17512 20534 17540 20946
rect 18144 20800 18196 20806
rect 18144 20742 18196 20748
rect 17500 20528 17552 20534
rect 17500 20470 17552 20476
rect 17132 20460 17184 20466
rect 17132 20402 17184 20408
rect 17408 20460 17460 20466
rect 17408 20402 17460 20408
rect 16396 20052 16448 20058
rect 16396 19994 16448 20000
rect 17144 19854 17172 20402
rect 17420 20058 17448 20402
rect 17868 20392 17920 20398
rect 17868 20334 17920 20340
rect 17880 20058 17908 20334
rect 17408 20052 17460 20058
rect 17408 19994 17460 20000
rect 17868 20052 17920 20058
rect 17868 19994 17920 20000
rect 17132 19848 17184 19854
rect 17132 19790 17184 19796
rect 16948 18964 17000 18970
rect 16948 18906 17000 18912
rect 16764 18692 16816 18698
rect 16764 18634 16816 18640
rect 16776 18358 16804 18634
rect 16764 18352 16816 18358
rect 16764 18294 16816 18300
rect 16960 18290 16988 18906
rect 17144 18766 17172 19790
rect 17500 19712 17552 19718
rect 17500 19654 17552 19660
rect 17684 19712 17736 19718
rect 17684 19654 17736 19660
rect 17224 19440 17276 19446
rect 17224 19382 17276 19388
rect 17132 18760 17184 18766
rect 17132 18702 17184 18708
rect 17040 18352 17092 18358
rect 17040 18294 17092 18300
rect 16948 18284 17000 18290
rect 16948 18226 17000 18232
rect 16672 18080 16724 18086
rect 16672 18022 16724 18028
rect 16856 18080 16908 18086
rect 16960 18068 16988 18226
rect 17052 18154 17080 18294
rect 17040 18148 17092 18154
rect 17040 18090 17092 18096
rect 16908 18040 16988 18068
rect 16856 18022 16908 18028
rect 16212 17196 16264 17202
rect 16212 17138 16264 17144
rect 16684 16794 16712 18022
rect 16960 17882 16988 18040
rect 16948 17876 17000 17882
rect 16948 17818 17000 17824
rect 17052 17678 17080 18090
rect 17132 17740 17184 17746
rect 17132 17682 17184 17688
rect 17040 17672 17092 17678
rect 17040 17614 17092 17620
rect 16764 17196 16816 17202
rect 16764 17138 16816 17144
rect 16948 17196 17000 17202
rect 17052 17184 17080 17614
rect 17144 17202 17172 17682
rect 17000 17156 17080 17184
rect 17132 17196 17184 17202
rect 16948 17138 17000 17144
rect 17132 17138 17184 17144
rect 16028 16788 16080 16794
rect 16028 16730 16080 16736
rect 16672 16788 16724 16794
rect 16672 16730 16724 16736
rect 15844 16720 15896 16726
rect 15844 16662 15896 16668
rect 15752 16516 15804 16522
rect 15752 16458 15804 16464
rect 15660 16244 15712 16250
rect 15660 16186 15712 16192
rect 15292 16108 15344 16114
rect 15292 16050 15344 16056
rect 15672 16046 15700 16186
rect 15856 16046 15884 16662
rect 15936 16652 15988 16658
rect 15936 16594 15988 16600
rect 14740 16040 14792 16046
rect 14740 15982 14792 15988
rect 15660 16040 15712 16046
rect 15660 15982 15712 15988
rect 15844 16040 15896 16046
rect 15844 15982 15896 15988
rect 13544 15496 13596 15502
rect 13544 15438 13596 15444
rect 13556 15026 13584 15438
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 14280 14816 14332 14822
rect 14280 14758 14332 14764
rect 14292 14482 14320 14758
rect 14280 14476 14332 14482
rect 14280 14418 14332 14424
rect 14004 14408 14056 14414
rect 14004 14350 14056 14356
rect 14016 14074 14044 14350
rect 14004 14068 14056 14074
rect 14004 14010 14056 14016
rect 13096 6886 13308 6914
rect 12992 3596 13044 3602
rect 12992 3538 13044 3544
rect 13096 3466 13124 6886
rect 14752 6866 14780 15982
rect 15672 15706 15700 15982
rect 15660 15700 15712 15706
rect 15660 15642 15712 15648
rect 15856 15162 15884 15982
rect 15948 15706 15976 16594
rect 16040 16590 16068 16730
rect 16028 16584 16080 16590
rect 16028 16526 16080 16532
rect 16672 16584 16724 16590
rect 16776 16572 16804 17138
rect 16948 16992 17000 16998
rect 16948 16934 17000 16940
rect 16960 16590 16988 16934
rect 16724 16544 16804 16572
rect 16672 16526 16724 16532
rect 16040 16114 16068 16526
rect 16776 16182 16804 16544
rect 16948 16584 17000 16590
rect 16948 16526 17000 16532
rect 16764 16176 16816 16182
rect 16764 16118 16816 16124
rect 16028 16108 16080 16114
rect 16028 16050 16080 16056
rect 16672 16040 16724 16046
rect 16672 15982 16724 15988
rect 16580 15904 16632 15910
rect 16580 15846 16632 15852
rect 15936 15700 15988 15706
rect 15936 15642 15988 15648
rect 16592 15502 16620 15846
rect 16684 15706 16712 15982
rect 16776 15910 16804 16118
rect 17132 16108 17184 16114
rect 17052 16068 17132 16096
rect 16948 15972 17000 15978
rect 17052 15960 17080 16068
rect 17132 16050 17184 16056
rect 17000 15932 17080 15960
rect 16948 15914 17000 15920
rect 16764 15904 16816 15910
rect 16764 15846 16816 15852
rect 16672 15700 16724 15706
rect 16672 15642 16724 15648
rect 16672 15564 16724 15570
rect 16672 15506 16724 15512
rect 16580 15496 16632 15502
rect 16580 15438 16632 15444
rect 15844 15156 15896 15162
rect 15844 15098 15896 15104
rect 15936 14340 15988 14346
rect 15936 14282 15988 14288
rect 14740 6860 14792 6866
rect 14740 6802 14792 6808
rect 15476 3936 15528 3942
rect 15476 3878 15528 3884
rect 13268 3732 13320 3738
rect 13268 3674 13320 3680
rect 13084 3460 13136 3466
rect 13084 3402 13136 3408
rect 13280 3398 13308 3674
rect 15488 3602 15516 3878
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 13360 3528 13412 3534
rect 13360 3470 13412 3476
rect 13176 3392 13228 3398
rect 13176 3334 13228 3340
rect 13268 3392 13320 3398
rect 13268 3334 13320 3340
rect 13188 3126 13216 3334
rect 13176 3120 13228 3126
rect 13176 3062 13228 3068
rect 13372 3058 13400 3470
rect 15752 3460 15804 3466
rect 15752 3402 15804 3408
rect 15764 3194 15792 3402
rect 15752 3188 15804 3194
rect 15752 3130 15804 3136
rect 13360 3052 13412 3058
rect 13360 2994 13412 3000
rect 15948 2650 15976 14282
rect 16684 13938 16712 15506
rect 16672 13932 16724 13938
rect 16672 13874 16724 13880
rect 16948 13932 17000 13938
rect 16948 13874 17000 13880
rect 16684 11694 16712 13874
rect 16960 13530 16988 13874
rect 16948 13524 17000 13530
rect 16948 13466 17000 13472
rect 17236 13462 17264 19382
rect 17408 18760 17460 18766
rect 17408 18702 17460 18708
rect 17316 17808 17368 17814
rect 17316 17750 17368 17756
rect 17328 16658 17356 17750
rect 17420 17542 17448 18702
rect 17512 18698 17540 19654
rect 17696 18834 17724 19654
rect 17684 18828 17736 18834
rect 17684 18770 17736 18776
rect 17500 18692 17552 18698
rect 17500 18634 17552 18640
rect 17512 17678 17540 18634
rect 17592 18624 17644 18630
rect 17592 18566 17644 18572
rect 17604 18358 17632 18566
rect 17592 18352 17644 18358
rect 17592 18294 17644 18300
rect 17684 18284 17736 18290
rect 17684 18226 17736 18232
rect 17592 18080 17644 18086
rect 17592 18022 17644 18028
rect 17500 17672 17552 17678
rect 17500 17614 17552 17620
rect 17408 17536 17460 17542
rect 17408 17478 17460 17484
rect 17408 17332 17460 17338
rect 17408 17274 17460 17280
rect 17316 16652 17368 16658
rect 17316 16594 17368 16600
rect 17328 15638 17356 16594
rect 17420 16590 17448 17274
rect 17500 17196 17552 17202
rect 17500 17138 17552 17144
rect 17512 16794 17540 17138
rect 17500 16788 17552 16794
rect 17500 16730 17552 16736
rect 17408 16584 17460 16590
rect 17408 16526 17460 16532
rect 17420 16114 17448 16526
rect 17604 16114 17632 18022
rect 17696 16522 17724 18226
rect 17880 17746 17908 19994
rect 18156 19786 18184 20742
rect 18340 20466 18368 21898
rect 18328 20460 18380 20466
rect 18328 20402 18380 20408
rect 18144 19780 18196 19786
rect 18144 19722 18196 19728
rect 18328 19780 18380 19786
rect 18328 19722 18380 19728
rect 18052 18624 18104 18630
rect 18052 18566 18104 18572
rect 17868 17740 17920 17746
rect 17868 17682 17920 17688
rect 17880 17134 17908 17682
rect 17868 17128 17920 17134
rect 17868 17070 17920 17076
rect 17684 16516 17736 16522
rect 17684 16458 17736 16464
rect 17696 16250 17724 16458
rect 17880 16250 17908 17070
rect 18064 16454 18092 18566
rect 18156 18290 18184 19722
rect 18340 19446 18368 19722
rect 18328 19440 18380 19446
rect 18328 19382 18380 19388
rect 18616 18766 18644 22374
rect 19076 22094 19104 25230
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 19996 24954 20024 25842
rect 19984 24948 20036 24954
rect 19984 24890 20036 24896
rect 20180 24274 20208 27338
rect 20456 25362 20484 29106
rect 20916 29034 20944 30518
rect 21468 29850 21496 37742
rect 21548 36372 21600 36378
rect 21548 36314 21600 36320
rect 21560 36038 21588 36314
rect 21548 36032 21600 36038
rect 21548 35974 21600 35980
rect 21652 35766 21680 37810
rect 22008 36848 22060 36854
rect 22008 36790 22060 36796
rect 21732 36780 21784 36786
rect 21732 36722 21784 36728
rect 21744 36378 21772 36722
rect 21916 36644 21968 36650
rect 21916 36586 21968 36592
rect 21732 36372 21784 36378
rect 21732 36314 21784 36320
rect 21824 36304 21876 36310
rect 21824 36246 21876 36252
rect 21928 36258 21956 36586
rect 22020 36394 22048 36790
rect 22376 36712 22428 36718
rect 22376 36654 22428 36660
rect 22192 36576 22244 36582
rect 22192 36518 22244 36524
rect 22020 36378 22140 36394
rect 22020 36372 22152 36378
rect 22020 36366 22100 36372
rect 22100 36314 22152 36320
rect 21640 35760 21692 35766
rect 21640 35702 21692 35708
rect 21836 33930 21864 36246
rect 21928 36230 22048 36258
rect 22020 36174 22048 36230
rect 22008 36168 22060 36174
rect 22008 36110 22060 36116
rect 21916 36100 21968 36106
rect 21916 36042 21968 36048
rect 21928 35834 21956 36042
rect 21916 35828 21968 35834
rect 21916 35770 21968 35776
rect 22204 34678 22232 36518
rect 22388 36174 22416 36654
rect 22376 36168 22428 36174
rect 22376 36110 22428 36116
rect 22284 35284 22336 35290
rect 22284 35226 22336 35232
rect 22192 34672 22244 34678
rect 22192 34614 22244 34620
rect 22100 33992 22152 33998
rect 22204 33980 22232 34614
rect 22296 34474 22324 35226
rect 22284 34468 22336 34474
rect 22284 34410 22336 34416
rect 22296 33998 22324 34410
rect 22388 34134 22416 36110
rect 22376 34128 22428 34134
rect 22376 34070 22428 34076
rect 22152 33952 22232 33980
rect 22284 33992 22336 33998
rect 22100 33934 22152 33940
rect 22284 33934 22336 33940
rect 22376 33992 22428 33998
rect 22376 33934 22428 33940
rect 21824 33924 21876 33930
rect 21824 33866 21876 33872
rect 21836 33386 21864 33866
rect 22192 33856 22244 33862
rect 22192 33798 22244 33804
rect 22204 33454 22232 33798
rect 22388 33590 22416 33934
rect 22376 33584 22428 33590
rect 22376 33526 22428 33532
rect 22468 33516 22520 33522
rect 22468 33458 22520 33464
rect 22192 33448 22244 33454
rect 22192 33390 22244 33396
rect 21824 33380 21876 33386
rect 21824 33322 21876 33328
rect 22100 32224 22152 32230
rect 22100 32166 22152 32172
rect 21824 31272 21876 31278
rect 21824 31214 21876 31220
rect 21456 29844 21508 29850
rect 21456 29786 21508 29792
rect 21272 29232 21324 29238
rect 21272 29174 21324 29180
rect 20536 29028 20588 29034
rect 20536 28970 20588 28976
rect 20904 29028 20956 29034
rect 20904 28970 20956 28976
rect 20444 25356 20496 25362
rect 20444 25298 20496 25304
rect 20352 25152 20404 25158
rect 20352 25094 20404 25100
rect 20364 24818 20392 25094
rect 20352 24812 20404 24818
rect 20352 24754 20404 24760
rect 20456 24274 20484 25298
rect 20168 24268 20220 24274
rect 20168 24210 20220 24216
rect 20444 24268 20496 24274
rect 20444 24210 20496 24216
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 19432 23860 19484 23866
rect 19432 23802 19484 23808
rect 19156 23724 19208 23730
rect 19156 23666 19208 23672
rect 19168 22778 19196 23666
rect 19444 23254 19472 23802
rect 20456 23798 20484 24210
rect 19708 23792 19760 23798
rect 19708 23734 19760 23740
rect 20444 23792 20496 23798
rect 20444 23734 20496 23740
rect 19432 23248 19484 23254
rect 19432 23190 19484 23196
rect 19720 23118 19748 23734
rect 20076 23724 20128 23730
rect 20076 23666 20128 23672
rect 19984 23520 20036 23526
rect 19984 23462 20036 23468
rect 19340 23112 19392 23118
rect 19340 23054 19392 23060
rect 19708 23112 19760 23118
rect 19708 23054 19760 23060
rect 19248 22976 19300 22982
rect 19248 22918 19300 22924
rect 19156 22772 19208 22778
rect 19156 22714 19208 22720
rect 19260 22642 19288 22918
rect 19248 22636 19300 22642
rect 19248 22578 19300 22584
rect 19352 22098 19380 23054
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19432 22704 19484 22710
rect 19432 22646 19484 22652
rect 19076 22066 19196 22094
rect 18972 21956 19024 21962
rect 18972 21898 19024 21904
rect 18984 21554 19012 21898
rect 18972 21548 19024 21554
rect 18972 21490 19024 21496
rect 19064 21548 19116 21554
rect 19064 21490 19116 21496
rect 18696 20596 18748 20602
rect 18696 20538 18748 20544
rect 18708 19378 18736 20538
rect 19076 20534 19104 21490
rect 19064 20528 19116 20534
rect 19064 20470 19116 20476
rect 19076 19718 19104 20470
rect 19168 20466 19196 22066
rect 19340 22092 19392 22098
rect 19340 22034 19392 22040
rect 19340 21956 19392 21962
rect 19340 21898 19392 21904
rect 19248 21888 19300 21894
rect 19248 21830 19300 21836
rect 19260 21622 19288 21830
rect 19248 21616 19300 21622
rect 19248 21558 19300 21564
rect 19352 20602 19380 21898
rect 19444 21690 19472 22646
rect 19996 22030 20024 23462
rect 20088 23118 20116 23666
rect 20444 23180 20496 23186
rect 20444 23122 20496 23128
rect 20076 23112 20128 23118
rect 20076 23054 20128 23060
rect 20088 22438 20116 23054
rect 20352 23044 20404 23050
rect 20352 22986 20404 22992
rect 20076 22432 20128 22438
rect 20076 22374 20128 22380
rect 19984 22024 20036 22030
rect 19984 21966 20036 21972
rect 20260 22024 20312 22030
rect 20260 21966 20312 21972
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19432 21684 19484 21690
rect 19432 21626 19484 21632
rect 19444 21010 19472 21626
rect 20272 21554 20300 21966
rect 20076 21548 20128 21554
rect 20076 21490 20128 21496
rect 20260 21548 20312 21554
rect 20260 21490 20312 21496
rect 19524 21480 19576 21486
rect 19524 21422 19576 21428
rect 19432 21004 19484 21010
rect 19432 20946 19484 20952
rect 19536 20890 19564 21422
rect 19444 20862 19564 20890
rect 19984 20868 20036 20874
rect 19340 20596 19392 20602
rect 19340 20538 19392 20544
rect 19156 20460 19208 20466
rect 19156 20402 19208 20408
rect 19340 20460 19392 20466
rect 19340 20402 19392 20408
rect 19352 20058 19380 20402
rect 19340 20052 19392 20058
rect 19340 19994 19392 20000
rect 19064 19712 19116 19718
rect 19064 19654 19116 19660
rect 19444 19378 19472 20862
rect 19984 20810 20036 20816
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19996 20602 20024 20810
rect 19984 20596 20036 20602
rect 19984 20538 20036 20544
rect 19984 20460 20036 20466
rect 19984 20402 20036 20408
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 18696 19372 18748 19378
rect 18696 19314 18748 19320
rect 19432 19372 19484 19378
rect 19432 19314 19484 19320
rect 19340 19168 19392 19174
rect 19340 19110 19392 19116
rect 19352 18970 19380 19110
rect 19340 18964 19392 18970
rect 19340 18906 19392 18912
rect 18328 18760 18380 18766
rect 18328 18702 18380 18708
rect 18604 18760 18656 18766
rect 18604 18702 18656 18708
rect 18144 18284 18196 18290
rect 18144 18226 18196 18232
rect 18340 18222 18368 18702
rect 19432 18692 19484 18698
rect 19432 18634 19484 18640
rect 19444 18358 19472 18634
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19432 18352 19484 18358
rect 19432 18294 19484 18300
rect 18696 18284 18748 18290
rect 18696 18226 18748 18232
rect 18328 18216 18380 18222
rect 18328 18158 18380 18164
rect 18708 16454 18736 18226
rect 19444 18222 19472 18294
rect 19432 18216 19484 18222
rect 19432 18158 19484 18164
rect 19432 18080 19484 18086
rect 19432 18022 19484 18028
rect 19444 17678 19472 18022
rect 19432 17672 19484 17678
rect 19432 17614 19484 17620
rect 19432 17536 19484 17542
rect 19432 17478 19484 17484
rect 19444 17202 19472 17478
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 19432 17196 19484 17202
rect 19432 17138 19484 17144
rect 19616 17196 19668 17202
rect 19616 17138 19668 17144
rect 19524 17128 19576 17134
rect 19524 17070 19576 17076
rect 19536 16658 19564 17070
rect 19524 16652 19576 16658
rect 19524 16594 19576 16600
rect 19248 16584 19300 16590
rect 19248 16526 19300 16532
rect 19260 16454 19288 16526
rect 19628 16522 19656 17138
rect 19616 16516 19668 16522
rect 19616 16458 19668 16464
rect 18052 16448 18104 16454
rect 18052 16390 18104 16396
rect 18696 16448 18748 16454
rect 18696 16390 18748 16396
rect 19248 16448 19300 16454
rect 19248 16390 19300 16396
rect 17684 16244 17736 16250
rect 17684 16186 17736 16192
rect 17868 16244 17920 16250
rect 17868 16186 17920 16192
rect 17408 16108 17460 16114
rect 17408 16050 17460 16056
rect 17592 16108 17644 16114
rect 17592 16050 17644 16056
rect 18512 16108 18564 16114
rect 18512 16050 18564 16056
rect 17316 15632 17368 15638
rect 17316 15574 17368 15580
rect 17604 15502 17632 16050
rect 17592 15496 17644 15502
rect 17592 15438 17644 15444
rect 18144 15156 18196 15162
rect 18144 15098 18196 15104
rect 18052 14816 18104 14822
rect 18052 14758 18104 14764
rect 18064 14414 18092 14758
rect 18052 14408 18104 14414
rect 18052 14350 18104 14356
rect 18156 14346 18184 15098
rect 18524 15026 18552 16050
rect 19260 15502 19288 16390
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 19340 15972 19392 15978
rect 19340 15914 19392 15920
rect 19248 15496 19300 15502
rect 19248 15438 19300 15444
rect 19248 15360 19300 15366
rect 19248 15302 19300 15308
rect 19064 15088 19116 15094
rect 19064 15030 19116 15036
rect 18512 15020 18564 15026
rect 18512 14962 18564 14968
rect 18524 14618 18552 14962
rect 18788 14952 18840 14958
rect 18788 14894 18840 14900
rect 18512 14612 18564 14618
rect 18512 14554 18564 14560
rect 18800 14482 18828 14894
rect 18788 14476 18840 14482
rect 18788 14418 18840 14424
rect 18328 14408 18380 14414
rect 18328 14350 18380 14356
rect 18144 14340 18196 14346
rect 18144 14282 18196 14288
rect 17960 14068 18012 14074
rect 17960 14010 18012 14016
rect 17224 13456 17276 13462
rect 17224 13398 17276 13404
rect 17236 12434 17264 13398
rect 17972 13326 18000 14010
rect 18052 14000 18104 14006
rect 18052 13942 18104 13948
rect 18064 13530 18092 13942
rect 18052 13524 18104 13530
rect 18052 13466 18104 13472
rect 17960 13320 18012 13326
rect 17960 13262 18012 13268
rect 18156 12986 18184 14282
rect 18340 13870 18368 14350
rect 18328 13864 18380 13870
rect 18328 13806 18380 13812
rect 18800 13530 18828 14418
rect 19076 14006 19104 15030
rect 19260 14822 19288 15302
rect 19248 14816 19300 14822
rect 19248 14758 19300 14764
rect 19064 14000 19116 14006
rect 19064 13942 19116 13948
rect 19076 13870 19104 13942
rect 19064 13864 19116 13870
rect 19064 13806 19116 13812
rect 18788 13524 18840 13530
rect 18788 13466 18840 13472
rect 19076 13462 19104 13806
rect 19260 13734 19288 14758
rect 19352 14414 19380 15914
rect 19996 15706 20024 20402
rect 20088 20058 20116 21490
rect 20364 21418 20392 22986
rect 20456 22506 20484 23122
rect 20444 22500 20496 22506
rect 20444 22442 20496 22448
rect 20352 21412 20404 21418
rect 20352 21354 20404 21360
rect 20260 20460 20312 20466
rect 20364 20448 20392 21354
rect 20456 21350 20484 22442
rect 20444 21344 20496 21350
rect 20444 21286 20496 21292
rect 20456 20890 20484 21286
rect 20548 21026 20576 28970
rect 21284 28762 21312 29174
rect 21732 29164 21784 29170
rect 21732 29106 21784 29112
rect 21272 28756 21324 28762
rect 21272 28698 21324 28704
rect 20720 28484 20772 28490
rect 20720 28426 20772 28432
rect 20732 27606 20760 28426
rect 21284 28218 21312 28698
rect 21640 28416 21692 28422
rect 21640 28358 21692 28364
rect 21272 28212 21324 28218
rect 21272 28154 21324 28160
rect 20904 27872 20956 27878
rect 20904 27814 20956 27820
rect 20720 27600 20772 27606
rect 20626 27568 20682 27577
rect 20720 27542 20772 27548
rect 20626 27503 20682 27512
rect 20640 27402 20668 27503
rect 20916 27470 20944 27814
rect 21284 27538 21312 28154
rect 21272 27532 21324 27538
rect 21272 27474 21324 27480
rect 21652 27470 21680 28358
rect 21744 27606 21772 29106
rect 21836 29102 21864 31214
rect 22112 30326 22140 32166
rect 22204 31958 22232 33390
rect 22376 33312 22428 33318
rect 22376 33254 22428 33260
rect 22388 32434 22416 33254
rect 22376 32428 22428 32434
rect 22376 32370 22428 32376
rect 22284 32360 22336 32366
rect 22284 32302 22336 32308
rect 22296 32230 22324 32302
rect 22284 32224 22336 32230
rect 22284 32166 22336 32172
rect 22192 31952 22244 31958
rect 22192 31894 22244 31900
rect 22204 31822 22232 31894
rect 22480 31822 22508 33458
rect 22192 31816 22244 31822
rect 22468 31816 22520 31822
rect 22192 31758 22244 31764
rect 22296 31776 22468 31804
rect 22296 31482 22324 31776
rect 22468 31758 22520 31764
rect 22284 31476 22336 31482
rect 22284 31418 22336 31424
rect 22284 31340 22336 31346
rect 22284 31282 22336 31288
rect 22296 30938 22324 31282
rect 22284 30932 22336 30938
rect 22284 30874 22336 30880
rect 22100 30320 22152 30326
rect 22100 30262 22152 30268
rect 21824 29096 21876 29102
rect 21824 29038 21876 29044
rect 21836 28558 21864 29038
rect 22192 28756 22244 28762
rect 22192 28698 22244 28704
rect 21824 28552 21876 28558
rect 21824 28494 21876 28500
rect 21916 28416 21968 28422
rect 21916 28358 21968 28364
rect 21928 28150 21956 28358
rect 22204 28218 22232 28698
rect 22284 28552 22336 28558
rect 22284 28494 22336 28500
rect 22192 28212 22244 28218
rect 22192 28154 22244 28160
rect 21916 28144 21968 28150
rect 21916 28086 21968 28092
rect 22296 28082 22324 28494
rect 22284 28076 22336 28082
rect 22284 28018 22336 28024
rect 22296 27674 22324 28018
rect 22284 27668 22336 27674
rect 22284 27610 22336 27616
rect 21732 27600 21784 27606
rect 21732 27542 21784 27548
rect 20904 27464 20956 27470
rect 20904 27406 20956 27412
rect 21640 27464 21692 27470
rect 21640 27406 21692 27412
rect 20628 27396 20680 27402
rect 20628 27338 20680 27344
rect 22376 26512 22428 26518
rect 22376 26454 22428 26460
rect 22100 26376 22152 26382
rect 22100 26318 22152 26324
rect 22284 26376 22336 26382
rect 22284 26318 22336 26324
rect 20812 26240 20864 26246
rect 20812 26182 20864 26188
rect 20996 26240 21048 26246
rect 20996 26182 21048 26188
rect 21272 26240 21324 26246
rect 21272 26182 21324 26188
rect 20824 25294 20852 26182
rect 21008 25702 21036 26182
rect 20996 25696 21048 25702
rect 20996 25638 21048 25644
rect 21008 25294 21036 25638
rect 21284 25498 21312 26182
rect 22112 25498 22140 26318
rect 22192 26240 22244 26246
rect 22192 26182 22244 26188
rect 22204 25906 22232 26182
rect 22192 25900 22244 25906
rect 22192 25842 22244 25848
rect 21272 25492 21324 25498
rect 21272 25434 21324 25440
rect 22100 25492 22152 25498
rect 22100 25434 22152 25440
rect 20812 25288 20864 25294
rect 20812 25230 20864 25236
rect 20996 25288 21048 25294
rect 20996 25230 21048 25236
rect 22296 24750 22324 26318
rect 22388 25226 22416 26454
rect 22376 25220 22428 25226
rect 22376 25162 22428 25168
rect 22388 24818 22416 25162
rect 22376 24812 22428 24818
rect 22376 24754 22428 24760
rect 22284 24744 22336 24750
rect 22284 24686 22336 24692
rect 22376 24200 22428 24206
rect 22376 24142 22428 24148
rect 22388 23798 22416 24142
rect 22376 23792 22428 23798
rect 22376 23734 22428 23740
rect 22100 23588 22152 23594
rect 22100 23530 22152 23536
rect 21272 23520 21324 23526
rect 21272 23462 21324 23468
rect 21284 23118 21312 23462
rect 21272 23112 21324 23118
rect 21272 23054 21324 23060
rect 21456 22976 21508 22982
rect 21456 22918 21508 22924
rect 20812 22636 20864 22642
rect 20812 22578 20864 22584
rect 20628 22432 20680 22438
rect 20628 22374 20680 22380
rect 20640 21486 20668 22374
rect 20824 21554 20852 22578
rect 20904 22432 20956 22438
rect 20904 22374 20956 22380
rect 20916 22030 20944 22374
rect 21468 22030 21496 22918
rect 20904 22024 20956 22030
rect 20904 21966 20956 21972
rect 21456 22024 21508 22030
rect 21456 21966 21508 21972
rect 20812 21548 20864 21554
rect 20812 21490 20864 21496
rect 21468 21486 21496 21966
rect 20628 21480 20680 21486
rect 20628 21422 20680 21428
rect 21456 21480 21508 21486
rect 21456 21422 21508 21428
rect 20548 20998 20668 21026
rect 21468 21010 21496 21422
rect 22112 21418 22140 23530
rect 22468 22636 22520 22642
rect 22468 22578 22520 22584
rect 22480 21622 22508 22578
rect 22572 22094 22600 41550
rect 22848 40934 22876 41550
rect 24412 41414 24440 41550
rect 24136 41386 24440 41414
rect 22836 40928 22888 40934
rect 22836 40870 22888 40876
rect 23388 40928 23440 40934
rect 23388 40870 23440 40876
rect 22928 39432 22980 39438
rect 22928 39374 22980 39380
rect 22940 38758 22968 39374
rect 22928 38752 22980 38758
rect 22928 38694 22980 38700
rect 22940 38214 22968 38694
rect 23020 38344 23072 38350
rect 23020 38286 23072 38292
rect 22928 38208 22980 38214
rect 22928 38150 22980 38156
rect 22652 36168 22704 36174
rect 22652 36110 22704 36116
rect 22664 35290 22692 36110
rect 22744 35828 22796 35834
rect 22744 35770 22796 35776
rect 22756 35494 22784 35770
rect 22744 35488 22796 35494
rect 22744 35430 22796 35436
rect 22652 35284 22704 35290
rect 22652 35226 22704 35232
rect 22756 35154 22784 35430
rect 22836 35284 22888 35290
rect 22836 35226 22888 35232
rect 22744 35148 22796 35154
rect 22744 35090 22796 35096
rect 22652 35080 22704 35086
rect 22652 35022 22704 35028
rect 22664 34746 22692 35022
rect 22652 34740 22704 34746
rect 22652 34682 22704 34688
rect 22756 34678 22784 35090
rect 22848 34746 22876 35226
rect 22836 34740 22888 34746
rect 22836 34682 22888 34688
rect 22744 34672 22796 34678
rect 22744 34614 22796 34620
rect 22836 34604 22888 34610
rect 22836 34546 22888 34552
rect 22848 34202 22876 34546
rect 22836 34196 22888 34202
rect 22836 34138 22888 34144
rect 22744 33448 22796 33454
rect 22744 33390 22796 33396
rect 22756 32502 22784 33390
rect 22836 32836 22888 32842
rect 22836 32778 22888 32784
rect 22848 32570 22876 32778
rect 22836 32564 22888 32570
rect 22836 32506 22888 32512
rect 22744 32496 22796 32502
rect 22744 32438 22796 32444
rect 22756 31754 22784 32438
rect 22744 31748 22796 31754
rect 22744 31690 22796 31696
rect 22756 30802 22784 31690
rect 22744 30796 22796 30802
rect 22744 30738 22796 30744
rect 22652 28620 22704 28626
rect 22652 28562 22704 28568
rect 22664 28082 22692 28562
rect 22744 28144 22796 28150
rect 22744 28086 22796 28092
rect 22652 28076 22704 28082
rect 22652 28018 22704 28024
rect 22664 27334 22692 28018
rect 22756 27606 22784 28086
rect 22744 27600 22796 27606
rect 22744 27542 22796 27548
rect 22652 27328 22704 27334
rect 22652 27270 22704 27276
rect 22940 26382 22968 38150
rect 23032 35154 23060 38286
rect 23204 37868 23256 37874
rect 23204 37810 23256 37816
rect 23216 37466 23244 37810
rect 23204 37460 23256 37466
rect 23204 37402 23256 37408
rect 23400 35834 23428 40870
rect 24136 40497 24164 41386
rect 24122 40488 24178 40497
rect 24122 40423 24178 40432
rect 26424 40452 26476 40458
rect 23756 36848 23808 36854
rect 23756 36790 23808 36796
rect 23664 36780 23716 36786
rect 23664 36722 23716 36728
rect 23480 36168 23532 36174
rect 23480 36110 23532 36116
rect 23388 35828 23440 35834
rect 23388 35770 23440 35776
rect 23492 35290 23520 36110
rect 23676 35766 23704 36722
rect 23664 35760 23716 35766
rect 23664 35702 23716 35708
rect 23676 35290 23704 35702
rect 23480 35284 23532 35290
rect 23480 35226 23532 35232
rect 23664 35284 23716 35290
rect 23664 35226 23716 35232
rect 23020 35148 23072 35154
rect 23020 35090 23072 35096
rect 23032 35034 23060 35090
rect 23032 35018 23152 35034
rect 23032 35012 23164 35018
rect 23032 35006 23112 35012
rect 23112 34954 23164 34960
rect 23020 34740 23072 34746
rect 23020 34682 23072 34688
rect 23032 34610 23060 34682
rect 23020 34604 23072 34610
rect 23020 34546 23072 34552
rect 23204 34604 23256 34610
rect 23204 34546 23256 34552
rect 23388 34604 23440 34610
rect 23388 34546 23440 34552
rect 23216 33454 23244 34546
rect 23400 34202 23428 34546
rect 23388 34196 23440 34202
rect 23388 34138 23440 34144
rect 23296 34128 23348 34134
rect 23296 34070 23348 34076
rect 23308 33590 23336 34070
rect 23296 33584 23348 33590
rect 23296 33526 23348 33532
rect 23204 33448 23256 33454
rect 23204 33390 23256 33396
rect 23308 32450 23336 33526
rect 23664 33516 23716 33522
rect 23664 33458 23716 33464
rect 23676 33114 23704 33458
rect 23664 33108 23716 33114
rect 23664 33050 23716 33056
rect 23216 32434 23336 32450
rect 23204 32428 23336 32434
rect 23256 32422 23336 32428
rect 23204 32370 23256 32376
rect 23296 32360 23348 32366
rect 23296 32302 23348 32308
rect 23308 31754 23336 32302
rect 23388 31816 23440 31822
rect 23388 31758 23440 31764
rect 23296 31748 23348 31754
rect 23296 31690 23348 31696
rect 23112 31680 23164 31686
rect 23112 31622 23164 31628
rect 23124 30734 23152 31622
rect 23400 31482 23428 31758
rect 23388 31476 23440 31482
rect 23388 31418 23440 31424
rect 23768 30938 23796 36790
rect 23848 36032 23900 36038
rect 23848 35974 23900 35980
rect 23860 35766 23888 35974
rect 23848 35760 23900 35766
rect 23848 35702 23900 35708
rect 23848 34944 23900 34950
rect 23848 34886 23900 34892
rect 23860 34746 23888 34886
rect 23848 34740 23900 34746
rect 23848 34682 23900 34688
rect 24032 34604 24084 34610
rect 24032 34546 24084 34552
rect 24044 34066 24072 34546
rect 24032 34060 24084 34066
rect 24032 34002 24084 34008
rect 23848 32768 23900 32774
rect 23848 32710 23900 32716
rect 23756 30932 23808 30938
rect 23756 30874 23808 30880
rect 23860 30870 23888 32710
rect 23848 30864 23900 30870
rect 23848 30806 23900 30812
rect 23112 30728 23164 30734
rect 23112 30670 23164 30676
rect 23204 28960 23256 28966
rect 23204 28902 23256 28908
rect 23020 28552 23072 28558
rect 23020 28494 23072 28500
rect 23032 27674 23060 28494
rect 23216 28218 23244 28902
rect 23296 28552 23348 28558
rect 23296 28494 23348 28500
rect 23204 28212 23256 28218
rect 23204 28154 23256 28160
rect 23020 27668 23072 27674
rect 23020 27610 23072 27616
rect 23112 27464 23164 27470
rect 23112 27406 23164 27412
rect 23020 26784 23072 26790
rect 23020 26726 23072 26732
rect 22928 26376 22980 26382
rect 22928 26318 22980 26324
rect 23032 26314 23060 26726
rect 23020 26308 23072 26314
rect 23020 26250 23072 26256
rect 23032 25430 23060 26250
rect 23020 25424 23072 25430
rect 23020 25366 23072 25372
rect 23124 25158 23152 27406
rect 23216 27402 23244 28154
rect 23308 27470 23336 28494
rect 23388 28416 23440 28422
rect 23388 28358 23440 28364
rect 23400 28082 23428 28358
rect 23388 28076 23440 28082
rect 23388 28018 23440 28024
rect 23296 27464 23348 27470
rect 23296 27406 23348 27412
rect 23388 27464 23440 27470
rect 23388 27406 23440 27412
rect 23204 27396 23256 27402
rect 23204 27338 23256 27344
rect 23112 25152 23164 25158
rect 23112 25094 23164 25100
rect 23216 24614 23244 27338
rect 23400 27334 23428 27406
rect 23388 27328 23440 27334
rect 23388 27270 23440 27276
rect 23296 26988 23348 26994
rect 23296 26930 23348 26936
rect 23308 25770 23336 26930
rect 23400 26382 23428 27270
rect 24032 27056 24084 27062
rect 24032 26998 24084 27004
rect 23480 26920 23532 26926
rect 23480 26862 23532 26868
rect 23388 26376 23440 26382
rect 23388 26318 23440 26324
rect 23296 25764 23348 25770
rect 23296 25706 23348 25712
rect 23308 24818 23336 25706
rect 23400 25294 23428 26318
rect 23492 26246 23520 26862
rect 23756 26512 23808 26518
rect 23756 26454 23808 26460
rect 23480 26240 23532 26246
rect 23480 26182 23532 26188
rect 23664 25900 23716 25906
rect 23664 25842 23716 25848
rect 23572 25696 23624 25702
rect 23572 25638 23624 25644
rect 23584 25362 23612 25638
rect 23572 25356 23624 25362
rect 23572 25298 23624 25304
rect 23388 25288 23440 25294
rect 23388 25230 23440 25236
rect 23296 24812 23348 24818
rect 23296 24754 23348 24760
rect 23204 24608 23256 24614
rect 23204 24550 23256 24556
rect 23480 24132 23532 24138
rect 23480 24074 23532 24080
rect 23492 23322 23520 24074
rect 23572 24064 23624 24070
rect 23572 24006 23624 24012
rect 23584 23866 23612 24006
rect 23572 23860 23624 23866
rect 23572 23802 23624 23808
rect 23676 23730 23704 25842
rect 23768 24206 23796 26454
rect 24044 25974 24072 26998
rect 24032 25968 24084 25974
rect 24032 25910 24084 25916
rect 24044 24750 24072 25910
rect 24032 24744 24084 24750
rect 24032 24686 24084 24692
rect 23756 24200 23808 24206
rect 23756 24142 23808 24148
rect 23664 23724 23716 23730
rect 23584 23684 23664 23712
rect 23480 23316 23532 23322
rect 23480 23258 23532 23264
rect 23584 23050 23612 23684
rect 23664 23666 23716 23672
rect 23768 23322 23796 24142
rect 24044 24138 24072 24686
rect 24032 24132 24084 24138
rect 24032 24074 24084 24080
rect 23756 23316 23808 23322
rect 23756 23258 23808 23264
rect 23848 23180 23900 23186
rect 23848 23122 23900 23128
rect 23572 23044 23624 23050
rect 23572 22986 23624 22992
rect 23296 22976 23348 22982
rect 23296 22918 23348 22924
rect 22572 22066 22784 22094
rect 22284 21616 22336 21622
rect 22284 21558 22336 21564
rect 22468 21616 22520 21622
rect 22468 21558 22520 21564
rect 22100 21412 22152 21418
rect 22100 21354 22152 21360
rect 21732 21344 21784 21350
rect 21732 21286 21784 21292
rect 20456 20862 20576 20890
rect 20444 20800 20496 20806
rect 20444 20742 20496 20748
rect 20456 20466 20484 20742
rect 20312 20420 20392 20448
rect 20444 20460 20496 20466
rect 20260 20402 20312 20408
rect 20444 20402 20496 20408
rect 20076 20052 20128 20058
rect 20076 19994 20128 20000
rect 20088 19854 20116 19994
rect 20076 19848 20128 19854
rect 20076 19790 20128 19796
rect 20260 19712 20312 19718
rect 20260 19654 20312 19660
rect 20352 19712 20404 19718
rect 20352 19654 20404 19660
rect 20076 19372 20128 19378
rect 20076 19314 20128 19320
rect 20088 17202 20116 19314
rect 20272 19242 20300 19654
rect 20364 19378 20392 19654
rect 20352 19372 20404 19378
rect 20352 19314 20404 19320
rect 20548 19258 20576 20862
rect 20260 19236 20312 19242
rect 20260 19178 20312 19184
rect 20364 19230 20576 19258
rect 20364 17678 20392 19230
rect 20352 17672 20404 17678
rect 20352 17614 20404 17620
rect 20076 17196 20128 17202
rect 20076 17138 20128 17144
rect 20364 17134 20392 17614
rect 20640 17338 20668 20998
rect 21456 21004 21508 21010
rect 21456 20946 21508 20952
rect 21744 20942 21772 21286
rect 21732 20936 21784 20942
rect 21732 20878 21784 20884
rect 22008 20460 22060 20466
rect 21928 20420 22008 20448
rect 20904 20392 20956 20398
rect 20904 20334 20956 20340
rect 20916 19854 20944 20334
rect 21824 20052 21876 20058
rect 21824 19994 21876 20000
rect 21180 19984 21232 19990
rect 21180 19926 21232 19932
rect 20904 19848 20956 19854
rect 20904 19790 20956 19796
rect 20916 19514 20944 19790
rect 20904 19508 20956 19514
rect 20904 19450 20956 19456
rect 21088 19236 21140 19242
rect 21088 19178 21140 19184
rect 21100 18290 21128 19178
rect 21192 19174 21220 19926
rect 21640 19712 21692 19718
rect 21640 19654 21692 19660
rect 21548 19372 21600 19378
rect 21548 19314 21600 19320
rect 21180 19168 21232 19174
rect 21180 19110 21232 19116
rect 21560 18834 21588 19314
rect 21548 18828 21600 18834
rect 21548 18770 21600 18776
rect 21560 18290 21588 18770
rect 21088 18284 21140 18290
rect 21088 18226 21140 18232
rect 21548 18284 21600 18290
rect 21548 18226 21600 18232
rect 20628 17332 20680 17338
rect 20628 17274 20680 17280
rect 20536 17196 20588 17202
rect 20536 17138 20588 17144
rect 20352 17128 20404 17134
rect 20352 17070 20404 17076
rect 20260 16992 20312 16998
rect 20260 16934 20312 16940
rect 20272 16114 20300 16934
rect 20260 16108 20312 16114
rect 20260 16050 20312 16056
rect 19984 15700 20036 15706
rect 19984 15642 20036 15648
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 19996 15026 20024 15642
rect 20548 15502 20576 17138
rect 21180 17060 21232 17066
rect 21180 17002 21232 17008
rect 20812 16720 20864 16726
rect 20812 16662 20864 16668
rect 20824 16114 20852 16662
rect 20996 16652 21048 16658
rect 20996 16594 21048 16600
rect 20812 16108 20864 16114
rect 20812 16050 20864 16056
rect 20824 15706 20852 16050
rect 21008 15978 21036 16594
rect 21088 16448 21140 16454
rect 21088 16390 21140 16396
rect 21100 15978 21128 16390
rect 20996 15972 21048 15978
rect 20996 15914 21048 15920
rect 21088 15972 21140 15978
rect 21088 15914 21140 15920
rect 20812 15700 20864 15706
rect 20812 15642 20864 15648
rect 21100 15570 21128 15914
rect 21192 15706 21220 17002
rect 21560 16182 21588 18226
rect 21652 16590 21680 19654
rect 21836 18834 21864 19994
rect 21824 18828 21876 18834
rect 21824 18770 21876 18776
rect 21824 17196 21876 17202
rect 21824 17138 21876 17144
rect 21640 16584 21692 16590
rect 21640 16526 21692 16532
rect 21548 16176 21600 16182
rect 21548 16118 21600 16124
rect 21180 15700 21232 15706
rect 21180 15642 21232 15648
rect 21560 15570 21588 16118
rect 21640 15904 21692 15910
rect 21640 15846 21692 15852
rect 21088 15564 21140 15570
rect 21088 15506 21140 15512
rect 21548 15564 21600 15570
rect 21548 15506 21600 15512
rect 20536 15496 20588 15502
rect 20536 15438 20588 15444
rect 21180 15088 21232 15094
rect 21180 15030 21232 15036
rect 19984 15020 20036 15026
rect 19984 14962 20036 14968
rect 20904 15020 20956 15026
rect 20956 14980 21036 15008
rect 20904 14962 20956 14968
rect 19432 14816 19484 14822
rect 19432 14758 19484 14764
rect 19708 14816 19760 14822
rect 19708 14758 19760 14764
rect 19340 14408 19392 14414
rect 19340 14350 19392 14356
rect 19248 13728 19300 13734
rect 19248 13670 19300 13676
rect 19064 13456 19116 13462
rect 19064 13398 19116 13404
rect 18420 13388 18472 13394
rect 18420 13330 18472 13336
rect 18144 12980 18196 12986
rect 18144 12922 18196 12928
rect 18432 12442 18460 13330
rect 19260 13326 19288 13670
rect 19248 13320 19300 13326
rect 19248 13262 19300 13268
rect 18512 13252 18564 13258
rect 18512 13194 18564 13200
rect 18524 12850 18552 13194
rect 18696 12912 18748 12918
rect 18696 12854 18748 12860
rect 18512 12844 18564 12850
rect 18512 12786 18564 12792
rect 18708 12782 18736 12854
rect 18696 12776 18748 12782
rect 18696 12718 18748 12724
rect 17144 12406 17264 12434
rect 18420 12436 18472 12442
rect 16672 11688 16724 11694
rect 16672 11630 16724 11636
rect 17144 11218 17172 12406
rect 18420 12378 18472 12384
rect 17868 12232 17920 12238
rect 17868 12174 17920 12180
rect 17500 11756 17552 11762
rect 17500 11698 17552 11704
rect 17132 11212 17184 11218
rect 17132 11154 17184 11160
rect 17512 10538 17540 11698
rect 17684 11552 17736 11558
rect 17684 11494 17736 11500
rect 17696 11218 17724 11494
rect 17684 11212 17736 11218
rect 17684 11154 17736 11160
rect 17592 11008 17644 11014
rect 17592 10950 17644 10956
rect 17604 10742 17632 10950
rect 17592 10736 17644 10742
rect 17592 10678 17644 10684
rect 17500 10532 17552 10538
rect 17500 10474 17552 10480
rect 17696 10266 17724 11154
rect 17880 11150 17908 12174
rect 18328 12164 18380 12170
rect 18328 12106 18380 12112
rect 18236 11280 18288 11286
rect 18236 11222 18288 11228
rect 17776 11144 17828 11150
rect 17776 11086 17828 11092
rect 17868 11144 17920 11150
rect 17868 11086 17920 11092
rect 17788 11014 17816 11086
rect 17776 11008 17828 11014
rect 17776 10950 17828 10956
rect 17788 10674 17816 10950
rect 17880 10810 17908 11086
rect 17868 10804 17920 10810
rect 17868 10746 17920 10752
rect 17776 10668 17828 10674
rect 17776 10610 17828 10616
rect 17684 10260 17736 10266
rect 17684 10202 17736 10208
rect 17684 9988 17736 9994
rect 17684 9930 17736 9936
rect 17696 9722 17724 9930
rect 17684 9716 17736 9722
rect 17684 9658 17736 9664
rect 17788 9586 17816 10610
rect 17776 9580 17828 9586
rect 17776 9522 17828 9528
rect 18248 9518 18276 11222
rect 18340 11082 18368 12106
rect 18604 12096 18656 12102
rect 18604 12038 18656 12044
rect 18512 11620 18564 11626
rect 18512 11562 18564 11568
rect 18524 11354 18552 11562
rect 18512 11348 18564 11354
rect 18512 11290 18564 11296
rect 18616 11234 18644 12038
rect 18708 11354 18736 12718
rect 19064 11688 19116 11694
rect 19064 11630 19116 11636
rect 18696 11348 18748 11354
rect 18696 11290 18748 11296
rect 18616 11206 18736 11234
rect 18328 11076 18380 11082
rect 18328 11018 18380 11024
rect 18420 10668 18472 10674
rect 18420 10610 18472 10616
rect 18432 9586 18460 10610
rect 18708 10606 18736 11206
rect 19076 11150 19104 11630
rect 19352 11218 19380 14350
rect 19444 13938 19472 14758
rect 19720 14414 19748 14758
rect 19708 14408 19760 14414
rect 19708 14350 19760 14356
rect 20720 14272 20772 14278
rect 20720 14214 20772 14220
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19432 13932 19484 13938
rect 19432 13874 19484 13880
rect 19444 12986 19472 13874
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 20732 12918 20760 14214
rect 21008 13326 21036 14980
rect 21088 14816 21140 14822
rect 21088 14758 21140 14764
rect 20904 13320 20956 13326
rect 20904 13262 20956 13268
rect 20996 13320 21048 13326
rect 20996 13262 21048 13268
rect 20916 12918 20944 13262
rect 20720 12912 20772 12918
rect 20720 12854 20772 12860
rect 20904 12912 20956 12918
rect 20904 12854 20956 12860
rect 19892 12844 19944 12850
rect 19892 12786 19944 12792
rect 19904 12306 19932 12786
rect 20916 12594 20944 12854
rect 20732 12566 20944 12594
rect 19892 12300 19944 12306
rect 19892 12242 19944 12248
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 20260 11824 20312 11830
rect 20260 11766 20312 11772
rect 19616 11552 19668 11558
rect 19616 11494 19668 11500
rect 19432 11280 19484 11286
rect 19432 11222 19484 11228
rect 19340 11212 19392 11218
rect 19340 11154 19392 11160
rect 19064 11144 19116 11150
rect 19064 11086 19116 11092
rect 19076 10742 19104 11086
rect 19064 10736 19116 10742
rect 19064 10678 19116 10684
rect 18696 10600 18748 10606
rect 18696 10542 18748 10548
rect 18708 10266 18736 10542
rect 18696 10260 18748 10266
rect 18696 10202 18748 10208
rect 18708 9586 18736 10202
rect 19352 9586 19380 11154
rect 19444 10130 19472 11222
rect 19628 11150 19656 11494
rect 19616 11144 19668 11150
rect 19616 11086 19668 11092
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 20272 10810 20300 11766
rect 20732 11558 20760 12566
rect 21008 12434 21036 13262
rect 21100 12646 21128 14758
rect 21192 14074 21220 15030
rect 21652 14278 21680 15846
rect 21836 15638 21864 17138
rect 21824 15632 21876 15638
rect 21824 15574 21876 15580
rect 21640 14272 21692 14278
rect 21640 14214 21692 14220
rect 21180 14068 21232 14074
rect 21180 14010 21232 14016
rect 21836 14006 21864 15574
rect 21928 14346 21956 20420
rect 22008 20402 22060 20408
rect 22112 20330 22140 21354
rect 22192 20528 22244 20534
rect 22192 20470 22244 20476
rect 22100 20324 22152 20330
rect 22100 20266 22152 20272
rect 22204 19446 22232 20470
rect 22296 20058 22324 21558
rect 22376 21548 22428 21554
rect 22376 21490 22428 21496
rect 22284 20052 22336 20058
rect 22284 19994 22336 20000
rect 22192 19440 22244 19446
rect 22192 19382 22244 19388
rect 22008 16992 22060 16998
rect 22008 16934 22060 16940
rect 22020 16114 22048 16934
rect 22204 16522 22232 19382
rect 22192 16516 22244 16522
rect 22192 16458 22244 16464
rect 22388 16250 22416 21490
rect 22756 20058 22784 22066
rect 22928 21888 22980 21894
rect 22928 21830 22980 21836
rect 22940 20942 22968 21830
rect 23308 21146 23336 22918
rect 23584 22710 23612 22986
rect 23572 22704 23624 22710
rect 23624 22652 23704 22658
rect 23572 22646 23704 22652
rect 23584 22630 23704 22646
rect 23572 22568 23624 22574
rect 23572 22510 23624 22516
rect 23296 21140 23348 21146
rect 23296 21082 23348 21088
rect 22928 20936 22980 20942
rect 22928 20878 22980 20884
rect 23296 20868 23348 20874
rect 23296 20810 23348 20816
rect 22836 20256 22888 20262
rect 22836 20198 22888 20204
rect 22744 20052 22796 20058
rect 22744 19994 22796 20000
rect 22848 19854 22876 20198
rect 22836 19848 22888 19854
rect 22836 19790 22888 19796
rect 23020 19712 23072 19718
rect 23020 19654 23072 19660
rect 23032 19446 23060 19654
rect 23020 19440 23072 19446
rect 23020 19382 23072 19388
rect 23112 19304 23164 19310
rect 23112 19246 23164 19252
rect 23020 19168 23072 19174
rect 23020 19110 23072 19116
rect 23032 18766 23060 19110
rect 23020 18760 23072 18766
rect 23020 18702 23072 18708
rect 23124 18290 23152 19246
rect 23112 18284 23164 18290
rect 23112 18226 23164 18232
rect 23308 17882 23336 20810
rect 23388 20800 23440 20806
rect 23388 20742 23440 20748
rect 23400 20330 23428 20742
rect 23480 20392 23532 20398
rect 23480 20334 23532 20340
rect 23388 20324 23440 20330
rect 23388 20266 23440 20272
rect 23492 19378 23520 20334
rect 23480 19372 23532 19378
rect 23480 19314 23532 19320
rect 23492 18358 23520 19314
rect 23584 18442 23612 22510
rect 23676 21486 23704 22630
rect 23664 21480 23716 21486
rect 23664 21422 23716 21428
rect 23860 18902 23888 23122
rect 24044 23118 24072 24074
rect 24032 23112 24084 23118
rect 24032 23054 24084 23060
rect 24136 22094 24164 40423
rect 26424 40394 26476 40400
rect 24584 40044 24636 40050
rect 24584 39986 24636 39992
rect 24308 39840 24360 39846
rect 24308 39782 24360 39788
rect 24320 36922 24348 39782
rect 24596 39642 24624 39986
rect 25320 39840 25372 39846
rect 25320 39782 25372 39788
rect 24584 39636 24636 39642
rect 24584 39578 24636 39584
rect 24492 39364 24544 39370
rect 24492 39306 24544 39312
rect 24504 39098 24532 39306
rect 24492 39092 24544 39098
rect 24492 39034 24544 39040
rect 25332 38962 25360 39782
rect 26436 39506 26464 40394
rect 27068 40044 27120 40050
rect 27068 39986 27120 39992
rect 26976 39976 27028 39982
rect 26976 39918 27028 39924
rect 26424 39500 26476 39506
rect 26424 39442 26476 39448
rect 26988 39438 27016 39918
rect 27080 39642 27108 39986
rect 27068 39636 27120 39642
rect 27068 39578 27120 39584
rect 25504 39432 25556 39438
rect 25504 39374 25556 39380
rect 25596 39432 25648 39438
rect 25596 39374 25648 39380
rect 26884 39432 26936 39438
rect 26884 39374 26936 39380
rect 26976 39432 27028 39438
rect 26976 39374 27028 39380
rect 25412 39364 25464 39370
rect 25412 39306 25464 39312
rect 25424 39030 25452 39306
rect 25412 39024 25464 39030
rect 25412 38966 25464 38972
rect 24400 38956 24452 38962
rect 24400 38898 24452 38904
rect 25320 38956 25372 38962
rect 25320 38898 25372 38904
rect 24412 37806 24440 38898
rect 25044 38752 25096 38758
rect 25044 38694 25096 38700
rect 24768 38276 24820 38282
rect 24768 38218 24820 38224
rect 24400 37800 24452 37806
rect 24400 37742 24452 37748
rect 24676 37800 24728 37806
rect 24676 37742 24728 37748
rect 24688 37262 24716 37742
rect 24780 37262 24808 38218
rect 24952 38208 25004 38214
rect 24952 38150 25004 38156
rect 24860 37664 24912 37670
rect 24860 37606 24912 37612
rect 24872 37330 24900 37606
rect 24964 37330 24992 38150
rect 25056 37670 25084 38694
rect 25332 38418 25360 38898
rect 25320 38412 25372 38418
rect 25320 38354 25372 38360
rect 25044 37664 25096 37670
rect 25044 37606 25096 37612
rect 25056 37398 25084 37606
rect 25228 37460 25280 37466
rect 25228 37402 25280 37408
rect 25044 37392 25096 37398
rect 25044 37334 25096 37340
rect 24860 37324 24912 37330
rect 24860 37266 24912 37272
rect 24952 37324 25004 37330
rect 24952 37266 25004 37272
rect 24676 37256 24728 37262
rect 24676 37198 24728 37204
rect 24768 37256 24820 37262
rect 24768 37198 24820 37204
rect 24308 36916 24360 36922
rect 24308 36858 24360 36864
rect 24320 35698 24348 36858
rect 24688 36718 24716 37198
rect 25044 36780 25096 36786
rect 25044 36722 25096 36728
rect 24676 36712 24728 36718
rect 24676 36654 24728 36660
rect 25056 35698 25084 36722
rect 24308 35692 24360 35698
rect 24308 35634 24360 35640
rect 25044 35692 25096 35698
rect 25044 35634 25096 35640
rect 24320 34610 24348 35634
rect 24860 35080 24912 35086
rect 24860 35022 24912 35028
rect 24492 35012 24544 35018
rect 24492 34954 24544 34960
rect 24308 34604 24360 34610
rect 24308 34546 24360 34552
rect 24504 33590 24532 34954
rect 24872 34202 24900 35022
rect 25136 35012 25188 35018
rect 25136 34954 25188 34960
rect 24952 34944 25004 34950
rect 24952 34886 25004 34892
rect 24964 34678 24992 34886
rect 24952 34672 25004 34678
rect 24952 34614 25004 34620
rect 24860 34196 24912 34202
rect 24860 34138 24912 34144
rect 25148 33998 25176 34954
rect 25136 33992 25188 33998
rect 25136 33934 25188 33940
rect 24492 33584 24544 33590
rect 24492 33526 24544 33532
rect 24504 32502 24532 33526
rect 24768 33380 24820 33386
rect 24768 33322 24820 33328
rect 24492 32496 24544 32502
rect 24492 32438 24544 32444
rect 24676 32428 24728 32434
rect 24676 32370 24728 32376
rect 24216 32292 24268 32298
rect 24216 32234 24268 32240
rect 24228 31890 24256 32234
rect 24688 32026 24716 32370
rect 24676 32020 24728 32026
rect 24676 31962 24728 31968
rect 24216 31884 24268 31890
rect 24216 31826 24268 31832
rect 24228 31414 24256 31826
rect 24216 31408 24268 31414
rect 24216 31350 24268 31356
rect 24780 30802 24808 33322
rect 24952 32836 25004 32842
rect 24952 32778 25004 32784
rect 24964 32570 24992 32778
rect 24952 32564 25004 32570
rect 24952 32506 25004 32512
rect 25136 32360 25188 32366
rect 25136 32302 25188 32308
rect 25148 32026 25176 32302
rect 25136 32020 25188 32026
rect 25136 31962 25188 31968
rect 25044 31816 25096 31822
rect 25044 31758 25096 31764
rect 24768 30796 24820 30802
rect 24768 30738 24820 30744
rect 24308 30660 24360 30666
rect 24308 30602 24360 30608
rect 24320 30258 24348 30602
rect 24780 30258 24808 30738
rect 24308 30252 24360 30258
rect 24308 30194 24360 30200
rect 24768 30252 24820 30258
rect 24768 30194 24820 30200
rect 24860 30116 24912 30122
rect 24860 30058 24912 30064
rect 24676 30048 24728 30054
rect 24676 29990 24728 29996
rect 24688 29850 24716 29990
rect 24676 29844 24728 29850
rect 24676 29786 24728 29792
rect 24584 29232 24636 29238
rect 24584 29174 24636 29180
rect 24216 29028 24268 29034
rect 24216 28970 24268 28976
rect 24228 28626 24256 28970
rect 24216 28620 24268 28626
rect 24216 28562 24268 28568
rect 24228 28218 24256 28562
rect 24216 28212 24268 28218
rect 24216 28154 24268 28160
rect 24596 27470 24624 29174
rect 24872 29034 24900 30058
rect 24860 29028 24912 29034
rect 24860 28970 24912 28976
rect 24872 28626 24900 28970
rect 24860 28620 24912 28626
rect 24860 28562 24912 28568
rect 24860 27940 24912 27946
rect 24860 27882 24912 27888
rect 24584 27464 24636 27470
rect 24584 27406 24636 27412
rect 24492 26376 24544 26382
rect 24492 26318 24544 26324
rect 24504 26246 24532 26318
rect 24492 26240 24544 26246
rect 24492 26182 24544 26188
rect 24504 25974 24532 26182
rect 24492 25968 24544 25974
rect 24492 25910 24544 25916
rect 24504 25498 24532 25910
rect 24492 25492 24544 25498
rect 24492 25434 24544 25440
rect 24504 24682 24532 25434
rect 24492 24676 24544 24682
rect 24492 24618 24544 24624
rect 24584 23180 24636 23186
rect 24584 23122 24636 23128
rect 24400 23112 24452 23118
rect 24400 23054 24452 23060
rect 24412 22642 24440 23054
rect 24596 22982 24624 23122
rect 24872 23118 24900 27882
rect 24952 25288 25004 25294
rect 24952 25230 25004 25236
rect 24964 24818 24992 25230
rect 24952 24812 25004 24818
rect 24952 24754 25004 24760
rect 25056 23322 25084 31758
rect 25240 31482 25268 37402
rect 25424 31754 25452 38966
rect 25516 38214 25544 39374
rect 25608 39030 25636 39374
rect 26896 39098 26924 39374
rect 26884 39092 26936 39098
rect 26884 39034 26936 39040
rect 25596 39024 25648 39030
rect 25596 38966 25648 38972
rect 27172 38962 27200 43046
rect 27816 42226 27844 43046
rect 27804 42220 27856 42226
rect 27804 42162 27856 42168
rect 28368 42158 28396 45200
rect 30472 43104 30524 43110
rect 30472 43046 30524 43052
rect 30484 42770 30512 43046
rect 30944 42770 30972 45200
rect 33520 43246 33548 45200
rect 33324 43240 33376 43246
rect 33324 43182 33376 43188
rect 33508 43240 33560 43246
rect 33508 43182 33560 43188
rect 33140 43172 33192 43178
rect 33140 43114 33192 43120
rect 33152 42770 33180 43114
rect 30472 42764 30524 42770
rect 30472 42706 30524 42712
rect 30932 42764 30984 42770
rect 30932 42706 30984 42712
rect 33140 42764 33192 42770
rect 33140 42706 33192 42712
rect 30656 42628 30708 42634
rect 30656 42570 30708 42576
rect 30668 42362 30696 42570
rect 33336 42362 33364 43182
rect 33968 42696 34020 42702
rect 33968 42638 34020 42644
rect 33416 42560 33468 42566
rect 33416 42502 33468 42508
rect 30656 42356 30708 42362
rect 30656 42298 30708 42304
rect 33324 42356 33376 42362
rect 33324 42298 33376 42304
rect 33428 42226 33456 42502
rect 33980 42226 34008 42638
rect 34164 42362 34192 45200
rect 34520 43104 34572 43110
rect 34520 43046 34572 43052
rect 34152 42356 34204 42362
rect 34152 42298 34204 42304
rect 30564 42220 30616 42226
rect 30564 42162 30616 42168
rect 33416 42220 33468 42226
rect 33416 42162 33468 42168
rect 33968 42220 34020 42226
rect 33968 42162 34020 42168
rect 28080 42152 28132 42158
rect 28080 42094 28132 42100
rect 28356 42152 28408 42158
rect 28356 42094 28408 42100
rect 28092 41818 28120 42094
rect 28080 41812 28132 41818
rect 28080 41754 28132 41760
rect 30576 41750 30604 42162
rect 30564 41744 30616 41750
rect 30564 41686 30616 41692
rect 28172 41608 28224 41614
rect 28172 41550 28224 41556
rect 28080 40384 28132 40390
rect 28080 40326 28132 40332
rect 27436 40180 27488 40186
rect 27436 40122 27488 40128
rect 27448 39506 27476 40122
rect 27436 39500 27488 39506
rect 27436 39442 27488 39448
rect 25872 38956 25924 38962
rect 25872 38898 25924 38904
rect 27160 38956 27212 38962
rect 27160 38898 27212 38904
rect 25884 38350 25912 38898
rect 25872 38344 25924 38350
rect 25872 38286 25924 38292
rect 25504 38208 25556 38214
rect 25504 38150 25556 38156
rect 25504 37868 25556 37874
rect 25556 37828 25636 37856
rect 25504 37810 25556 37816
rect 25608 37466 25636 37828
rect 25596 37460 25648 37466
rect 25596 37402 25648 37408
rect 25608 36038 25636 37402
rect 25884 37194 25912 38286
rect 27172 38282 27200 38898
rect 27448 38894 27476 39442
rect 27896 39364 27948 39370
rect 27896 39306 27948 39312
rect 27908 39098 27936 39306
rect 27896 39092 27948 39098
rect 27896 39034 27948 39040
rect 28092 38962 28120 40326
rect 28184 39030 28212 41550
rect 30576 41002 30604 41686
rect 34532 41614 34560 43046
rect 34934 43004 35242 43024
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42928 35242 42948
rect 35440 42696 35492 42702
rect 35440 42638 35492 42644
rect 34888 42356 34940 42362
rect 34888 42298 34940 42304
rect 34900 42158 34928 42298
rect 34796 42152 34848 42158
rect 34796 42094 34848 42100
rect 34888 42152 34940 42158
rect 34888 42094 34940 42100
rect 34808 41818 34836 42094
rect 35348 42084 35400 42090
rect 35348 42026 35400 42032
rect 34934 41916 35242 41936
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41840 35242 41860
rect 34796 41812 34848 41818
rect 34796 41754 34848 41760
rect 35256 41676 35308 41682
rect 35360 41664 35388 42026
rect 35452 41682 35480 42638
rect 35624 42016 35676 42022
rect 35624 41958 35676 41964
rect 35636 41682 35664 41958
rect 36096 41682 36124 45200
rect 37384 42770 37412 45200
rect 37372 42764 37424 42770
rect 37372 42706 37424 42712
rect 37832 42628 37884 42634
rect 37832 42570 37884 42576
rect 36452 42220 36504 42226
rect 36452 42162 36504 42168
rect 35308 41636 35388 41664
rect 35440 41676 35492 41682
rect 35256 41618 35308 41624
rect 35440 41618 35492 41624
rect 35624 41676 35676 41682
rect 35624 41618 35676 41624
rect 36084 41676 36136 41682
rect 36084 41618 36136 41624
rect 34520 41608 34572 41614
rect 34520 41550 34572 41556
rect 32496 41132 32548 41138
rect 32496 41074 32548 41080
rect 32588 41132 32640 41138
rect 32588 41074 32640 41080
rect 33048 41132 33100 41138
rect 33048 41074 33100 41080
rect 33416 41132 33468 41138
rect 33416 41074 33468 41080
rect 30564 40996 30616 41002
rect 30564 40938 30616 40944
rect 32508 40730 32536 41074
rect 32312 40724 32364 40730
rect 32312 40666 32364 40672
rect 32496 40724 32548 40730
rect 32496 40666 32548 40672
rect 28908 40588 28960 40594
rect 28908 40530 28960 40536
rect 28920 39642 28948 40530
rect 31116 40520 31168 40526
rect 31116 40462 31168 40468
rect 32128 40520 32180 40526
rect 32128 40462 32180 40468
rect 30748 40452 30800 40458
rect 30748 40394 30800 40400
rect 29828 40112 29880 40118
rect 29828 40054 29880 40060
rect 28908 39636 28960 39642
rect 28908 39578 28960 39584
rect 28172 39024 28224 39030
rect 28172 38966 28224 38972
rect 28080 38956 28132 38962
rect 28080 38898 28132 38904
rect 27436 38888 27488 38894
rect 27436 38830 27488 38836
rect 26240 38276 26292 38282
rect 26240 38218 26292 38224
rect 27160 38276 27212 38282
rect 27160 38218 27212 38224
rect 26148 38208 26200 38214
rect 26148 38150 26200 38156
rect 25872 37188 25924 37194
rect 25872 37130 25924 37136
rect 26056 36712 26108 36718
rect 26160 36700 26188 38150
rect 26252 37874 26280 38218
rect 26240 37868 26292 37874
rect 26240 37810 26292 37816
rect 26108 36672 26188 36700
rect 26056 36654 26108 36660
rect 26068 36106 26096 36654
rect 26148 36576 26200 36582
rect 26148 36518 26200 36524
rect 26160 36174 26188 36518
rect 26252 36378 26280 37810
rect 27448 37738 27476 38830
rect 27804 38820 27856 38826
rect 27804 38762 27856 38768
rect 27816 37874 27844 38762
rect 27988 38208 28040 38214
rect 27988 38150 28040 38156
rect 28816 38208 28868 38214
rect 28816 38150 28868 38156
rect 27804 37868 27856 37874
rect 27804 37810 27856 37816
rect 27712 37800 27764 37806
rect 27712 37742 27764 37748
rect 27436 37732 27488 37738
rect 27436 37674 27488 37680
rect 26332 37664 26384 37670
rect 26332 37606 26384 37612
rect 26344 36786 26372 37606
rect 27448 37398 27476 37674
rect 27528 37664 27580 37670
rect 27528 37606 27580 37612
rect 27436 37392 27488 37398
rect 27436 37334 27488 37340
rect 27540 37330 27568 37606
rect 27528 37324 27580 37330
rect 27528 37266 27580 37272
rect 27528 37188 27580 37194
rect 27528 37130 27580 37136
rect 27252 37120 27304 37126
rect 27252 37062 27304 37068
rect 26332 36780 26384 36786
rect 26332 36722 26384 36728
rect 26424 36780 26476 36786
rect 26424 36722 26476 36728
rect 26332 36644 26384 36650
rect 26332 36586 26384 36592
rect 26240 36372 26292 36378
rect 26240 36314 26292 36320
rect 26344 36310 26372 36586
rect 26332 36304 26384 36310
rect 26332 36246 26384 36252
rect 26344 36174 26372 36246
rect 26148 36168 26200 36174
rect 26148 36110 26200 36116
rect 26332 36168 26384 36174
rect 26332 36110 26384 36116
rect 26056 36100 26108 36106
rect 26056 36042 26108 36048
rect 25596 36032 25648 36038
rect 25596 35974 25648 35980
rect 25608 35086 25636 35974
rect 25688 35692 25740 35698
rect 25688 35634 25740 35640
rect 25596 35080 25648 35086
rect 25596 35022 25648 35028
rect 25700 33998 25728 35634
rect 25964 35080 26016 35086
rect 25964 35022 26016 35028
rect 26344 35034 26372 36110
rect 26436 35222 26464 36722
rect 27264 36378 27292 37062
rect 27436 36576 27488 36582
rect 27436 36518 27488 36524
rect 27252 36372 27304 36378
rect 27252 36314 27304 36320
rect 27448 36212 27476 36518
rect 27540 36310 27568 37130
rect 27620 37120 27672 37126
rect 27620 37062 27672 37068
rect 27528 36304 27580 36310
rect 27528 36246 27580 36252
rect 27436 36206 27488 36212
rect 27436 36148 27488 36154
rect 27436 36032 27488 36038
rect 27436 35974 27488 35980
rect 27160 35692 27212 35698
rect 27160 35634 27212 35640
rect 26424 35216 26476 35222
rect 26424 35158 26476 35164
rect 26792 35148 26844 35154
rect 26792 35090 26844 35096
rect 25872 34740 25924 34746
rect 25872 34682 25924 34688
rect 25780 34604 25832 34610
rect 25780 34546 25832 34552
rect 25504 33992 25556 33998
rect 25504 33934 25556 33940
rect 25688 33992 25740 33998
rect 25688 33934 25740 33940
rect 25332 31726 25452 31754
rect 25228 31476 25280 31482
rect 25228 31418 25280 31424
rect 25240 30938 25268 31418
rect 25332 31142 25360 31726
rect 25320 31136 25372 31142
rect 25318 31104 25320 31113
rect 25372 31104 25374 31113
rect 25318 31039 25374 31048
rect 25228 30932 25280 30938
rect 25228 30874 25280 30880
rect 25412 30592 25464 30598
rect 25412 30534 25464 30540
rect 25228 30252 25280 30258
rect 25228 30194 25280 30200
rect 25240 29578 25268 30194
rect 25424 30054 25452 30534
rect 25412 30048 25464 30054
rect 25412 29990 25464 29996
rect 25228 29572 25280 29578
rect 25228 29514 25280 29520
rect 25240 29186 25268 29514
rect 25320 29232 25372 29238
rect 25240 29180 25320 29186
rect 25240 29174 25372 29180
rect 25240 29158 25360 29174
rect 25136 27328 25188 27334
rect 25136 27270 25188 27276
rect 25148 25226 25176 27270
rect 25136 25220 25188 25226
rect 25136 25162 25188 25168
rect 25044 23316 25096 23322
rect 25044 23258 25096 23264
rect 24860 23112 24912 23118
rect 24860 23054 24912 23060
rect 24584 22976 24636 22982
rect 24584 22918 24636 22924
rect 24596 22778 24624 22918
rect 24584 22772 24636 22778
rect 24584 22714 24636 22720
rect 25240 22710 25268 29158
rect 25412 28960 25464 28966
rect 25412 28902 25464 28908
rect 25424 28694 25452 28902
rect 25412 28688 25464 28694
rect 25412 28630 25464 28636
rect 25320 27872 25372 27878
rect 25320 27814 25372 27820
rect 25332 27402 25360 27814
rect 25320 27396 25372 27402
rect 25320 27338 25372 27344
rect 25516 26382 25544 33934
rect 25700 33454 25728 33934
rect 25688 33448 25740 33454
rect 25688 33390 25740 33396
rect 25792 33386 25820 34546
rect 25884 33998 25912 34682
rect 25872 33992 25924 33998
rect 25872 33934 25924 33940
rect 25976 33522 26004 35022
rect 26344 35006 26556 35034
rect 26148 34944 26200 34950
rect 26148 34886 26200 34892
rect 25964 33516 26016 33522
rect 25964 33458 26016 33464
rect 25780 33380 25832 33386
rect 25780 33322 25832 33328
rect 25688 32904 25740 32910
rect 25688 32846 25740 32852
rect 25700 31890 25728 32846
rect 25688 31884 25740 31890
rect 25688 31826 25740 31832
rect 25700 31210 25728 31826
rect 25976 31754 26004 33458
rect 26056 33448 26108 33454
rect 26056 33390 26108 33396
rect 26068 33114 26096 33390
rect 26056 33108 26108 33114
rect 26056 33050 26108 33056
rect 26068 32366 26096 33050
rect 26056 32360 26108 32366
rect 26056 32302 26108 32308
rect 26160 31754 26188 34886
rect 26332 32428 26384 32434
rect 26332 32370 26384 32376
rect 25964 31748 26016 31754
rect 25964 31690 26016 31696
rect 26148 31748 26200 31754
rect 26148 31690 26200 31696
rect 26344 31464 26372 32370
rect 26424 32224 26476 32230
rect 26424 32166 26476 32172
rect 26436 31822 26464 32166
rect 26424 31816 26476 31822
rect 26424 31758 26476 31764
rect 26344 31436 26464 31464
rect 25780 31408 25832 31414
rect 25780 31350 25832 31356
rect 25688 31204 25740 31210
rect 25688 31146 25740 31152
rect 25596 30660 25648 30666
rect 25596 30602 25648 30608
rect 25608 30122 25636 30602
rect 25700 30190 25728 31146
rect 25792 30734 25820 31350
rect 25872 31340 25924 31346
rect 25872 31282 25924 31288
rect 26332 31340 26384 31346
rect 26332 31282 26384 31288
rect 25780 30728 25832 30734
rect 25780 30670 25832 30676
rect 25792 30326 25820 30670
rect 25780 30320 25832 30326
rect 25780 30262 25832 30268
rect 25688 30184 25740 30190
rect 25884 30138 25912 31282
rect 25964 31136 26016 31142
rect 25964 31078 26016 31084
rect 25688 30126 25740 30132
rect 25596 30116 25648 30122
rect 25596 30058 25648 30064
rect 25700 29646 25728 30126
rect 25792 30110 25912 30138
rect 25688 29640 25740 29646
rect 25688 29582 25740 29588
rect 25700 28150 25728 29582
rect 25792 28694 25820 30110
rect 25976 29646 26004 31078
rect 26344 30394 26372 31282
rect 26436 31210 26464 31436
rect 26424 31204 26476 31210
rect 26424 31146 26476 31152
rect 26424 30660 26476 30666
rect 26424 30602 26476 30608
rect 26332 30388 26384 30394
rect 26332 30330 26384 30336
rect 26056 30048 26108 30054
rect 26056 29990 26108 29996
rect 25964 29640 26016 29646
rect 25964 29582 26016 29588
rect 25780 28688 25832 28694
rect 25780 28630 25832 28636
rect 25688 28144 25740 28150
rect 25688 28086 25740 28092
rect 25700 27538 25728 28086
rect 25688 27532 25740 27538
rect 25688 27474 25740 27480
rect 25504 26376 25556 26382
rect 25504 26318 25556 26324
rect 25412 25356 25464 25362
rect 25412 25298 25464 25304
rect 25424 24750 25452 25298
rect 25412 24744 25464 24750
rect 25412 24686 25464 24692
rect 25424 24206 25452 24686
rect 25412 24200 25464 24206
rect 25412 24142 25464 24148
rect 25228 22704 25280 22710
rect 25228 22646 25280 22652
rect 24400 22636 24452 22642
rect 24400 22578 24452 22584
rect 24136 22066 24256 22094
rect 23848 18896 23900 18902
rect 23848 18838 23900 18844
rect 23584 18414 23704 18442
rect 23480 18352 23532 18358
rect 23480 18294 23532 18300
rect 23572 18284 23624 18290
rect 23572 18226 23624 18232
rect 23584 18170 23612 18226
rect 23492 18142 23612 18170
rect 23296 17876 23348 17882
rect 23296 17818 23348 17824
rect 23308 17338 23336 17818
rect 23492 17678 23520 18142
rect 23480 17672 23532 17678
rect 23480 17614 23532 17620
rect 23296 17332 23348 17338
rect 23296 17274 23348 17280
rect 22744 17196 22796 17202
rect 22744 17138 22796 17144
rect 22756 16726 22784 17138
rect 23492 17134 23520 17614
rect 23296 17128 23348 17134
rect 23296 17070 23348 17076
rect 23480 17128 23532 17134
rect 23480 17070 23532 17076
rect 23112 16788 23164 16794
rect 23112 16730 23164 16736
rect 22744 16720 22796 16726
rect 22744 16662 22796 16668
rect 22376 16244 22428 16250
rect 22376 16186 22428 16192
rect 22008 16108 22060 16114
rect 22008 16050 22060 16056
rect 22560 15904 22612 15910
rect 22560 15846 22612 15852
rect 22572 15706 22600 15846
rect 22756 15706 22784 16662
rect 22192 15700 22244 15706
rect 22192 15642 22244 15648
rect 22560 15700 22612 15706
rect 22560 15642 22612 15648
rect 22744 15700 22796 15706
rect 22744 15642 22796 15648
rect 22204 15026 22232 15642
rect 22284 15496 22336 15502
rect 22284 15438 22336 15444
rect 22192 15020 22244 15026
rect 22192 14962 22244 14968
rect 22008 14612 22060 14618
rect 22008 14554 22060 14560
rect 22020 14482 22048 14554
rect 22204 14550 22232 14962
rect 22192 14544 22244 14550
rect 22192 14486 22244 14492
rect 22008 14476 22060 14482
rect 22008 14418 22060 14424
rect 21916 14340 21968 14346
rect 21916 14282 21968 14288
rect 21824 14000 21876 14006
rect 21824 13942 21876 13948
rect 21272 13932 21324 13938
rect 21272 13874 21324 13880
rect 21284 12850 21312 13874
rect 21928 13462 21956 14282
rect 21916 13456 21968 13462
rect 21836 13404 21916 13410
rect 21836 13398 21968 13404
rect 21836 13382 21956 13398
rect 21732 13184 21784 13190
rect 21836 13138 21864 13382
rect 21916 13320 21968 13326
rect 21916 13262 21968 13268
rect 21784 13132 21864 13138
rect 21732 13126 21864 13132
rect 21744 13110 21864 13126
rect 21272 12844 21324 12850
rect 21272 12786 21324 12792
rect 21836 12782 21864 13110
rect 21928 12918 21956 13262
rect 21916 12912 21968 12918
rect 21916 12854 21968 12860
rect 22020 12850 22048 14418
rect 22296 14346 22324 15438
rect 22756 15094 22784 15642
rect 22928 15564 22980 15570
rect 22928 15506 22980 15512
rect 22940 15094 22968 15506
rect 22744 15088 22796 15094
rect 22744 15030 22796 15036
rect 22928 15088 22980 15094
rect 22928 15030 22980 15036
rect 22836 14884 22888 14890
rect 22836 14826 22888 14832
rect 22652 14408 22704 14414
rect 22652 14350 22704 14356
rect 22100 14340 22152 14346
rect 22100 14282 22152 14288
rect 22284 14340 22336 14346
rect 22284 14282 22336 14288
rect 22112 13870 22140 14282
rect 22664 14074 22692 14350
rect 22652 14068 22704 14074
rect 22652 14010 22704 14016
rect 22284 13932 22336 13938
rect 22284 13874 22336 13880
rect 22100 13864 22152 13870
rect 22100 13806 22152 13812
rect 22296 13530 22324 13874
rect 22284 13524 22336 13530
rect 22284 13466 22336 13472
rect 22664 13326 22692 14010
rect 22848 14006 22876 14826
rect 22940 14618 22968 15030
rect 22928 14612 22980 14618
rect 22928 14554 22980 14560
rect 23124 14260 23152 16730
rect 23308 16726 23336 17070
rect 23296 16720 23348 16726
rect 23296 16662 23348 16668
rect 23480 16448 23532 16454
rect 23480 16390 23532 16396
rect 23492 15910 23520 16390
rect 23480 15904 23532 15910
rect 23480 15846 23532 15852
rect 23296 15564 23348 15570
rect 23296 15506 23348 15512
rect 23308 14958 23336 15506
rect 23676 15162 23704 18414
rect 23756 18080 23808 18086
rect 23756 18022 23808 18028
rect 23768 17270 23796 18022
rect 23756 17264 23808 17270
rect 23756 17206 23808 17212
rect 23848 16992 23900 16998
rect 23848 16934 23900 16940
rect 23860 16046 23888 16934
rect 23940 16652 23992 16658
rect 23940 16594 23992 16600
rect 23848 16040 23900 16046
rect 23848 15982 23900 15988
rect 23664 15156 23716 15162
rect 23664 15098 23716 15104
rect 23296 14952 23348 14958
rect 23296 14894 23348 14900
rect 23296 14272 23348 14278
rect 23124 14232 23296 14260
rect 23296 14214 23348 14220
rect 22836 14000 22888 14006
rect 22836 13942 22888 13948
rect 22652 13320 22704 13326
rect 22652 13262 22704 13268
rect 22008 12844 22060 12850
rect 22008 12786 22060 12792
rect 21824 12776 21876 12782
rect 21824 12718 21876 12724
rect 21088 12640 21140 12646
rect 21088 12582 21140 12588
rect 22020 12442 22048 12786
rect 22652 12640 22704 12646
rect 22652 12582 22704 12588
rect 20824 12406 21036 12434
rect 22008 12436 22060 12442
rect 20824 12306 20852 12406
rect 22008 12378 22060 12384
rect 20812 12300 20864 12306
rect 20812 12242 20864 12248
rect 20824 11762 20852 12242
rect 22664 12238 22692 12582
rect 22848 12238 22876 13942
rect 23308 12714 23336 14214
rect 23676 12850 23704 15098
rect 23860 14890 23888 15982
rect 23952 15094 23980 16594
rect 23940 15088 23992 15094
rect 23940 15030 23992 15036
rect 24228 15026 24256 22066
rect 24584 21548 24636 21554
rect 24584 21490 24636 21496
rect 24308 21480 24360 21486
rect 24308 21422 24360 21428
rect 24320 20398 24348 21422
rect 24596 21146 24624 21490
rect 24584 21140 24636 21146
rect 24584 21082 24636 21088
rect 24400 20936 24452 20942
rect 24400 20878 24452 20884
rect 24308 20392 24360 20398
rect 24308 20334 24360 20340
rect 24412 20262 24440 20878
rect 24952 20460 25004 20466
rect 24952 20402 25004 20408
rect 24768 20392 24820 20398
rect 24768 20334 24820 20340
rect 24400 20256 24452 20262
rect 24400 20198 24452 20204
rect 24780 19922 24808 20334
rect 24768 19916 24820 19922
rect 24768 19858 24820 19864
rect 24860 19168 24912 19174
rect 24860 19110 24912 19116
rect 24872 18766 24900 19110
rect 24860 18760 24912 18766
rect 24860 18702 24912 18708
rect 24860 17604 24912 17610
rect 24860 17546 24912 17552
rect 24872 17338 24900 17546
rect 24860 17332 24912 17338
rect 24860 17274 24912 17280
rect 24768 17196 24820 17202
rect 24768 17138 24820 17144
rect 24780 16658 24808 17138
rect 24768 16652 24820 16658
rect 24768 16594 24820 16600
rect 24964 16590 24992 20402
rect 25320 19780 25372 19786
rect 25320 19722 25372 19728
rect 25136 18624 25188 18630
rect 25136 18566 25188 18572
rect 25148 18358 25176 18566
rect 25136 18352 25188 18358
rect 25136 18294 25188 18300
rect 25332 17270 25360 19722
rect 25320 17264 25372 17270
rect 25320 17206 25372 17212
rect 24400 16584 24452 16590
rect 24400 16526 24452 16532
rect 24952 16584 25004 16590
rect 24952 16526 25004 16532
rect 24412 15366 24440 16526
rect 24400 15360 24452 15366
rect 24400 15302 24452 15308
rect 24216 15020 24268 15026
rect 24216 14962 24268 14968
rect 23848 14884 23900 14890
rect 23848 14826 23900 14832
rect 25516 13802 25544 26318
rect 25596 24812 25648 24818
rect 25596 24754 25648 24760
rect 25608 24274 25636 24754
rect 25596 24268 25648 24274
rect 25596 24210 25648 24216
rect 25608 23866 25636 24210
rect 25596 23860 25648 23866
rect 25596 23802 25648 23808
rect 25688 18760 25740 18766
rect 25688 18702 25740 18708
rect 25700 18290 25728 18702
rect 25688 18284 25740 18290
rect 25688 18226 25740 18232
rect 25792 15094 25820 28630
rect 26068 28558 26096 29990
rect 26436 29578 26464 30602
rect 26528 30258 26556 35006
rect 26516 30252 26568 30258
rect 26516 30194 26568 30200
rect 26424 29572 26476 29578
rect 26424 29514 26476 29520
rect 26056 28552 26108 28558
rect 26056 28494 26108 28500
rect 26068 28014 26096 28494
rect 26056 28008 26108 28014
rect 26056 27950 26108 27956
rect 26608 27872 26660 27878
rect 26608 27814 26660 27820
rect 26332 26240 26384 26246
rect 26332 26182 26384 26188
rect 26344 25974 26372 26182
rect 26332 25968 26384 25974
rect 26332 25910 26384 25916
rect 26516 25764 26568 25770
rect 26516 25706 26568 25712
rect 26148 25696 26200 25702
rect 26148 25638 26200 25644
rect 26160 25294 26188 25638
rect 26528 25362 26556 25706
rect 26516 25356 26568 25362
rect 26516 25298 26568 25304
rect 26148 25288 26200 25294
rect 26148 25230 26200 25236
rect 26160 24818 26188 25230
rect 26148 24812 26200 24818
rect 26148 24754 26200 24760
rect 25870 24712 25926 24721
rect 25870 24647 25872 24656
rect 25924 24647 25926 24656
rect 25872 24618 25924 24624
rect 26160 24410 26188 24754
rect 26148 24404 26200 24410
rect 26148 24346 26200 24352
rect 26240 24200 26292 24206
rect 26240 24142 26292 24148
rect 26252 23866 26280 24142
rect 26240 23860 26292 23866
rect 26240 23802 26292 23808
rect 26424 23180 26476 23186
rect 26424 23122 26476 23128
rect 26240 23044 26292 23050
rect 26240 22986 26292 22992
rect 26252 22574 26280 22986
rect 26436 22642 26464 23122
rect 26424 22636 26476 22642
rect 26424 22578 26476 22584
rect 26240 22568 26292 22574
rect 26240 22510 26292 22516
rect 25872 22160 25924 22166
rect 25872 22102 25924 22108
rect 25884 21350 25912 22102
rect 25964 22092 26016 22098
rect 25964 22034 26016 22040
rect 25976 21486 26004 22034
rect 26056 21888 26108 21894
rect 26056 21830 26108 21836
rect 25964 21480 26016 21486
rect 25964 21422 26016 21428
rect 25872 21344 25924 21350
rect 25924 21304 26004 21332
rect 25872 21286 25924 21292
rect 25884 21221 25912 21286
rect 25976 20874 26004 21304
rect 26068 20942 26096 21830
rect 26252 21146 26280 22510
rect 26332 22024 26384 22030
rect 26332 21966 26384 21972
rect 26344 21690 26372 21966
rect 26424 21956 26476 21962
rect 26424 21898 26476 21904
rect 26332 21684 26384 21690
rect 26332 21626 26384 21632
rect 26240 21140 26292 21146
rect 26240 21082 26292 21088
rect 26148 21072 26200 21078
rect 26148 21014 26200 21020
rect 26056 20936 26108 20942
rect 26056 20878 26108 20884
rect 25964 20868 26016 20874
rect 25964 20810 26016 20816
rect 25964 18692 26016 18698
rect 25964 18634 26016 18640
rect 25976 17610 26004 18634
rect 26056 18284 26108 18290
rect 26056 18226 26108 18232
rect 26068 17678 26096 18226
rect 26056 17672 26108 17678
rect 26056 17614 26108 17620
rect 25964 17604 26016 17610
rect 25964 17546 26016 17552
rect 25964 15360 26016 15366
rect 25964 15302 26016 15308
rect 25976 15094 26004 15302
rect 25780 15088 25832 15094
rect 25780 15030 25832 15036
rect 25964 15088 26016 15094
rect 25964 15030 26016 15036
rect 25792 14600 25820 15030
rect 25792 14572 25912 14600
rect 25780 14476 25832 14482
rect 25780 14418 25832 14424
rect 25688 14340 25740 14346
rect 25688 14282 25740 14288
rect 24584 13796 24636 13802
rect 24584 13738 24636 13744
rect 25504 13796 25556 13802
rect 25504 13738 25556 13744
rect 24400 13320 24452 13326
rect 24400 13262 24452 13268
rect 23664 12844 23716 12850
rect 23664 12786 23716 12792
rect 23848 12844 23900 12850
rect 23848 12786 23900 12792
rect 23296 12708 23348 12714
rect 23296 12650 23348 12656
rect 23676 12434 23704 12786
rect 23860 12442 23888 12786
rect 24412 12782 24440 13262
rect 24596 12986 24624 13738
rect 25700 13530 25728 14282
rect 25688 13524 25740 13530
rect 25688 13466 25740 13472
rect 24676 13252 24728 13258
rect 24676 13194 24728 13200
rect 24584 12980 24636 12986
rect 24584 12922 24636 12928
rect 24400 12776 24452 12782
rect 24400 12718 24452 12724
rect 23848 12436 23900 12442
rect 23676 12406 23796 12434
rect 22652 12232 22704 12238
rect 22652 12174 22704 12180
rect 22836 12232 22888 12238
rect 22836 12174 22888 12180
rect 23664 12232 23716 12238
rect 23664 12174 23716 12180
rect 21640 12164 21692 12170
rect 21640 12106 21692 12112
rect 20812 11756 20864 11762
rect 20812 11698 20864 11704
rect 20720 11552 20772 11558
rect 20720 11494 20772 11500
rect 20260 10804 20312 10810
rect 20260 10746 20312 10752
rect 20732 10266 20760 11494
rect 21652 11354 21680 12106
rect 21640 11348 21692 11354
rect 21640 11290 21692 11296
rect 20812 11076 20864 11082
rect 20812 11018 20864 11024
rect 20824 10606 20852 11018
rect 21652 10606 21680 11290
rect 20812 10600 20864 10606
rect 20812 10542 20864 10548
rect 21640 10600 21692 10606
rect 21640 10542 21692 10548
rect 20824 10470 20852 10542
rect 21916 10532 21968 10538
rect 21916 10474 21968 10480
rect 20812 10464 20864 10470
rect 20812 10406 20864 10412
rect 20720 10260 20772 10266
rect 20720 10202 20772 10208
rect 21928 10198 21956 10474
rect 21916 10192 21968 10198
rect 21916 10134 21968 10140
rect 19432 10124 19484 10130
rect 19432 10066 19484 10072
rect 20352 10056 20404 10062
rect 20352 9998 20404 10004
rect 19432 9920 19484 9926
rect 19432 9862 19484 9868
rect 18420 9580 18472 9586
rect 18420 9522 18472 9528
rect 18696 9580 18748 9586
rect 18696 9522 18748 9528
rect 19340 9580 19392 9586
rect 19340 9522 19392 9528
rect 18236 9512 18288 9518
rect 18236 9454 18288 9460
rect 19444 8974 19472 9862
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19616 9580 19668 9586
rect 19616 9522 19668 9528
rect 19628 9178 19656 9522
rect 20364 9450 20392 9998
rect 20536 9988 20588 9994
rect 20536 9930 20588 9936
rect 20548 9518 20576 9930
rect 20996 9920 21048 9926
rect 20996 9862 21048 9868
rect 22284 9920 22336 9926
rect 22284 9862 22336 9868
rect 20536 9512 20588 9518
rect 20536 9454 20588 9460
rect 20352 9444 20404 9450
rect 20352 9386 20404 9392
rect 19616 9172 19668 9178
rect 19616 9114 19668 9120
rect 19432 8968 19484 8974
rect 19432 8910 19484 8916
rect 20364 8906 20392 9386
rect 20548 8974 20576 9454
rect 20536 8968 20588 8974
rect 20536 8910 20588 8916
rect 20352 8900 20404 8906
rect 20352 8842 20404 8848
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 21008 8498 21036 9862
rect 22296 9178 22324 9862
rect 22376 9580 22428 9586
rect 22376 9522 22428 9528
rect 22284 9172 22336 9178
rect 22284 9114 22336 9120
rect 21180 8900 21232 8906
rect 21180 8842 21232 8848
rect 21192 8634 21220 8842
rect 22388 8838 22416 9522
rect 22848 8974 22876 12174
rect 23480 11144 23532 11150
rect 23480 11086 23532 11092
rect 23112 10668 23164 10674
rect 23112 10610 23164 10616
rect 23124 10266 23152 10610
rect 23112 10260 23164 10266
rect 23112 10202 23164 10208
rect 22928 10056 22980 10062
rect 23124 10010 23152 10202
rect 22928 9998 22980 10004
rect 22940 8974 22968 9998
rect 23032 9982 23152 10010
rect 23032 9450 23060 9982
rect 23112 9920 23164 9926
rect 23112 9862 23164 9868
rect 23124 9586 23152 9862
rect 23112 9580 23164 9586
rect 23112 9522 23164 9528
rect 23492 9518 23520 11086
rect 23676 10810 23704 12174
rect 23768 11762 23796 12406
rect 23848 12378 23900 12384
rect 24596 12306 24624 12922
rect 24584 12300 24636 12306
rect 24584 12242 24636 12248
rect 24688 11898 24716 13194
rect 25792 12986 25820 14418
rect 25884 14074 25912 14572
rect 25976 14414 26004 15030
rect 26160 14550 26188 21014
rect 26436 20330 26464 21898
rect 26620 20534 26648 27814
rect 26804 26518 26832 35090
rect 26884 35012 26936 35018
rect 26884 34954 26936 34960
rect 26896 34202 26924 34954
rect 27172 34746 27200 35634
rect 27160 34740 27212 34746
rect 27160 34682 27212 34688
rect 26884 34196 26936 34202
rect 26884 34138 26936 34144
rect 26896 33998 26924 34138
rect 27172 33998 27200 34682
rect 27448 34610 27476 35974
rect 27632 35698 27660 37062
rect 27724 36786 27752 37742
rect 27712 36780 27764 36786
rect 27816 36768 27844 37810
rect 28000 37330 28028 38150
rect 27988 37324 28040 37330
rect 27988 37266 28040 37272
rect 28448 37256 28500 37262
rect 28448 37198 28500 37204
rect 27896 36780 27948 36786
rect 27816 36740 27896 36768
rect 27712 36722 27764 36728
rect 27896 36722 27948 36728
rect 28080 36780 28132 36786
rect 28080 36722 28132 36728
rect 27804 36372 27856 36378
rect 27804 36314 27856 36320
rect 27712 36304 27764 36310
rect 27712 36246 27764 36252
rect 27620 35692 27672 35698
rect 27620 35634 27672 35640
rect 27528 35488 27580 35494
rect 27528 35430 27580 35436
rect 27436 34604 27488 34610
rect 27436 34546 27488 34552
rect 26884 33992 26936 33998
rect 26884 33934 26936 33940
rect 27160 33992 27212 33998
rect 27160 33934 27212 33940
rect 26976 33924 27028 33930
rect 26976 33866 27028 33872
rect 26988 33386 27016 33866
rect 27448 33862 27476 34546
rect 27540 34474 27568 35430
rect 27724 35154 27752 36246
rect 27816 36174 27844 36314
rect 27804 36168 27856 36174
rect 27804 36110 27856 36116
rect 28092 36038 28120 36722
rect 28356 36576 28408 36582
rect 28356 36518 28408 36524
rect 28080 36032 28132 36038
rect 28080 35974 28132 35980
rect 27804 35692 27856 35698
rect 27804 35634 27856 35640
rect 27712 35148 27764 35154
rect 27712 35090 27764 35096
rect 27620 35080 27672 35086
rect 27620 35022 27672 35028
rect 27632 34746 27660 35022
rect 27620 34740 27672 34746
rect 27620 34682 27672 34688
rect 27528 34468 27580 34474
rect 27528 34410 27580 34416
rect 27540 33998 27568 34410
rect 27816 34202 27844 35634
rect 28080 35284 28132 35290
rect 28080 35226 28132 35232
rect 27988 34604 28040 34610
rect 27988 34546 28040 34552
rect 27804 34196 27856 34202
rect 27804 34138 27856 34144
rect 27528 33992 27580 33998
rect 27528 33934 27580 33940
rect 27436 33856 27488 33862
rect 27436 33798 27488 33804
rect 27816 33522 27844 34138
rect 27160 33516 27212 33522
rect 27160 33458 27212 33464
rect 27804 33516 27856 33522
rect 27804 33458 27856 33464
rect 26976 33380 27028 33386
rect 26976 33322 27028 33328
rect 27068 33312 27120 33318
rect 27068 33254 27120 33260
rect 26884 32768 26936 32774
rect 26884 32710 26936 32716
rect 26896 32570 26924 32710
rect 26884 32564 26936 32570
rect 26884 32506 26936 32512
rect 27080 32502 27108 33254
rect 27068 32496 27120 32502
rect 27068 32438 27120 32444
rect 26884 32428 26936 32434
rect 26884 32370 26936 32376
rect 26896 32026 26924 32370
rect 26976 32292 27028 32298
rect 26976 32234 27028 32240
rect 26884 32020 26936 32026
rect 26884 31962 26936 31968
rect 26988 31482 27016 32234
rect 26976 31476 27028 31482
rect 26976 31418 27028 31424
rect 27172 30870 27200 33458
rect 27252 33040 27304 33046
rect 27252 32982 27304 32988
rect 27620 33040 27672 33046
rect 27620 32982 27672 32988
rect 27264 31142 27292 32982
rect 27632 32910 27660 32982
rect 27816 32978 27844 33458
rect 28000 33454 28028 34546
rect 28092 33522 28120 35226
rect 28264 35080 28316 35086
rect 28264 35022 28316 35028
rect 28276 33998 28304 35022
rect 28368 34202 28396 36518
rect 28460 35290 28488 37198
rect 28724 37120 28776 37126
rect 28724 37062 28776 37068
rect 28736 36854 28764 37062
rect 28724 36848 28776 36854
rect 28724 36790 28776 36796
rect 28828 36786 28856 38150
rect 28920 37806 28948 39578
rect 29460 39432 29512 39438
rect 29460 39374 29512 39380
rect 29472 38962 29500 39374
rect 29460 38956 29512 38962
rect 29460 38898 29512 38904
rect 29736 38956 29788 38962
rect 29736 38898 29788 38904
rect 29748 38554 29776 38898
rect 29736 38548 29788 38554
rect 29736 38490 29788 38496
rect 28908 37800 28960 37806
rect 28908 37742 28960 37748
rect 28816 36780 28868 36786
rect 28816 36722 28868 36728
rect 28920 36582 28948 37742
rect 28908 36576 28960 36582
rect 28908 36518 28960 36524
rect 29552 36032 29604 36038
rect 29552 35974 29604 35980
rect 28632 35488 28684 35494
rect 28632 35430 28684 35436
rect 28448 35284 28500 35290
rect 28448 35226 28500 35232
rect 28644 34610 28672 35430
rect 29184 35284 29236 35290
rect 29184 35226 29236 35232
rect 28908 35148 28960 35154
rect 28908 35090 28960 35096
rect 28920 34678 28948 35090
rect 29196 34746 29224 35226
rect 29460 34944 29512 34950
rect 29460 34886 29512 34892
rect 29184 34740 29236 34746
rect 29184 34682 29236 34688
rect 28908 34672 28960 34678
rect 28908 34614 28960 34620
rect 28632 34604 28684 34610
rect 28632 34546 28684 34552
rect 29000 34604 29052 34610
rect 29000 34546 29052 34552
rect 28356 34196 28408 34202
rect 28356 34138 28408 34144
rect 28264 33992 28316 33998
rect 28264 33934 28316 33940
rect 28080 33516 28132 33522
rect 28080 33458 28132 33464
rect 27988 33448 28040 33454
rect 27988 33390 28040 33396
rect 27896 33312 27948 33318
rect 27896 33254 27948 33260
rect 27804 32972 27856 32978
rect 27804 32914 27856 32920
rect 27620 32904 27672 32910
rect 27620 32846 27672 32852
rect 27712 32904 27764 32910
rect 27712 32846 27764 32852
rect 27344 32836 27396 32842
rect 27344 32778 27396 32784
rect 27356 32298 27384 32778
rect 27724 32774 27752 32846
rect 27712 32768 27764 32774
rect 27712 32710 27764 32716
rect 27724 32502 27752 32710
rect 27712 32496 27764 32502
rect 27712 32438 27764 32444
rect 27816 32434 27844 32914
rect 27908 32910 27936 33254
rect 27896 32904 27948 32910
rect 27896 32846 27948 32852
rect 28000 32570 28028 33390
rect 28092 33046 28120 33458
rect 28276 33454 28304 33934
rect 28264 33448 28316 33454
rect 28264 33390 28316 33396
rect 28080 33040 28132 33046
rect 28080 32982 28132 32988
rect 27988 32564 28040 32570
rect 27988 32506 28040 32512
rect 28092 32434 28120 32982
rect 28368 32910 28396 34138
rect 29012 33930 29040 34546
rect 29472 33998 29500 34886
rect 29564 34626 29592 35974
rect 29840 35086 29868 40054
rect 30288 40044 30340 40050
rect 30288 39986 30340 39992
rect 30012 39840 30064 39846
rect 30012 39782 30064 39788
rect 30104 39840 30156 39846
rect 30104 39782 30156 39788
rect 30024 39302 30052 39782
rect 30012 39296 30064 39302
rect 30012 39238 30064 39244
rect 30116 38350 30144 39782
rect 30300 39438 30328 39986
rect 30760 39506 30788 40394
rect 31024 40384 31076 40390
rect 31024 40326 31076 40332
rect 30748 39500 30800 39506
rect 30748 39442 30800 39448
rect 30288 39432 30340 39438
rect 30288 39374 30340 39380
rect 30104 38344 30156 38350
rect 30104 38286 30156 38292
rect 30760 37262 30788 39442
rect 31036 39438 31064 40326
rect 31128 40186 31156 40462
rect 31116 40180 31168 40186
rect 31116 40122 31168 40128
rect 31300 40112 31352 40118
rect 31300 40054 31352 40060
rect 31024 39432 31076 39438
rect 31024 39374 31076 39380
rect 30840 39364 30892 39370
rect 30840 39306 30892 39312
rect 30852 39098 30880 39306
rect 31312 39098 31340 40054
rect 31760 39976 31812 39982
rect 31760 39918 31812 39924
rect 31484 39908 31536 39914
rect 31484 39850 31536 39856
rect 31496 39438 31524 39850
rect 31484 39432 31536 39438
rect 31484 39374 31536 39380
rect 30840 39092 30892 39098
rect 30840 39034 30892 39040
rect 31300 39092 31352 39098
rect 31300 39034 31352 39040
rect 31300 37664 31352 37670
rect 31300 37606 31352 37612
rect 31312 37262 31340 37606
rect 30748 37256 30800 37262
rect 30748 37198 30800 37204
rect 31300 37256 31352 37262
rect 31300 37198 31352 37204
rect 30760 36922 30788 37198
rect 30748 36916 30800 36922
rect 30748 36858 30800 36864
rect 30932 36916 30984 36922
rect 30932 36858 30984 36864
rect 30944 35154 30972 36858
rect 31300 36576 31352 36582
rect 31300 36518 31352 36524
rect 31312 36174 31340 36518
rect 31024 36168 31076 36174
rect 31024 36110 31076 36116
rect 31300 36168 31352 36174
rect 31300 36110 31352 36116
rect 31036 35834 31064 36110
rect 31496 35834 31524 39374
rect 31772 38962 31800 39918
rect 32140 39642 32168 40462
rect 32324 39982 32352 40666
rect 32600 40186 32628 41074
rect 33060 40390 33088 41074
rect 33324 40928 33376 40934
rect 33324 40870 33376 40876
rect 33048 40384 33100 40390
rect 33048 40326 33100 40332
rect 32588 40180 32640 40186
rect 32588 40122 32640 40128
rect 32312 39976 32364 39982
rect 32312 39918 32364 39924
rect 32324 39846 32352 39918
rect 32312 39840 32364 39846
rect 32312 39782 32364 39788
rect 32128 39636 32180 39642
rect 32128 39578 32180 39584
rect 32140 39438 32168 39578
rect 32600 39574 32628 40122
rect 33060 40118 33088 40326
rect 33048 40112 33100 40118
rect 33048 40054 33100 40060
rect 32956 39908 33008 39914
rect 32956 39850 33008 39856
rect 32588 39568 32640 39574
rect 32588 39510 32640 39516
rect 32128 39432 32180 39438
rect 32128 39374 32180 39380
rect 31852 39296 31904 39302
rect 31852 39238 31904 39244
rect 31864 38962 31892 39238
rect 32600 39030 32628 39510
rect 32968 39438 32996 39850
rect 32956 39432 33008 39438
rect 32956 39374 33008 39380
rect 33060 39302 33088 40054
rect 33336 39846 33364 40870
rect 33428 40186 33456 41074
rect 36464 41070 36492 42162
rect 37844 41818 37872 42570
rect 38672 42362 38700 45200
rect 42536 45098 42564 45200
rect 42168 45070 42564 45098
rect 41786 43616 41842 43625
rect 41786 43551 41842 43560
rect 40040 43104 40092 43110
rect 40040 43046 40092 43052
rect 40052 42838 40080 43046
rect 40040 42832 40092 42838
rect 40040 42774 40092 42780
rect 41800 42770 41828 43551
rect 41788 42764 41840 42770
rect 41788 42706 41840 42712
rect 39948 42628 40000 42634
rect 39948 42570 40000 42576
rect 38660 42356 38712 42362
rect 38660 42298 38712 42304
rect 38384 42152 38436 42158
rect 38384 42094 38436 42100
rect 38396 41818 38424 42094
rect 39960 41818 39988 42570
rect 37832 41812 37884 41818
rect 37832 41754 37884 41760
rect 38384 41812 38436 41818
rect 38384 41754 38436 41760
rect 39948 41812 40000 41818
rect 39948 41754 40000 41760
rect 37924 41608 37976 41614
rect 37924 41550 37976 41556
rect 39856 41608 39908 41614
rect 39856 41550 39908 41556
rect 41510 41576 41566 41585
rect 36452 41064 36504 41070
rect 36452 41006 36504 41012
rect 33600 40928 33652 40934
rect 33600 40870 33652 40876
rect 33612 40458 33640 40870
rect 34934 40828 35242 40848
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40752 35242 40772
rect 37372 40656 37424 40662
rect 37372 40598 37424 40604
rect 35348 40520 35400 40526
rect 35348 40462 35400 40468
rect 33600 40452 33652 40458
rect 33600 40394 33652 40400
rect 35256 40384 35308 40390
rect 35256 40326 35308 40332
rect 33416 40180 33468 40186
rect 33416 40122 33468 40128
rect 35268 40118 35296 40326
rect 34520 40112 34572 40118
rect 34520 40054 34572 40060
rect 35256 40112 35308 40118
rect 35256 40054 35308 40060
rect 33324 39840 33376 39846
rect 33324 39782 33376 39788
rect 33968 39840 34020 39846
rect 33968 39782 34020 39788
rect 33980 39438 34008 39782
rect 34532 39574 34560 40054
rect 34934 39740 35242 39760
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39664 35242 39684
rect 35360 39642 35388 40462
rect 37280 40452 37332 40458
rect 37280 40394 37332 40400
rect 36084 39976 36136 39982
rect 36084 39918 36136 39924
rect 35348 39636 35400 39642
rect 35348 39578 35400 39584
rect 34520 39568 34572 39574
rect 34520 39510 34572 39516
rect 33968 39432 34020 39438
rect 33968 39374 34020 39380
rect 33324 39364 33376 39370
rect 33324 39306 33376 39312
rect 33048 39296 33100 39302
rect 33048 39238 33100 39244
rect 33232 39296 33284 39302
rect 33232 39238 33284 39244
rect 32588 39024 32640 39030
rect 32588 38966 32640 38972
rect 31760 38956 31812 38962
rect 31760 38898 31812 38904
rect 31852 38956 31904 38962
rect 31852 38898 31904 38904
rect 33060 38758 33088 39238
rect 33048 38752 33100 38758
rect 33048 38694 33100 38700
rect 33244 38418 33272 39238
rect 33336 38962 33364 39306
rect 34532 39302 34560 39510
rect 34704 39432 34756 39438
rect 34704 39374 34756 39380
rect 34520 39296 34572 39302
rect 34520 39238 34572 39244
rect 33416 39024 33468 39030
rect 33416 38966 33468 38972
rect 33324 38956 33376 38962
rect 33324 38898 33376 38904
rect 33232 38412 33284 38418
rect 33232 38354 33284 38360
rect 33244 38010 33272 38354
rect 33232 38004 33284 38010
rect 33232 37946 33284 37952
rect 33428 37874 33456 38966
rect 34060 38956 34112 38962
rect 34060 38898 34112 38904
rect 33508 38752 33560 38758
rect 33508 38694 33560 38700
rect 32036 37868 32088 37874
rect 32036 37810 32088 37816
rect 32220 37868 32272 37874
rect 32220 37810 32272 37816
rect 32404 37868 32456 37874
rect 32404 37810 32456 37816
rect 33416 37868 33468 37874
rect 33416 37810 33468 37816
rect 32048 37466 32076 37810
rect 32036 37460 32088 37466
rect 32036 37402 32088 37408
rect 32232 36650 32260 37810
rect 32416 37126 32444 37810
rect 32496 37800 32548 37806
rect 32496 37742 32548 37748
rect 32404 37120 32456 37126
rect 32404 37062 32456 37068
rect 32312 36780 32364 36786
rect 32312 36722 32364 36728
rect 32220 36644 32272 36650
rect 32220 36586 32272 36592
rect 32324 36378 32352 36722
rect 32508 36582 32536 37742
rect 32680 37732 32732 37738
rect 32680 37674 32732 37680
rect 32588 37664 32640 37670
rect 32588 37606 32640 37612
rect 32600 37194 32628 37606
rect 32692 37466 32720 37674
rect 33048 37664 33100 37670
rect 33048 37606 33100 37612
rect 32680 37460 32732 37466
rect 32680 37402 32732 37408
rect 32588 37188 32640 37194
rect 32588 37130 32640 37136
rect 32496 36576 32548 36582
rect 32496 36518 32548 36524
rect 32312 36372 32364 36378
rect 32312 36314 32364 36320
rect 32508 36310 32536 36518
rect 32496 36304 32548 36310
rect 32496 36246 32548 36252
rect 32508 36174 32536 36246
rect 32496 36168 32548 36174
rect 32496 36110 32548 36116
rect 32692 35894 32720 37402
rect 33060 37330 33088 37606
rect 33428 37466 33456 37810
rect 33416 37460 33468 37466
rect 33416 37402 33468 37408
rect 33048 37324 33100 37330
rect 33048 37266 33100 37272
rect 32956 37188 33008 37194
rect 32956 37130 33008 37136
rect 32968 36718 32996 37130
rect 32956 36712 33008 36718
rect 32956 36654 33008 36660
rect 32692 35866 32812 35894
rect 31024 35828 31076 35834
rect 31024 35770 31076 35776
rect 31484 35828 31536 35834
rect 31484 35770 31536 35776
rect 31392 35692 31444 35698
rect 31392 35634 31444 35640
rect 30932 35148 30984 35154
rect 30932 35090 30984 35096
rect 29828 35080 29880 35086
rect 29828 35022 29880 35028
rect 29644 35012 29696 35018
rect 29644 34954 29696 34960
rect 30380 35012 30432 35018
rect 30380 34954 30432 34960
rect 29656 34746 29684 34954
rect 29644 34740 29696 34746
rect 29644 34682 29696 34688
rect 29564 34610 29684 34626
rect 29564 34604 29696 34610
rect 29564 34598 29644 34604
rect 29644 34546 29696 34552
rect 29656 34066 29684 34546
rect 30392 34202 30420 34954
rect 30472 34604 30524 34610
rect 30472 34546 30524 34552
rect 30380 34196 30432 34202
rect 30380 34138 30432 34144
rect 29644 34060 29696 34066
rect 29644 34002 29696 34008
rect 29460 33992 29512 33998
rect 29460 33934 29512 33940
rect 29000 33924 29052 33930
rect 29000 33866 29052 33872
rect 29460 33516 29512 33522
rect 29460 33458 29512 33464
rect 28632 33448 28684 33454
rect 28632 33390 28684 33396
rect 28356 32904 28408 32910
rect 28356 32846 28408 32852
rect 28356 32768 28408 32774
rect 28356 32710 28408 32716
rect 28368 32502 28396 32710
rect 28644 32570 28672 33390
rect 28632 32564 28684 32570
rect 28632 32506 28684 32512
rect 28356 32496 28408 32502
rect 28356 32438 28408 32444
rect 27804 32428 27856 32434
rect 27804 32370 27856 32376
rect 28080 32428 28132 32434
rect 28080 32370 28132 32376
rect 27344 32292 27396 32298
rect 27344 32234 27396 32240
rect 28092 32042 28120 32370
rect 28092 32026 28212 32042
rect 28092 32020 28224 32026
rect 28092 32014 28172 32020
rect 28172 31962 28224 31968
rect 28172 31408 28224 31414
rect 28172 31350 28224 31356
rect 27252 31136 27304 31142
rect 27252 31078 27304 31084
rect 28080 31136 28132 31142
rect 28080 31078 28132 31084
rect 27160 30864 27212 30870
rect 27160 30806 27212 30812
rect 27436 30728 27488 30734
rect 27436 30670 27488 30676
rect 27068 30592 27120 30598
rect 27068 30534 27120 30540
rect 27080 30326 27108 30534
rect 27068 30320 27120 30326
rect 27068 30262 27120 30268
rect 27448 29510 27476 30670
rect 28092 30326 28120 31078
rect 28184 30666 28212 31350
rect 28448 31340 28500 31346
rect 28448 31282 28500 31288
rect 28460 30938 28488 31282
rect 28264 30932 28316 30938
rect 28264 30874 28316 30880
rect 28448 30932 28500 30938
rect 28448 30874 28500 30880
rect 28172 30660 28224 30666
rect 28172 30602 28224 30608
rect 28080 30320 28132 30326
rect 28080 30262 28132 30268
rect 28276 29850 28304 30874
rect 28816 30592 28868 30598
rect 28816 30534 28868 30540
rect 28828 29850 28856 30534
rect 29000 30252 29052 30258
rect 29000 30194 29052 30200
rect 28908 30048 28960 30054
rect 28908 29990 28960 29996
rect 28264 29844 28316 29850
rect 28264 29786 28316 29792
rect 28816 29844 28868 29850
rect 28816 29786 28868 29792
rect 28540 29776 28592 29782
rect 28540 29718 28592 29724
rect 27712 29640 27764 29646
rect 27712 29582 27764 29588
rect 27436 29504 27488 29510
rect 27436 29446 27488 29452
rect 27068 28552 27120 28558
rect 27068 28494 27120 28500
rect 27344 28552 27396 28558
rect 27344 28494 27396 28500
rect 27080 28082 27108 28494
rect 27356 28218 27384 28494
rect 27344 28212 27396 28218
rect 27344 28154 27396 28160
rect 27448 28098 27476 29446
rect 27724 28762 27752 29582
rect 27712 28756 27764 28762
rect 27712 28698 27764 28704
rect 27896 28756 27948 28762
rect 27896 28698 27948 28704
rect 27528 28416 27580 28422
rect 27528 28358 27580 28364
rect 27540 28218 27568 28358
rect 27528 28212 27580 28218
rect 27528 28154 27580 28160
rect 27068 28076 27120 28082
rect 27448 28070 27568 28098
rect 27068 28018 27120 28024
rect 27540 26858 27568 28070
rect 27724 28014 27752 28698
rect 27712 28008 27764 28014
rect 27712 27950 27764 27956
rect 27908 27962 27936 28698
rect 28552 28626 28580 29718
rect 28920 29646 28948 29990
rect 28908 29640 28960 29646
rect 28908 29582 28960 29588
rect 28920 29170 28948 29582
rect 28908 29164 28960 29170
rect 28908 29106 28960 29112
rect 28724 29028 28776 29034
rect 28724 28970 28776 28976
rect 27988 28620 28040 28626
rect 27988 28562 28040 28568
rect 28540 28620 28592 28626
rect 28540 28562 28592 28568
rect 28000 28490 28028 28562
rect 27988 28484 28040 28490
rect 27988 28426 28040 28432
rect 28172 28416 28224 28422
rect 28172 28358 28224 28364
rect 27988 28008 28040 28014
rect 27908 27956 27988 27962
rect 27908 27950 28040 27956
rect 27908 27934 28028 27950
rect 27908 27674 27936 27934
rect 27896 27668 27948 27674
rect 27896 27610 27948 27616
rect 27528 26852 27580 26858
rect 27528 26794 27580 26800
rect 26792 26512 26844 26518
rect 26792 26454 26844 26460
rect 27068 25968 27120 25974
rect 27068 25910 27120 25916
rect 27080 24206 27108 25910
rect 27540 25294 27568 26794
rect 27908 26382 27936 27610
rect 28184 27470 28212 28358
rect 28552 28082 28580 28562
rect 28540 28076 28592 28082
rect 28540 28018 28592 28024
rect 28172 27464 28224 27470
rect 28172 27406 28224 27412
rect 28552 27062 28580 28018
rect 28736 27130 28764 28970
rect 28908 28484 28960 28490
rect 28908 28426 28960 28432
rect 28920 27334 28948 28426
rect 29012 27538 29040 30194
rect 29000 27532 29052 27538
rect 29000 27474 29052 27480
rect 28908 27328 28960 27334
rect 28908 27270 28960 27276
rect 28724 27124 28776 27130
rect 28724 27066 28776 27072
rect 28540 27056 28592 27062
rect 28540 26998 28592 27004
rect 28540 26852 28592 26858
rect 28540 26794 28592 26800
rect 27896 26376 27948 26382
rect 27896 26318 27948 26324
rect 27620 25832 27672 25838
rect 27620 25774 27672 25780
rect 27632 25498 27660 25774
rect 27620 25492 27672 25498
rect 27620 25434 27672 25440
rect 27896 25356 27948 25362
rect 27896 25298 27948 25304
rect 27436 25288 27488 25294
rect 27436 25230 27488 25236
rect 27528 25288 27580 25294
rect 27528 25230 27580 25236
rect 27448 24410 27476 25230
rect 27620 24676 27672 24682
rect 27620 24618 27672 24624
rect 27436 24404 27488 24410
rect 27436 24346 27488 24352
rect 27068 24200 27120 24206
rect 27528 24200 27580 24206
rect 27068 24142 27120 24148
rect 27356 24148 27528 24154
rect 27356 24142 27580 24148
rect 27356 24138 27568 24142
rect 27344 24132 27568 24138
rect 27396 24126 27568 24132
rect 27344 24074 27396 24080
rect 27448 23526 27476 24126
rect 27528 23860 27580 23866
rect 27528 23802 27580 23808
rect 27436 23520 27488 23526
rect 27436 23462 27488 23468
rect 26700 23316 26752 23322
rect 26700 23258 26752 23264
rect 26712 22710 26740 23258
rect 27344 23180 27396 23186
rect 27344 23122 27396 23128
rect 26700 22704 26752 22710
rect 26700 22646 26752 22652
rect 27068 22704 27120 22710
rect 27068 22646 27120 22652
rect 26608 20528 26660 20534
rect 26608 20470 26660 20476
rect 26424 20324 26476 20330
rect 26424 20266 26476 20272
rect 26332 19780 26384 19786
rect 26332 19722 26384 19728
rect 26240 18896 26292 18902
rect 26240 18838 26292 18844
rect 26252 18358 26280 18838
rect 26240 18352 26292 18358
rect 26240 18294 26292 18300
rect 26252 18154 26280 18294
rect 26240 18148 26292 18154
rect 26240 18090 26292 18096
rect 26252 17746 26280 18090
rect 26240 17740 26292 17746
rect 26240 17682 26292 17688
rect 26344 17066 26372 19722
rect 26712 19378 26740 22646
rect 26976 22024 27028 22030
rect 26976 21966 27028 21972
rect 26988 21690 27016 21966
rect 26976 21684 27028 21690
rect 26976 21626 27028 21632
rect 26988 21010 27016 21626
rect 27080 21078 27108 22646
rect 27252 22636 27304 22642
rect 27252 22578 27304 22584
rect 27160 21888 27212 21894
rect 27160 21830 27212 21836
rect 27068 21072 27120 21078
rect 27068 21014 27120 21020
rect 26792 21004 26844 21010
rect 26792 20946 26844 20952
rect 26976 21004 27028 21010
rect 26976 20946 27028 20952
rect 26700 19372 26752 19378
rect 26700 19314 26752 19320
rect 26424 18964 26476 18970
rect 26424 18906 26476 18912
rect 26436 18766 26464 18906
rect 26424 18760 26476 18766
rect 26424 18702 26476 18708
rect 26436 18290 26464 18702
rect 26424 18284 26476 18290
rect 26424 18226 26476 18232
rect 26436 18086 26464 18226
rect 26424 18080 26476 18086
rect 26424 18022 26476 18028
rect 26436 17882 26464 18022
rect 26424 17876 26476 17882
rect 26424 17818 26476 17824
rect 26712 17814 26740 19314
rect 26700 17808 26752 17814
rect 26700 17750 26752 17756
rect 26332 17060 26384 17066
rect 26332 17002 26384 17008
rect 26516 16176 26568 16182
rect 26516 16118 26568 16124
rect 26240 15972 26292 15978
rect 26240 15914 26292 15920
rect 26252 15026 26280 15914
rect 26528 15706 26556 16118
rect 26516 15700 26568 15706
rect 26516 15642 26568 15648
rect 26240 15020 26292 15026
rect 26240 14962 26292 14968
rect 26252 14618 26280 14962
rect 26424 14884 26476 14890
rect 26424 14826 26476 14832
rect 26240 14612 26292 14618
rect 26240 14554 26292 14560
rect 26148 14544 26200 14550
rect 26148 14486 26200 14492
rect 25964 14408 26016 14414
rect 25964 14350 26016 14356
rect 25872 14068 25924 14074
rect 25872 14010 25924 14016
rect 26436 13938 26464 14826
rect 26424 13932 26476 13938
rect 26424 13874 26476 13880
rect 25780 12980 25832 12986
rect 25780 12922 25832 12928
rect 24768 12640 24820 12646
rect 24768 12582 24820 12588
rect 24780 12102 24808 12582
rect 26436 12434 26464 13874
rect 26344 12406 26464 12434
rect 25688 12164 25740 12170
rect 25688 12106 25740 12112
rect 24768 12096 24820 12102
rect 24768 12038 24820 12044
rect 24676 11892 24728 11898
rect 24676 11834 24728 11840
rect 23756 11756 23808 11762
rect 23756 11698 23808 11704
rect 24400 11756 24452 11762
rect 24400 11698 24452 11704
rect 24216 11552 24268 11558
rect 24216 11494 24268 11500
rect 24228 11150 24256 11494
rect 24412 11354 24440 11698
rect 24400 11348 24452 11354
rect 24400 11290 24452 11296
rect 24780 11150 24808 12038
rect 25700 11898 25728 12106
rect 25872 12096 25924 12102
rect 25872 12038 25924 12044
rect 25688 11892 25740 11898
rect 25688 11834 25740 11840
rect 25884 11762 25912 12038
rect 25044 11756 25096 11762
rect 25044 11698 25096 11704
rect 25872 11756 25924 11762
rect 25872 11698 25924 11704
rect 25056 11354 25084 11698
rect 25412 11552 25464 11558
rect 25412 11494 25464 11500
rect 25044 11348 25096 11354
rect 25044 11290 25096 11296
rect 25424 11150 25452 11494
rect 24216 11144 24268 11150
rect 24216 11086 24268 11092
rect 24768 11144 24820 11150
rect 24768 11086 24820 11092
rect 25412 11144 25464 11150
rect 25412 11086 25464 11092
rect 23664 10804 23716 10810
rect 23664 10746 23716 10752
rect 24228 10674 24256 11086
rect 24216 10668 24268 10674
rect 24216 10610 24268 10616
rect 23664 10192 23716 10198
rect 23664 10134 23716 10140
rect 23676 9586 23704 10134
rect 24228 10130 24256 10610
rect 24780 10554 24808 11086
rect 24952 10668 25004 10674
rect 24952 10610 25004 10616
rect 24860 10600 24912 10606
rect 24780 10548 24860 10554
rect 24780 10542 24912 10548
rect 24780 10526 24900 10542
rect 24216 10124 24268 10130
rect 24216 10066 24268 10072
rect 24780 10010 24808 10526
rect 24860 10056 24912 10062
rect 24780 10004 24860 10010
rect 24780 9998 24912 10004
rect 24780 9982 24900 9998
rect 24676 9920 24728 9926
rect 24676 9862 24728 9868
rect 24688 9586 24716 9862
rect 23664 9580 23716 9586
rect 23664 9522 23716 9528
rect 24676 9580 24728 9586
rect 24676 9522 24728 9528
rect 23480 9512 23532 9518
rect 23480 9454 23532 9460
rect 23020 9444 23072 9450
rect 23020 9386 23072 9392
rect 22836 8968 22888 8974
rect 22836 8910 22888 8916
rect 22928 8968 22980 8974
rect 22928 8910 22980 8916
rect 22376 8832 22428 8838
rect 22376 8774 22428 8780
rect 22940 8634 22968 8910
rect 23032 8906 23060 9386
rect 23492 8974 23520 9454
rect 23848 9376 23900 9382
rect 23848 9318 23900 9324
rect 23480 8968 23532 8974
rect 23480 8910 23532 8916
rect 23020 8900 23072 8906
rect 23020 8842 23072 8848
rect 21180 8628 21232 8634
rect 21180 8570 21232 8576
rect 22928 8628 22980 8634
rect 22928 8570 22980 8576
rect 23860 8566 23888 9318
rect 23848 8560 23900 8566
rect 23848 8502 23900 8508
rect 24780 8498 24808 9982
rect 24964 9722 24992 10610
rect 25412 10464 25464 10470
rect 25412 10406 25464 10412
rect 24952 9716 25004 9722
rect 24952 9658 25004 9664
rect 25424 9586 25452 10406
rect 25596 9988 25648 9994
rect 25596 9930 25648 9936
rect 25608 9722 25636 9930
rect 25596 9716 25648 9722
rect 25596 9658 25648 9664
rect 25412 9580 25464 9586
rect 25412 9522 25464 9528
rect 20996 8492 21048 8498
rect 20996 8434 21048 8440
rect 24768 8492 24820 8498
rect 24768 8434 24820 8440
rect 26344 7750 26372 12406
rect 26804 11354 26832 20946
rect 27172 20942 27200 21830
rect 27264 21690 27292 22578
rect 27356 22030 27384 23122
rect 27540 22710 27568 23802
rect 27528 22704 27580 22710
rect 27528 22646 27580 22652
rect 27528 22568 27580 22574
rect 27528 22510 27580 22516
rect 27436 22092 27488 22098
rect 27436 22034 27488 22040
rect 27344 22024 27396 22030
rect 27344 21966 27396 21972
rect 27344 21888 27396 21894
rect 27344 21830 27396 21836
rect 27252 21684 27304 21690
rect 27252 21626 27304 21632
rect 27356 21486 27384 21830
rect 27344 21480 27396 21486
rect 27344 21422 27396 21428
rect 27448 21010 27476 22034
rect 27540 21962 27568 22510
rect 27528 21956 27580 21962
rect 27528 21898 27580 21904
rect 27540 21350 27568 21898
rect 27528 21344 27580 21350
rect 27528 21286 27580 21292
rect 27436 21004 27488 21010
rect 27436 20946 27488 20952
rect 27160 20936 27212 20942
rect 27160 20878 27212 20884
rect 27448 20058 27476 20946
rect 27436 20052 27488 20058
rect 27436 19994 27488 20000
rect 27068 19304 27120 19310
rect 27068 19246 27120 19252
rect 26976 18760 27028 18766
rect 26976 18702 27028 18708
rect 26988 18222 27016 18702
rect 27080 18630 27108 19246
rect 27068 18624 27120 18630
rect 27068 18566 27120 18572
rect 26976 18216 27028 18222
rect 26976 18158 27028 18164
rect 26988 17746 27016 18158
rect 26976 17740 27028 17746
rect 26976 17682 27028 17688
rect 27080 17134 27108 18566
rect 27252 17536 27304 17542
rect 27252 17478 27304 17484
rect 27068 17128 27120 17134
rect 27068 17070 27120 17076
rect 27264 16114 27292 17478
rect 27632 17270 27660 24618
rect 27908 24410 27936 25298
rect 27896 24404 27948 24410
rect 27896 24346 27948 24352
rect 27712 24200 27764 24206
rect 27712 24142 27764 24148
rect 27724 23798 27752 24142
rect 27712 23792 27764 23798
rect 27712 23734 27764 23740
rect 27804 23724 27856 23730
rect 27804 23666 27856 23672
rect 27988 23724 28040 23730
rect 27988 23666 28040 23672
rect 27816 23322 27844 23666
rect 27804 23316 27856 23322
rect 27804 23258 27856 23264
rect 28000 22642 28028 23666
rect 28552 23594 28580 26794
rect 28632 25764 28684 25770
rect 28632 25706 28684 25712
rect 28644 25498 28672 25706
rect 28632 25492 28684 25498
rect 28632 25434 28684 25440
rect 28644 25294 28672 25434
rect 28736 25378 28764 27066
rect 28816 26988 28868 26994
rect 28816 26930 28868 26936
rect 28828 26586 28856 26930
rect 28920 26926 28948 27270
rect 29012 27130 29040 27474
rect 29000 27124 29052 27130
rect 29000 27066 29052 27072
rect 28908 26920 28960 26926
rect 28908 26862 28960 26868
rect 28816 26580 28868 26586
rect 28816 26522 28868 26528
rect 28828 25888 28856 26522
rect 28908 25900 28960 25906
rect 28828 25860 28908 25888
rect 28908 25842 28960 25848
rect 29000 25696 29052 25702
rect 29000 25638 29052 25644
rect 28736 25362 28948 25378
rect 28736 25356 28960 25362
rect 28736 25350 28908 25356
rect 28908 25298 28960 25304
rect 29012 25294 29040 25638
rect 28632 25288 28684 25294
rect 28632 25230 28684 25236
rect 29000 25288 29052 25294
rect 29000 25230 29052 25236
rect 28644 24886 28672 25230
rect 28632 24880 28684 24886
rect 28632 24822 28684 24828
rect 28540 23588 28592 23594
rect 28540 23530 28592 23536
rect 28080 23112 28132 23118
rect 28080 23054 28132 23060
rect 27988 22636 28040 22642
rect 27988 22578 28040 22584
rect 28092 22166 28120 23054
rect 28644 22642 28672 24822
rect 29012 24750 29040 25230
rect 29092 24812 29144 24818
rect 29092 24754 29144 24760
rect 29000 24744 29052 24750
rect 29000 24686 29052 24692
rect 28724 24336 28776 24342
rect 28724 24278 28776 24284
rect 28736 24206 28764 24278
rect 28724 24200 28776 24206
rect 28724 24142 28776 24148
rect 28736 23798 28764 24142
rect 28724 23792 28776 23798
rect 28724 23734 28776 23740
rect 28632 22636 28684 22642
rect 28632 22578 28684 22584
rect 28080 22160 28132 22166
rect 28080 22102 28132 22108
rect 28092 21622 28120 22102
rect 29104 21894 29132 24754
rect 29472 24682 29500 33458
rect 30484 32722 30512 34546
rect 30944 34202 30972 35090
rect 31404 34746 31432 35634
rect 32784 35562 32812 35866
rect 32772 35556 32824 35562
rect 32772 35498 32824 35504
rect 32784 35154 32812 35498
rect 32956 35488 33008 35494
rect 32956 35430 33008 35436
rect 32772 35148 32824 35154
rect 32772 35090 32824 35096
rect 32496 35080 32548 35086
rect 32496 35022 32548 35028
rect 32312 34944 32364 34950
rect 32312 34886 32364 34892
rect 31392 34740 31444 34746
rect 31392 34682 31444 34688
rect 30932 34196 30984 34202
rect 30932 34138 30984 34144
rect 31668 34196 31720 34202
rect 31668 34138 31720 34144
rect 31484 33924 31536 33930
rect 31484 33866 31536 33872
rect 31496 33590 31524 33866
rect 31484 33584 31536 33590
rect 31484 33526 31536 33532
rect 31680 33522 31708 34138
rect 31944 34128 31996 34134
rect 31944 34070 31996 34076
rect 31668 33516 31720 33522
rect 31668 33458 31720 33464
rect 31956 32910 31984 34070
rect 32128 33992 32180 33998
rect 32128 33934 32180 33940
rect 32036 33448 32088 33454
rect 32036 33390 32088 33396
rect 32048 33114 32076 33390
rect 32036 33108 32088 33114
rect 32036 33050 32088 33056
rect 32140 32978 32168 33934
rect 32128 32972 32180 32978
rect 32128 32914 32180 32920
rect 32324 32910 32352 34886
rect 32508 34202 32536 35022
rect 32588 34740 32640 34746
rect 32588 34682 32640 34688
rect 32496 34196 32548 34202
rect 32496 34138 32548 34144
rect 32508 33590 32536 34138
rect 32600 33998 32628 34682
rect 32772 34672 32824 34678
rect 32968 34626 32996 35430
rect 33060 34746 33088 37266
rect 33324 36100 33376 36106
rect 33324 36042 33376 36048
rect 33336 35698 33364 36042
rect 33324 35692 33376 35698
rect 33324 35634 33376 35640
rect 33232 35216 33284 35222
rect 33232 35158 33284 35164
rect 33140 35080 33192 35086
rect 33140 35022 33192 35028
rect 33048 34740 33100 34746
rect 33048 34682 33100 34688
rect 32824 34620 32996 34626
rect 32772 34614 32996 34620
rect 32784 34598 32996 34614
rect 32968 34134 32996 34598
rect 33152 34474 33180 35022
rect 33140 34468 33192 34474
rect 33140 34410 33192 34416
rect 33048 34400 33100 34406
rect 33048 34342 33100 34348
rect 32956 34128 33008 34134
rect 32956 34070 33008 34076
rect 32588 33992 32640 33998
rect 32588 33934 32640 33940
rect 32496 33584 32548 33590
rect 32496 33526 32548 33532
rect 32680 33516 32732 33522
rect 32680 33458 32732 33464
rect 32692 33114 32720 33458
rect 33060 33436 33088 34342
rect 33152 33998 33180 34410
rect 33140 33992 33192 33998
rect 33140 33934 33192 33940
rect 33140 33448 33192 33454
rect 33060 33408 33140 33436
rect 32680 33108 32732 33114
rect 32680 33050 32732 33056
rect 33060 32910 33088 33408
rect 33140 33390 33192 33396
rect 33244 33318 33272 35158
rect 33336 35018 33364 35634
rect 33520 35630 33548 38694
rect 34072 38010 34100 38898
rect 34152 38752 34204 38758
rect 34152 38694 34204 38700
rect 34164 38214 34192 38694
rect 34152 38208 34204 38214
rect 34152 38150 34204 38156
rect 34060 38004 34112 38010
rect 34060 37946 34112 37952
rect 34072 37874 34100 37946
rect 33600 37868 33652 37874
rect 33600 37810 33652 37816
rect 34060 37868 34112 37874
rect 34060 37810 34112 37816
rect 33612 36378 33640 37810
rect 34164 37262 34192 38150
rect 34152 37256 34204 37262
rect 34152 37198 34204 37204
rect 34164 36922 34192 37198
rect 34152 36916 34204 36922
rect 34152 36858 34204 36864
rect 33600 36372 33652 36378
rect 33600 36314 33652 36320
rect 34164 36106 34192 36858
rect 34532 36854 34560 39238
rect 34716 38350 34744 39374
rect 34934 38652 35242 38672
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38576 35242 38596
rect 34980 38480 35032 38486
rect 34980 38422 35032 38428
rect 34704 38344 34756 38350
rect 34704 38286 34756 38292
rect 34796 38344 34848 38350
rect 34796 38286 34848 38292
rect 34716 37210 34744 38286
rect 34808 37466 34836 38286
rect 34992 37874 35020 38422
rect 36096 38418 36124 39918
rect 37292 39642 37320 40394
rect 37384 40050 37412 40598
rect 37740 40520 37792 40526
rect 37740 40462 37792 40468
rect 37648 40384 37700 40390
rect 37648 40326 37700 40332
rect 37660 40186 37688 40326
rect 37648 40180 37700 40186
rect 37648 40122 37700 40128
rect 37372 40044 37424 40050
rect 37372 39986 37424 39992
rect 37280 39636 37332 39642
rect 37280 39578 37332 39584
rect 37660 39438 37688 40122
rect 37752 39506 37780 40462
rect 37740 39500 37792 39506
rect 37740 39442 37792 39448
rect 37648 39432 37700 39438
rect 37648 39374 37700 39380
rect 37556 39296 37608 39302
rect 37556 39238 37608 39244
rect 37280 38956 37332 38962
rect 37280 38898 37332 38904
rect 37372 38956 37424 38962
rect 37372 38898 37424 38904
rect 36360 38752 36412 38758
rect 36360 38694 36412 38700
rect 36084 38412 36136 38418
rect 36084 38354 36136 38360
rect 34980 37868 35032 37874
rect 34980 37810 35032 37816
rect 36096 37806 36124 38354
rect 36372 38350 36400 38694
rect 36360 38344 36412 38350
rect 36360 38286 36412 38292
rect 37292 38010 37320 38898
rect 37384 38214 37412 38898
rect 37464 38752 37516 38758
rect 37464 38694 37516 38700
rect 37372 38208 37424 38214
rect 37372 38150 37424 38156
rect 37280 38004 37332 38010
rect 37280 37946 37332 37952
rect 37280 37868 37332 37874
rect 37280 37810 37332 37816
rect 36084 37800 36136 37806
rect 36084 37742 36136 37748
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 37292 37466 37320 37810
rect 34796 37460 34848 37466
rect 34796 37402 34848 37408
rect 37280 37460 37332 37466
rect 37280 37402 37332 37408
rect 35348 37324 35400 37330
rect 35348 37266 35400 37272
rect 34796 37256 34848 37262
rect 34716 37204 34796 37210
rect 34716 37198 34848 37204
rect 34716 37182 34836 37198
rect 34520 36848 34572 36854
rect 34520 36790 34572 36796
rect 34244 36372 34296 36378
rect 34244 36314 34296 36320
rect 33692 36100 33744 36106
rect 33692 36042 33744 36048
rect 34152 36100 34204 36106
rect 34152 36042 34204 36048
rect 33704 35698 33732 36042
rect 33692 35692 33744 35698
rect 33692 35634 33744 35640
rect 33508 35624 33560 35630
rect 33508 35566 33560 35572
rect 34060 35624 34112 35630
rect 34060 35566 34112 35572
rect 34072 35290 34100 35566
rect 34060 35284 34112 35290
rect 34060 35226 34112 35232
rect 34256 35086 34284 36314
rect 34532 36242 34560 36790
rect 34716 36786 34744 37182
rect 34704 36780 34756 36786
rect 34704 36722 34756 36728
rect 34520 36236 34572 36242
rect 34520 36178 34572 36184
rect 34716 36038 34744 36722
rect 34796 36576 34848 36582
rect 34796 36518 34848 36524
rect 34704 36032 34756 36038
rect 34704 35974 34756 35980
rect 34704 35760 34756 35766
rect 34704 35702 34756 35708
rect 34428 35488 34480 35494
rect 34428 35430 34480 35436
rect 34520 35488 34572 35494
rect 34520 35430 34572 35436
rect 34440 35290 34468 35430
rect 34428 35284 34480 35290
rect 34428 35226 34480 35232
rect 34244 35080 34296 35086
rect 34244 35022 34296 35028
rect 33324 35012 33376 35018
rect 33324 34954 33376 34960
rect 34532 34610 34560 35430
rect 34520 34604 34572 34610
rect 34520 34546 34572 34552
rect 34336 34128 34388 34134
rect 34336 34070 34388 34076
rect 33416 33992 33468 33998
rect 33416 33934 33468 33940
rect 34244 33992 34296 33998
rect 34244 33934 34296 33940
rect 33428 33386 33456 33934
rect 33968 33924 34020 33930
rect 33968 33866 34020 33872
rect 33980 33522 34008 33866
rect 34060 33856 34112 33862
rect 34060 33798 34112 33804
rect 34072 33522 34100 33798
rect 34256 33590 34284 33934
rect 34244 33584 34296 33590
rect 34244 33526 34296 33532
rect 33968 33516 34020 33522
rect 33968 33458 34020 33464
rect 34060 33516 34112 33522
rect 34060 33458 34112 33464
rect 33416 33380 33468 33386
rect 33416 33322 33468 33328
rect 33140 33312 33192 33318
rect 33140 33254 33192 33260
rect 33232 33312 33284 33318
rect 33232 33254 33284 33260
rect 33152 32910 33180 33254
rect 33244 32978 33272 33254
rect 33980 33046 34008 33458
rect 34348 33454 34376 34070
rect 34336 33448 34388 33454
rect 34336 33390 34388 33396
rect 34716 33114 34744 35702
rect 34808 35698 34836 36518
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 34796 35692 34848 35698
rect 34796 35634 34848 35640
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 35360 35222 35388 37266
rect 37384 37262 37412 38150
rect 37476 37670 37504 38694
rect 37464 37664 37516 37670
rect 37464 37606 37516 37612
rect 37372 37256 37424 37262
rect 37372 37198 37424 37204
rect 35992 36848 36044 36854
rect 35992 36790 36044 36796
rect 35440 36780 35492 36786
rect 35440 36722 35492 36728
rect 35452 36378 35480 36722
rect 35440 36372 35492 36378
rect 35440 36314 35492 36320
rect 35900 36100 35952 36106
rect 35900 36042 35952 36048
rect 35912 35562 35940 36042
rect 35900 35556 35952 35562
rect 35900 35498 35952 35504
rect 36004 35290 36032 36790
rect 36176 36712 36228 36718
rect 36176 36654 36228 36660
rect 36188 36242 36216 36654
rect 36176 36236 36228 36242
rect 36176 36178 36228 36184
rect 36728 36100 36780 36106
rect 36728 36042 36780 36048
rect 36740 35562 36768 36042
rect 37568 35894 37596 39238
rect 37660 38962 37688 39374
rect 37752 38962 37780 39442
rect 37648 38956 37700 38962
rect 37648 38898 37700 38904
rect 37740 38956 37792 38962
rect 37740 38898 37792 38904
rect 37660 38418 37688 38898
rect 37752 38826 37780 38898
rect 37740 38820 37792 38826
rect 37740 38762 37792 38768
rect 37648 38412 37700 38418
rect 37648 38354 37700 38360
rect 37660 37194 37688 38354
rect 37648 37188 37700 37194
rect 37648 37130 37700 37136
rect 37752 37126 37780 38762
rect 37740 37120 37792 37126
rect 37740 37062 37792 37068
rect 37476 35866 37596 35894
rect 37476 35630 37504 35866
rect 37464 35624 37516 35630
rect 37464 35566 37516 35572
rect 36728 35556 36780 35562
rect 36728 35498 36780 35504
rect 37648 35488 37700 35494
rect 37648 35430 37700 35436
rect 35992 35284 36044 35290
rect 35992 35226 36044 35232
rect 35348 35216 35400 35222
rect 35348 35158 35400 35164
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 35360 34066 35388 35158
rect 36084 35148 36136 35154
rect 36084 35090 36136 35096
rect 35900 35012 35952 35018
rect 35900 34954 35952 34960
rect 35348 34060 35400 34066
rect 35348 34002 35400 34008
rect 35440 33992 35492 33998
rect 35440 33934 35492 33940
rect 34796 33856 34848 33862
rect 34796 33798 34848 33804
rect 34704 33108 34756 33114
rect 34704 33050 34756 33056
rect 33968 33040 34020 33046
rect 33968 32982 34020 32988
rect 33232 32972 33284 32978
rect 33232 32914 33284 32920
rect 31944 32904 31996 32910
rect 31944 32846 31996 32852
rect 32312 32904 32364 32910
rect 32312 32846 32364 32852
rect 33048 32904 33100 32910
rect 33048 32846 33100 32852
rect 33140 32904 33192 32910
rect 33140 32846 33192 32852
rect 30932 32836 30984 32842
rect 30932 32778 30984 32784
rect 30300 32694 30512 32722
rect 30300 31822 30328 32694
rect 30656 32428 30708 32434
rect 30656 32370 30708 32376
rect 30472 32292 30524 32298
rect 30472 32234 30524 32240
rect 30380 31952 30432 31958
rect 30380 31894 30432 31900
rect 29644 31816 29696 31822
rect 29644 31758 29696 31764
rect 30288 31816 30340 31822
rect 30288 31758 30340 31764
rect 29656 31278 29684 31758
rect 30392 31278 30420 31894
rect 30484 31754 30512 32234
rect 30668 31958 30696 32370
rect 30656 31952 30708 31958
rect 30656 31894 30708 31900
rect 30472 31748 30524 31754
rect 30472 31690 30524 31696
rect 30840 31680 30892 31686
rect 30840 31622 30892 31628
rect 29644 31272 29696 31278
rect 29644 31214 29696 31220
rect 30380 31272 30432 31278
rect 30380 31214 30432 31220
rect 30748 31272 30800 31278
rect 30748 31214 30800 31220
rect 30472 30864 30524 30870
rect 30472 30806 30524 30812
rect 30012 30660 30064 30666
rect 30012 30602 30064 30608
rect 30024 30258 30052 30602
rect 30484 30394 30512 30806
rect 30656 30728 30708 30734
rect 30656 30670 30708 30676
rect 30472 30388 30524 30394
rect 30472 30330 30524 30336
rect 30668 30258 30696 30670
rect 30760 30410 30788 31214
rect 30852 30734 30880 31622
rect 30840 30728 30892 30734
rect 30840 30670 30892 30676
rect 30944 30682 30972 32778
rect 33980 32570 34008 32982
rect 33968 32564 34020 32570
rect 33968 32506 34020 32512
rect 34808 32502 34836 33798
rect 35452 33590 35480 33934
rect 35624 33856 35676 33862
rect 35624 33798 35676 33804
rect 35440 33584 35492 33590
rect 35440 33526 35492 33532
rect 35452 33454 35480 33526
rect 35440 33448 35492 33454
rect 35492 33408 35572 33436
rect 35440 33390 35492 33396
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 35348 33040 35400 33046
rect 35348 32982 35400 32988
rect 34796 32496 34848 32502
rect 34796 32438 34848 32444
rect 31760 32360 31812 32366
rect 31760 32302 31812 32308
rect 34796 32360 34848 32366
rect 34796 32302 34848 32308
rect 31772 31822 31800 32302
rect 32128 31884 32180 31890
rect 32128 31826 32180 31832
rect 31760 31816 31812 31822
rect 31760 31758 31812 31764
rect 32140 31482 32168 31826
rect 34808 31822 34836 32302
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 32772 31816 32824 31822
rect 32772 31758 32824 31764
rect 34796 31816 34848 31822
rect 34796 31758 34848 31764
rect 32128 31476 32180 31482
rect 32128 31418 32180 31424
rect 31300 31408 31352 31414
rect 31300 31350 31352 31356
rect 31116 31136 31168 31142
rect 31116 31078 31168 31084
rect 31128 30938 31156 31078
rect 31116 30932 31168 30938
rect 31116 30874 31168 30880
rect 31024 30728 31076 30734
rect 30944 30676 31024 30682
rect 30944 30670 31076 30676
rect 30852 30598 30880 30670
rect 30944 30654 31064 30670
rect 30840 30592 30892 30598
rect 30840 30534 30892 30540
rect 30760 30382 30880 30410
rect 30012 30252 30064 30258
rect 30012 30194 30064 30200
rect 30656 30252 30708 30258
rect 30656 30194 30708 30200
rect 29552 30048 29604 30054
rect 29552 29990 29604 29996
rect 30472 30048 30524 30054
rect 30472 29990 30524 29996
rect 29564 29306 29592 29990
rect 30484 29646 30512 29990
rect 30668 29714 30696 30194
rect 30656 29708 30708 29714
rect 30656 29650 30708 29656
rect 30472 29640 30524 29646
rect 30472 29582 30524 29588
rect 30564 29640 30616 29646
rect 30564 29582 30616 29588
rect 30380 29572 30432 29578
rect 30380 29514 30432 29520
rect 29552 29300 29604 29306
rect 29552 29242 29604 29248
rect 30392 29034 30420 29514
rect 30484 29306 30512 29582
rect 30472 29300 30524 29306
rect 30472 29242 30524 29248
rect 30484 29170 30512 29242
rect 30472 29164 30524 29170
rect 30472 29106 30524 29112
rect 30380 29028 30432 29034
rect 30380 28970 30432 28976
rect 29552 28076 29604 28082
rect 29552 28018 29604 28024
rect 29564 26858 29592 28018
rect 29828 27872 29880 27878
rect 29828 27814 29880 27820
rect 29840 27538 29868 27814
rect 30392 27606 30420 28970
rect 30472 28960 30524 28966
rect 30472 28902 30524 28908
rect 30484 28762 30512 28902
rect 30472 28756 30524 28762
rect 30472 28698 30524 28704
rect 30576 28558 30604 29582
rect 30748 29096 30800 29102
rect 30748 29038 30800 29044
rect 30760 28626 30788 29038
rect 30748 28620 30800 28626
rect 30748 28562 30800 28568
rect 30564 28552 30616 28558
rect 30564 28494 30616 28500
rect 30576 28082 30604 28494
rect 30564 28076 30616 28082
rect 30564 28018 30616 28024
rect 30760 28014 30788 28562
rect 30748 28008 30800 28014
rect 30748 27950 30800 27956
rect 30656 27940 30708 27946
rect 30656 27882 30708 27888
rect 30668 27674 30696 27882
rect 30656 27668 30708 27674
rect 30656 27610 30708 27616
rect 30380 27600 30432 27606
rect 30380 27542 30432 27548
rect 29828 27532 29880 27538
rect 29828 27474 29880 27480
rect 29552 26852 29604 26858
rect 29552 26794 29604 26800
rect 29840 26246 29868 27474
rect 30288 26308 30340 26314
rect 30288 26250 30340 26256
rect 29828 26240 29880 26246
rect 29828 26182 29880 26188
rect 30196 25152 30248 25158
rect 30196 25094 30248 25100
rect 29552 24812 29604 24818
rect 29552 24754 29604 24760
rect 29460 24676 29512 24682
rect 29460 24618 29512 24624
rect 29564 24410 29592 24754
rect 29552 24404 29604 24410
rect 29552 24346 29604 24352
rect 30208 24274 30236 25094
rect 30300 24614 30328 26250
rect 30564 26036 30616 26042
rect 30564 25978 30616 25984
rect 30472 25832 30524 25838
rect 30472 25774 30524 25780
rect 30484 25498 30512 25774
rect 30380 25492 30432 25498
rect 30380 25434 30432 25440
rect 30472 25492 30524 25498
rect 30472 25434 30524 25440
rect 30392 24954 30420 25434
rect 30380 24948 30432 24954
rect 30380 24890 30432 24896
rect 30288 24608 30340 24614
rect 30288 24550 30340 24556
rect 30380 24336 30432 24342
rect 30380 24278 30432 24284
rect 30196 24268 30248 24274
rect 30196 24210 30248 24216
rect 30392 23730 30420 24278
rect 30484 23866 30512 25434
rect 30576 25158 30604 25978
rect 30760 25226 30788 27950
rect 30852 27470 30880 30382
rect 30944 30258 30972 30654
rect 30932 30252 30984 30258
rect 30932 30194 30984 30200
rect 31208 30252 31260 30258
rect 31208 30194 31260 30200
rect 31024 29640 31076 29646
rect 31024 29582 31076 29588
rect 31036 28422 31064 29582
rect 31220 28626 31248 30194
rect 31312 29850 31340 31350
rect 31852 30864 31904 30870
rect 31772 30824 31852 30852
rect 31668 30660 31720 30666
rect 31772 30648 31800 30824
rect 31852 30806 31904 30812
rect 32784 30734 32812 31758
rect 35360 31414 35388 32982
rect 35544 32842 35572 33408
rect 35532 32836 35584 32842
rect 35532 32778 35584 32784
rect 35544 32434 35572 32778
rect 35636 32502 35664 33798
rect 35912 33046 35940 34954
rect 36096 34134 36124 35090
rect 37372 34604 37424 34610
rect 37372 34546 37424 34552
rect 37384 34202 37412 34546
rect 37660 34542 37688 35430
rect 37648 34536 37700 34542
rect 37648 34478 37700 34484
rect 37372 34196 37424 34202
rect 37372 34138 37424 34144
rect 36084 34128 36136 34134
rect 36084 34070 36136 34076
rect 35992 33652 36044 33658
rect 35992 33594 36044 33600
rect 36004 33386 36032 33594
rect 35992 33380 36044 33386
rect 35992 33322 36044 33328
rect 36096 33318 36124 34070
rect 36912 33992 36964 33998
rect 36912 33934 36964 33940
rect 37188 33992 37240 33998
rect 37188 33934 37240 33940
rect 36176 33924 36228 33930
rect 36176 33866 36228 33872
rect 36188 33522 36216 33866
rect 36268 33856 36320 33862
rect 36268 33798 36320 33804
rect 36360 33856 36412 33862
rect 36360 33798 36412 33804
rect 36280 33658 36308 33798
rect 36268 33652 36320 33658
rect 36268 33594 36320 33600
rect 36176 33516 36228 33522
rect 36176 33458 36228 33464
rect 36084 33312 36136 33318
rect 36084 33254 36136 33260
rect 36280 33114 36308 33594
rect 36268 33108 36320 33114
rect 36268 33050 36320 33056
rect 36372 33046 36400 33798
rect 36452 33448 36504 33454
rect 36452 33390 36504 33396
rect 36464 33114 36492 33390
rect 36924 33386 36952 33934
rect 37200 33454 37228 33934
rect 37280 33856 37332 33862
rect 37280 33798 37332 33804
rect 37188 33448 37240 33454
rect 37188 33390 37240 33396
rect 36912 33380 36964 33386
rect 36912 33322 36964 33328
rect 36636 33312 36688 33318
rect 36636 33254 36688 33260
rect 36452 33108 36504 33114
rect 36452 33050 36504 33056
rect 35900 33040 35952 33046
rect 35900 32982 35952 32988
rect 36360 33040 36412 33046
rect 36360 32982 36412 32988
rect 36372 32910 36400 32982
rect 35716 32904 35768 32910
rect 35716 32846 35768 32852
rect 36360 32904 36412 32910
rect 36360 32846 36412 32852
rect 35624 32496 35676 32502
rect 35624 32438 35676 32444
rect 35728 32434 35756 32846
rect 36084 32496 36136 32502
rect 36084 32438 36136 32444
rect 35532 32428 35584 32434
rect 35532 32370 35584 32376
rect 35716 32428 35768 32434
rect 35716 32370 35768 32376
rect 35440 32224 35492 32230
rect 35440 32166 35492 32172
rect 35452 31822 35480 32166
rect 35728 32026 35756 32370
rect 35716 32020 35768 32026
rect 35716 31962 35768 31968
rect 35440 31816 35492 31822
rect 35440 31758 35492 31764
rect 36096 31754 36124 32438
rect 36648 31822 36676 33254
rect 36924 32842 36952 33322
rect 36912 32836 36964 32842
rect 36912 32778 36964 32784
rect 36924 32570 36952 32778
rect 36912 32564 36964 32570
rect 36912 32506 36964 32512
rect 37292 32434 37320 33798
rect 37556 33652 37608 33658
rect 37556 33594 37608 33600
rect 37568 33522 37596 33594
rect 37556 33516 37608 33522
rect 37556 33458 37608 33464
rect 37568 33114 37596 33458
rect 37556 33108 37608 33114
rect 37556 33050 37608 33056
rect 37372 32836 37424 32842
rect 37372 32778 37424 32784
rect 37384 32570 37412 32778
rect 37372 32564 37424 32570
rect 37372 32506 37424 32512
rect 37280 32428 37332 32434
rect 37280 32370 37332 32376
rect 36636 31816 36688 31822
rect 36636 31758 36688 31764
rect 36004 31726 36124 31754
rect 35348 31408 35400 31414
rect 35348 31350 35400 31356
rect 34796 31204 34848 31210
rect 34796 31146 34848 31152
rect 32772 30728 32824 30734
rect 31852 30706 31904 30712
rect 32772 30670 32824 30676
rect 31852 30648 31904 30654
rect 31720 30620 31800 30648
rect 31668 30602 31720 30608
rect 31484 30252 31536 30258
rect 31484 30194 31536 30200
rect 31300 29844 31352 29850
rect 31300 29786 31352 29792
rect 31392 29844 31444 29850
rect 31392 29786 31444 29792
rect 31300 29096 31352 29102
rect 31404 29084 31432 29786
rect 31496 29170 31524 30194
rect 31484 29164 31536 29170
rect 31484 29106 31536 29112
rect 31668 29164 31720 29170
rect 31668 29106 31720 29112
rect 31352 29056 31432 29084
rect 31300 29038 31352 29044
rect 31576 29028 31628 29034
rect 31576 28970 31628 28976
rect 31300 28756 31352 28762
rect 31300 28698 31352 28704
rect 31208 28620 31260 28626
rect 31208 28562 31260 28568
rect 31024 28416 31076 28422
rect 31024 28358 31076 28364
rect 31116 28416 31168 28422
rect 31116 28358 31168 28364
rect 31036 27946 31064 28358
rect 31024 27940 31076 27946
rect 31024 27882 31076 27888
rect 31128 27674 31156 28358
rect 31220 28218 31248 28562
rect 31208 28212 31260 28218
rect 31208 28154 31260 28160
rect 31312 28082 31340 28698
rect 31588 28558 31616 28970
rect 31680 28762 31708 29106
rect 31772 28994 31800 30620
rect 31864 30258 31892 30648
rect 31852 30252 31904 30258
rect 31852 30194 31904 30200
rect 32312 30252 32364 30258
rect 32312 30194 32364 30200
rect 31864 29714 31892 30194
rect 31852 29708 31904 29714
rect 31852 29650 31904 29656
rect 32324 29306 32352 30194
rect 32784 30190 32812 30670
rect 33692 30592 33744 30598
rect 33692 30534 33744 30540
rect 33876 30592 33928 30598
rect 33876 30534 33928 30540
rect 32772 30184 32824 30190
rect 32772 30126 32824 30132
rect 32784 29510 32812 30126
rect 33600 29844 33652 29850
rect 33600 29786 33652 29792
rect 33324 29572 33376 29578
rect 33324 29514 33376 29520
rect 32772 29504 32824 29510
rect 32772 29446 32824 29452
rect 33232 29504 33284 29510
rect 33232 29446 33284 29452
rect 32312 29300 32364 29306
rect 32312 29242 32364 29248
rect 32588 29164 32640 29170
rect 32588 29106 32640 29112
rect 32600 29034 32628 29106
rect 32588 29028 32640 29034
rect 31772 28966 31984 28994
rect 32588 28970 32640 28976
rect 31668 28756 31720 28762
rect 31668 28698 31720 28704
rect 31576 28552 31628 28558
rect 31576 28494 31628 28500
rect 31956 28490 31984 28966
rect 32128 28960 32180 28966
rect 32128 28902 32180 28908
rect 32312 28960 32364 28966
rect 32312 28902 32364 28908
rect 32140 28626 32168 28902
rect 32128 28620 32180 28626
rect 32128 28562 32180 28568
rect 32324 28558 32352 28902
rect 32312 28552 32364 28558
rect 32312 28494 32364 28500
rect 31760 28484 31812 28490
rect 31760 28426 31812 28432
rect 31944 28484 31996 28490
rect 31944 28426 31996 28432
rect 31300 28076 31352 28082
rect 31300 28018 31352 28024
rect 31116 27668 31168 27674
rect 31116 27610 31168 27616
rect 30840 27464 30892 27470
rect 30840 27406 30892 27412
rect 30852 26994 30880 27406
rect 31128 27334 31156 27610
rect 31116 27328 31168 27334
rect 31116 27270 31168 27276
rect 30840 26988 30892 26994
rect 30840 26930 30892 26936
rect 31300 26920 31352 26926
rect 31300 26862 31352 26868
rect 31024 26512 31076 26518
rect 31024 26454 31076 26460
rect 31036 25906 31064 26454
rect 31024 25900 31076 25906
rect 31024 25842 31076 25848
rect 30840 25696 30892 25702
rect 30840 25638 30892 25644
rect 30748 25220 30800 25226
rect 30748 25162 30800 25168
rect 30564 25152 30616 25158
rect 30564 25094 30616 25100
rect 30576 24682 30604 25094
rect 30564 24676 30616 24682
rect 30564 24618 30616 24624
rect 30576 24410 30604 24618
rect 30564 24404 30616 24410
rect 30564 24346 30616 24352
rect 30656 24200 30708 24206
rect 30656 24142 30708 24148
rect 30564 24064 30616 24070
rect 30564 24006 30616 24012
rect 30472 23860 30524 23866
rect 30472 23802 30524 23808
rect 30576 23730 30604 24006
rect 30380 23724 30432 23730
rect 30564 23724 30616 23730
rect 30432 23684 30512 23712
rect 30380 23666 30432 23672
rect 29276 23520 29328 23526
rect 29276 23462 29328 23468
rect 29092 21888 29144 21894
rect 29092 21830 29144 21836
rect 28080 21616 28132 21622
rect 28080 21558 28132 21564
rect 28632 21480 28684 21486
rect 28632 21422 28684 21428
rect 27896 21344 27948 21350
rect 27896 21286 27948 21292
rect 27908 21146 27936 21286
rect 28644 21146 28672 21422
rect 27896 21140 27948 21146
rect 27896 21082 27948 21088
rect 28632 21140 28684 21146
rect 28632 21082 28684 21088
rect 28356 19372 28408 19378
rect 28356 19314 28408 19320
rect 28368 18766 28396 19314
rect 28356 18760 28408 18766
rect 28356 18702 28408 18708
rect 27804 18624 27856 18630
rect 27804 18566 27856 18572
rect 27816 18358 27844 18566
rect 27804 18352 27856 18358
rect 27804 18294 27856 18300
rect 27712 18080 27764 18086
rect 27712 18022 27764 18028
rect 28540 18080 28592 18086
rect 28540 18022 28592 18028
rect 28632 18080 28684 18086
rect 28632 18022 28684 18028
rect 27724 17678 27752 18022
rect 28552 17814 28580 18022
rect 28540 17808 28592 17814
rect 28540 17750 28592 17756
rect 27712 17672 27764 17678
rect 27712 17614 27764 17620
rect 28080 17604 28132 17610
rect 28080 17546 28132 17552
rect 27620 17264 27672 17270
rect 27620 17206 27672 17212
rect 28092 17202 28120 17546
rect 28080 17196 28132 17202
rect 28080 17138 28132 17144
rect 28552 17134 28580 17750
rect 28644 17678 28672 18022
rect 28632 17672 28684 17678
rect 28632 17614 28684 17620
rect 28816 17536 28868 17542
rect 28816 17478 28868 17484
rect 28828 17202 28856 17478
rect 28816 17196 28868 17202
rect 28816 17138 28868 17144
rect 28540 17128 28592 17134
rect 28540 17070 28592 17076
rect 27620 17060 27672 17066
rect 27620 17002 27672 17008
rect 27632 16182 27660 17002
rect 27620 16176 27672 16182
rect 27620 16118 27672 16124
rect 28552 16114 28580 17070
rect 27068 16108 27120 16114
rect 26988 16068 27068 16096
rect 26988 15026 27016 16068
rect 27068 16050 27120 16056
rect 27252 16108 27304 16114
rect 27252 16050 27304 16056
rect 28540 16108 28592 16114
rect 28540 16050 28592 16056
rect 27068 15904 27120 15910
rect 27068 15846 27120 15852
rect 27620 15904 27672 15910
rect 27620 15846 27672 15852
rect 26976 15020 27028 15026
rect 26976 14962 27028 14968
rect 27080 14958 27108 15846
rect 27632 15434 27660 15846
rect 27528 15428 27580 15434
rect 27528 15370 27580 15376
rect 27620 15428 27672 15434
rect 27620 15370 27672 15376
rect 27436 15020 27488 15026
rect 27436 14962 27488 14968
rect 27068 14952 27120 14958
rect 27068 14894 27120 14900
rect 26976 14816 27028 14822
rect 26976 14758 27028 14764
rect 26988 14414 27016 14758
rect 27080 14618 27108 14894
rect 27448 14618 27476 14962
rect 27068 14612 27120 14618
rect 27068 14554 27120 14560
rect 27436 14612 27488 14618
rect 27436 14554 27488 14560
rect 26976 14408 27028 14414
rect 26976 14350 27028 14356
rect 27540 13954 27568 15370
rect 28448 14952 28500 14958
rect 28448 14894 28500 14900
rect 28356 14816 28408 14822
rect 28356 14758 28408 14764
rect 27448 13938 27568 13954
rect 28368 13938 28396 14758
rect 27448 13932 27580 13938
rect 27448 13926 27528 13932
rect 27448 12986 27476 13926
rect 27528 13874 27580 13880
rect 28356 13932 28408 13938
rect 28356 13874 28408 13880
rect 27528 13796 27580 13802
rect 27528 13738 27580 13744
rect 27436 12980 27488 12986
rect 27436 12922 27488 12928
rect 27448 12434 27476 12922
rect 27540 12918 27568 13738
rect 27804 13728 27856 13734
rect 27804 13670 27856 13676
rect 27528 12912 27580 12918
rect 27528 12854 27580 12860
rect 27816 12850 27844 13670
rect 27804 12844 27856 12850
rect 27804 12786 27856 12792
rect 27988 12844 28040 12850
rect 27988 12786 28040 12792
rect 27356 12406 27476 12434
rect 27356 12238 27384 12406
rect 27344 12232 27396 12238
rect 27344 12174 27396 12180
rect 26792 11348 26844 11354
rect 26792 11290 26844 11296
rect 27344 11348 27396 11354
rect 27344 11290 27396 11296
rect 27356 10810 27384 11290
rect 27816 11082 27844 12786
rect 28000 12238 28028 12786
rect 28460 12238 28488 14894
rect 29288 13870 29316 23462
rect 30380 23180 30432 23186
rect 30380 23122 30432 23128
rect 30012 23044 30064 23050
rect 30012 22986 30064 22992
rect 29828 22636 29880 22642
rect 29828 22578 29880 22584
rect 29840 21622 29868 22578
rect 30024 22574 30052 22986
rect 30196 22976 30248 22982
rect 30196 22918 30248 22924
rect 30012 22568 30064 22574
rect 30012 22510 30064 22516
rect 30208 22098 30236 22918
rect 30392 22166 30420 23122
rect 30484 22438 30512 23684
rect 30564 23666 30616 23672
rect 30472 22432 30524 22438
rect 30472 22374 30524 22380
rect 30380 22160 30432 22166
rect 30380 22102 30432 22108
rect 30196 22092 30248 22098
rect 30576 22094 30604 23666
rect 30668 23254 30696 24142
rect 30748 24132 30800 24138
rect 30748 24074 30800 24080
rect 30760 23526 30788 24074
rect 30748 23520 30800 23526
rect 30748 23462 30800 23468
rect 30656 23248 30708 23254
rect 30656 23190 30708 23196
rect 30760 22642 30788 23462
rect 30748 22636 30800 22642
rect 30748 22578 30800 22584
rect 30576 22066 30788 22094
rect 30196 22034 30248 22040
rect 30564 21888 30616 21894
rect 30564 21830 30616 21836
rect 29828 21616 29880 21622
rect 29828 21558 29880 21564
rect 30576 21554 30604 21830
rect 30760 21622 30788 22066
rect 30852 21622 30880 25638
rect 31024 25288 31076 25294
rect 31024 25230 31076 25236
rect 31036 24818 31064 25230
rect 31208 25220 31260 25226
rect 31208 25162 31260 25168
rect 31024 24812 31076 24818
rect 31024 24754 31076 24760
rect 31116 24744 31168 24750
rect 31114 24712 31116 24721
rect 31168 24712 31170 24721
rect 31114 24647 31170 24656
rect 30932 23860 30984 23866
rect 30932 23802 30984 23808
rect 30944 23186 30972 23802
rect 31116 23724 31168 23730
rect 31220 23712 31248 25162
rect 31312 24818 31340 26862
rect 31484 26376 31536 26382
rect 31484 26318 31536 26324
rect 31392 25696 31444 25702
rect 31392 25638 31444 25644
rect 31300 24812 31352 24818
rect 31300 24754 31352 24760
rect 31404 24410 31432 25638
rect 31496 25294 31524 26318
rect 31772 25906 31800 28426
rect 32324 28370 32352 28494
rect 32600 28422 32628 28970
rect 32232 28342 32352 28370
rect 32496 28416 32548 28422
rect 32496 28358 32548 28364
rect 32588 28416 32640 28422
rect 32588 28358 32640 28364
rect 31852 27872 31904 27878
rect 31852 27814 31904 27820
rect 31864 27606 31892 27814
rect 31852 27600 31904 27606
rect 31852 27542 31904 27548
rect 31852 27464 31904 27470
rect 31852 27406 31904 27412
rect 32036 27464 32088 27470
rect 32036 27406 32088 27412
rect 31864 26858 31892 27406
rect 31852 26852 31904 26858
rect 31852 26794 31904 26800
rect 31864 26586 31892 26794
rect 31852 26580 31904 26586
rect 31852 26522 31904 26528
rect 32048 26518 32076 27406
rect 32036 26512 32088 26518
rect 32036 26454 32088 26460
rect 32128 26376 32180 26382
rect 32128 26318 32180 26324
rect 31944 26308 31996 26314
rect 31944 26250 31996 26256
rect 31760 25900 31812 25906
rect 31760 25842 31812 25848
rect 31484 25288 31536 25294
rect 31484 25230 31536 25236
rect 31392 24404 31444 24410
rect 31392 24346 31444 24352
rect 31300 24064 31352 24070
rect 31300 24006 31352 24012
rect 31168 23684 31248 23712
rect 31116 23666 31168 23672
rect 30932 23180 30984 23186
rect 30932 23122 30984 23128
rect 31024 23112 31076 23118
rect 31024 23054 31076 23060
rect 30932 22636 30984 22642
rect 30932 22578 30984 22584
rect 30944 21690 30972 22578
rect 31036 22166 31064 23054
rect 31024 22160 31076 22166
rect 31024 22102 31076 22108
rect 30932 21684 30984 21690
rect 30932 21626 30984 21632
rect 30748 21616 30800 21622
rect 30748 21558 30800 21564
rect 30840 21616 30892 21622
rect 30840 21558 30892 21564
rect 29368 21548 29420 21554
rect 29368 21490 29420 21496
rect 30564 21548 30616 21554
rect 30564 21490 30616 21496
rect 29380 21350 29408 21490
rect 30196 21480 30248 21486
rect 30196 21422 30248 21428
rect 29368 21344 29420 21350
rect 29368 21286 29420 21292
rect 29380 20534 29408 21286
rect 30208 21146 30236 21422
rect 30380 21344 30432 21350
rect 30380 21286 30432 21292
rect 30196 21140 30248 21146
rect 30196 21082 30248 21088
rect 30392 20942 30420 21286
rect 30380 20936 30432 20942
rect 30380 20878 30432 20884
rect 29368 20528 29420 20534
rect 29368 20470 29420 20476
rect 29552 20460 29604 20466
rect 29552 20402 29604 20408
rect 29564 19310 29592 20402
rect 30392 19786 30420 20878
rect 30576 20874 30604 21490
rect 30760 20890 30788 21558
rect 30852 21350 30880 21558
rect 30840 21344 30892 21350
rect 30840 21286 30892 21292
rect 30932 21344 30984 21350
rect 30932 21286 30984 21292
rect 30944 20942 30972 21286
rect 31312 20942 31340 24006
rect 31392 23588 31444 23594
rect 31392 23530 31444 23536
rect 31404 23050 31432 23530
rect 31392 23044 31444 23050
rect 31392 22986 31444 22992
rect 31404 22710 31432 22986
rect 31392 22704 31444 22710
rect 31392 22646 31444 22652
rect 31496 22094 31524 25230
rect 31760 25152 31812 25158
rect 31760 25094 31812 25100
rect 31772 24886 31800 25094
rect 31760 24880 31812 24886
rect 31760 24822 31812 24828
rect 31760 24404 31812 24410
rect 31760 24346 31812 24352
rect 31576 24132 31628 24138
rect 31576 24074 31628 24080
rect 31588 23866 31616 24074
rect 31668 24064 31720 24070
rect 31668 24006 31720 24012
rect 31576 23860 31628 23866
rect 31576 23802 31628 23808
rect 31680 23798 31708 24006
rect 31668 23792 31720 23798
rect 31668 23734 31720 23740
rect 31576 23656 31628 23662
rect 31576 23598 31628 23604
rect 31588 23526 31616 23598
rect 31576 23520 31628 23526
rect 31576 23462 31628 23468
rect 31496 22066 31616 22094
rect 31392 21956 31444 21962
rect 31392 21898 31444 21904
rect 31404 21010 31432 21898
rect 31588 21418 31616 22066
rect 31772 21962 31800 24346
rect 31956 23730 31984 26250
rect 32140 25974 32168 26318
rect 32036 25968 32088 25974
rect 32036 25910 32088 25916
rect 32128 25968 32180 25974
rect 32128 25910 32180 25916
rect 32048 25770 32076 25910
rect 32036 25764 32088 25770
rect 32036 25706 32088 25712
rect 32140 25362 32168 25910
rect 32128 25356 32180 25362
rect 32128 25298 32180 25304
rect 32036 24608 32088 24614
rect 32036 24550 32088 24556
rect 32048 24274 32076 24550
rect 32036 24268 32088 24274
rect 32036 24210 32088 24216
rect 32232 24206 32260 28342
rect 32508 27470 32536 28358
rect 32600 28218 32628 28358
rect 32588 28212 32640 28218
rect 32588 28154 32640 28160
rect 32784 28150 32812 29446
rect 33244 29102 33272 29446
rect 33336 29345 33364 29514
rect 33322 29336 33378 29345
rect 33322 29271 33378 29280
rect 33324 29164 33376 29170
rect 33324 29106 33376 29112
rect 33232 29096 33284 29102
rect 33232 29038 33284 29044
rect 32772 28144 32824 28150
rect 32772 28086 32824 28092
rect 32680 28076 32732 28082
rect 32680 28018 32732 28024
rect 32692 27674 32720 28018
rect 32680 27668 32732 27674
rect 32680 27610 32732 27616
rect 32496 27464 32548 27470
rect 32496 27406 32548 27412
rect 32956 27056 33008 27062
rect 32956 26998 33008 27004
rect 32968 26246 32996 26998
rect 32956 26240 33008 26246
rect 32956 26182 33008 26188
rect 33244 25922 33272 29038
rect 33336 28558 33364 29106
rect 33612 28626 33640 29786
rect 33704 29510 33732 30534
rect 33888 30190 33916 30534
rect 34808 30326 34836 31146
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 36004 30734 36032 31726
rect 36636 31680 36688 31686
rect 36636 31622 36688 31628
rect 36648 30734 36676 31622
rect 37568 30938 37596 33050
rect 37556 30932 37608 30938
rect 37556 30874 37608 30880
rect 35992 30728 36044 30734
rect 35992 30670 36044 30676
rect 36636 30728 36688 30734
rect 36636 30670 36688 30676
rect 34796 30320 34848 30326
rect 34796 30262 34848 30268
rect 34520 30252 34572 30258
rect 34520 30194 34572 30200
rect 33876 30184 33928 30190
rect 33876 30126 33928 30132
rect 33888 29578 33916 30126
rect 33968 30048 34020 30054
rect 33968 29990 34020 29996
rect 33876 29572 33928 29578
rect 33876 29514 33928 29520
rect 33692 29504 33744 29510
rect 33692 29446 33744 29452
rect 33704 28966 33732 29446
rect 33888 29170 33916 29514
rect 33980 29170 34008 29990
rect 33876 29164 33928 29170
rect 33876 29106 33928 29112
rect 33968 29164 34020 29170
rect 33968 29106 34020 29112
rect 33980 29034 34008 29106
rect 33968 29028 34020 29034
rect 33968 28970 34020 28976
rect 33692 28960 33744 28966
rect 33692 28902 33744 28908
rect 33600 28620 33652 28626
rect 33600 28562 33652 28568
rect 33324 28552 33376 28558
rect 33324 28494 33376 28500
rect 33336 28218 33364 28494
rect 34532 28490 34560 30194
rect 34808 29646 34836 30262
rect 36004 30122 36032 30670
rect 37464 30252 37516 30258
rect 37464 30194 37516 30200
rect 35992 30116 36044 30122
rect 35992 30058 36044 30064
rect 37188 30116 37240 30122
rect 37188 30058 37240 30064
rect 36820 30048 36872 30054
rect 36820 29990 36872 29996
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 36832 29646 36860 29990
rect 37200 29646 37228 30058
rect 34796 29640 34848 29646
rect 34796 29582 34848 29588
rect 36820 29640 36872 29646
rect 36820 29582 36872 29588
rect 37188 29640 37240 29646
rect 37188 29582 37240 29588
rect 35624 29572 35676 29578
rect 35624 29514 35676 29520
rect 35532 29164 35584 29170
rect 35532 29106 35584 29112
rect 34796 29028 34848 29034
rect 34796 28970 34848 28976
rect 34808 28626 34836 28970
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 35544 28762 35572 29106
rect 35532 28756 35584 28762
rect 35532 28698 35584 28704
rect 34888 28688 34940 28694
rect 34888 28630 34940 28636
rect 34796 28620 34848 28626
rect 34796 28562 34848 28568
rect 34520 28484 34572 28490
rect 34520 28426 34572 28432
rect 34428 28416 34480 28422
rect 34428 28358 34480 28364
rect 33324 28212 33376 28218
rect 33324 28154 33376 28160
rect 34060 28144 34112 28150
rect 34060 28086 34112 28092
rect 33600 28008 33652 28014
rect 33600 27950 33652 27956
rect 33508 27328 33560 27334
rect 33508 27270 33560 27276
rect 33324 26444 33376 26450
rect 33324 26386 33376 26392
rect 33336 26246 33364 26386
rect 33324 26240 33376 26246
rect 33324 26182 33376 26188
rect 33060 25894 33272 25922
rect 33336 25906 33364 26182
rect 33324 25900 33376 25906
rect 33060 25838 33088 25894
rect 33324 25842 33376 25848
rect 33048 25832 33100 25838
rect 33048 25774 33100 25780
rect 32312 24812 32364 24818
rect 32364 24772 32444 24800
rect 32312 24754 32364 24760
rect 32416 24682 32444 24772
rect 32404 24676 32456 24682
rect 32404 24618 32456 24624
rect 32312 24608 32364 24614
rect 32312 24550 32364 24556
rect 32220 24200 32272 24206
rect 32220 24142 32272 24148
rect 31944 23724 31996 23730
rect 31944 23666 31996 23672
rect 31944 22636 31996 22642
rect 31944 22578 31996 22584
rect 31956 22098 31984 22578
rect 31944 22092 31996 22098
rect 31944 22034 31996 22040
rect 31956 21962 31984 22034
rect 31760 21956 31812 21962
rect 31760 21898 31812 21904
rect 31944 21956 31996 21962
rect 31944 21898 31996 21904
rect 31668 21888 31720 21894
rect 31668 21830 31720 21836
rect 31680 21622 31708 21830
rect 31668 21616 31720 21622
rect 31668 21558 31720 21564
rect 31944 21548 31996 21554
rect 31944 21490 31996 21496
rect 31576 21412 31628 21418
rect 31576 21354 31628 21360
rect 31956 21146 31984 21490
rect 32324 21486 32352 24550
rect 32416 23730 32444 24618
rect 32956 24608 33008 24614
rect 32956 24550 33008 24556
rect 32968 24410 32996 24550
rect 32956 24404 33008 24410
rect 32956 24346 33008 24352
rect 32404 23724 32456 23730
rect 32404 23666 32456 23672
rect 33324 23656 33376 23662
rect 33324 23598 33376 23604
rect 33336 22778 33364 23598
rect 33416 23520 33468 23526
rect 33416 23462 33468 23468
rect 33428 23118 33456 23462
rect 33416 23112 33468 23118
rect 33416 23054 33468 23060
rect 33324 22772 33376 22778
rect 33324 22714 33376 22720
rect 33140 22500 33192 22506
rect 33140 22442 33192 22448
rect 32772 22432 32824 22438
rect 32772 22374 32824 22380
rect 32784 22030 32812 22374
rect 32496 22024 32548 22030
rect 32496 21966 32548 21972
rect 32772 22024 32824 22030
rect 32772 21966 32824 21972
rect 32508 21690 32536 21966
rect 32680 21888 32732 21894
rect 32680 21830 32732 21836
rect 32496 21684 32548 21690
rect 32496 21626 32548 21632
rect 32312 21480 32364 21486
rect 32312 21422 32364 21428
rect 31944 21140 31996 21146
rect 31944 21082 31996 21088
rect 31392 21004 31444 21010
rect 31392 20946 31444 20952
rect 30932 20936 30984 20942
rect 30564 20868 30616 20874
rect 30760 20862 30880 20890
rect 31300 20936 31352 20942
rect 30932 20878 30984 20884
rect 31220 20896 31300 20924
rect 30564 20810 30616 20816
rect 30576 20466 30604 20810
rect 30852 20806 30880 20862
rect 30748 20800 30800 20806
rect 30748 20742 30800 20748
rect 30840 20800 30892 20806
rect 30840 20742 30892 20748
rect 30564 20460 30616 20466
rect 30564 20402 30616 20408
rect 30576 19854 30604 20402
rect 30564 19848 30616 19854
rect 30564 19790 30616 19796
rect 30380 19780 30432 19786
rect 30380 19722 30432 19728
rect 29552 19304 29604 19310
rect 29552 19246 29604 19252
rect 29564 18698 29592 19246
rect 29460 18692 29512 18698
rect 29460 18634 29512 18640
rect 29552 18692 29604 18698
rect 29552 18634 29604 18640
rect 30564 18692 30616 18698
rect 30564 18634 30616 18640
rect 29472 17610 29500 18634
rect 29564 17746 29592 18634
rect 30196 18284 30248 18290
rect 30196 18226 30248 18232
rect 29552 17740 29604 17746
rect 29552 17682 29604 17688
rect 29460 17604 29512 17610
rect 29460 17546 29512 17552
rect 29472 17270 29500 17546
rect 30208 17338 30236 18226
rect 30472 18216 30524 18222
rect 30472 18158 30524 18164
rect 30484 17882 30512 18158
rect 30472 17876 30524 17882
rect 30472 17818 30524 17824
rect 30576 17610 30604 18634
rect 30656 18080 30708 18086
rect 30656 18022 30708 18028
rect 30564 17604 30616 17610
rect 30564 17546 30616 17552
rect 30576 17338 30604 17546
rect 29644 17332 29696 17338
rect 29644 17274 29696 17280
rect 30196 17332 30248 17338
rect 30196 17274 30248 17280
rect 30564 17332 30616 17338
rect 30564 17274 30616 17280
rect 29460 17264 29512 17270
rect 29460 17206 29512 17212
rect 29552 15904 29604 15910
rect 29552 15846 29604 15852
rect 29564 15162 29592 15846
rect 29656 15502 29684 17274
rect 29736 17196 29788 17202
rect 29736 17138 29788 17144
rect 29644 15496 29696 15502
rect 29644 15438 29696 15444
rect 29748 15366 29776 17138
rect 29920 15904 29972 15910
rect 29920 15846 29972 15852
rect 29736 15360 29788 15366
rect 29736 15302 29788 15308
rect 29552 15156 29604 15162
rect 29552 15098 29604 15104
rect 29644 14340 29696 14346
rect 29644 14282 29696 14288
rect 29656 14074 29684 14282
rect 29644 14068 29696 14074
rect 29644 14010 29696 14016
rect 29748 14006 29776 15302
rect 29932 14482 29960 15846
rect 30196 14884 30248 14890
rect 30196 14826 30248 14832
rect 30012 14816 30064 14822
rect 30012 14758 30064 14764
rect 30024 14618 30052 14758
rect 30208 14618 30236 14826
rect 30668 14822 30696 18022
rect 30760 16590 30788 20742
rect 30944 19446 30972 20878
rect 31220 20466 31248 20896
rect 31300 20878 31352 20884
rect 31668 20936 31720 20942
rect 31668 20878 31720 20884
rect 31680 20466 31708 20878
rect 32324 20466 32352 21422
rect 32496 20528 32548 20534
rect 32496 20470 32548 20476
rect 31208 20460 31260 20466
rect 31208 20402 31260 20408
rect 31300 20460 31352 20466
rect 31300 20402 31352 20408
rect 31576 20460 31628 20466
rect 31576 20402 31628 20408
rect 31668 20460 31720 20466
rect 31668 20402 31720 20408
rect 32312 20460 32364 20466
rect 32312 20402 32364 20408
rect 31208 20256 31260 20262
rect 31208 20198 31260 20204
rect 30932 19440 30984 19446
rect 30932 19382 30984 19388
rect 31024 17536 31076 17542
rect 31024 17478 31076 17484
rect 31036 16658 31064 17478
rect 31024 16652 31076 16658
rect 31024 16594 31076 16600
rect 30748 16584 30800 16590
rect 30748 16526 30800 16532
rect 31036 15502 31064 16594
rect 31220 15502 31248 20198
rect 31312 18766 31340 20402
rect 31588 20058 31616 20402
rect 31576 20052 31628 20058
rect 31576 19994 31628 20000
rect 32508 19922 32536 20470
rect 32496 19916 32548 19922
rect 32496 19858 32548 19864
rect 32692 19854 32720 21830
rect 33048 21412 33100 21418
rect 33048 21354 33100 21360
rect 33060 20806 33088 21354
rect 33152 21146 33180 22442
rect 33520 22438 33548 27270
rect 33612 26994 33640 27950
rect 33600 26988 33652 26994
rect 33600 26930 33652 26936
rect 33968 26988 34020 26994
rect 33968 26930 34020 26936
rect 33600 26376 33652 26382
rect 33600 26318 33652 26324
rect 33784 26376 33836 26382
rect 33784 26318 33836 26324
rect 33612 25974 33640 26318
rect 33796 26042 33824 26318
rect 33876 26240 33928 26246
rect 33876 26182 33928 26188
rect 33784 26036 33836 26042
rect 33784 25978 33836 25984
rect 33600 25968 33652 25974
rect 33600 25910 33652 25916
rect 33888 25294 33916 26182
rect 33980 25906 34008 26930
rect 33968 25900 34020 25906
rect 33968 25842 34020 25848
rect 34072 25294 34100 28086
rect 34440 28082 34468 28358
rect 34428 28076 34480 28082
rect 34428 28018 34480 28024
rect 34900 27962 34928 28630
rect 35532 28484 35584 28490
rect 35532 28426 35584 28432
rect 35544 28082 35572 28426
rect 35532 28076 35584 28082
rect 35532 28018 35584 28024
rect 34808 27934 34928 27962
rect 34704 27464 34756 27470
rect 34704 27406 34756 27412
rect 34612 27396 34664 27402
rect 34612 27338 34664 27344
rect 34428 27328 34480 27334
rect 34428 27270 34480 27276
rect 34152 27056 34204 27062
rect 34152 26998 34204 27004
rect 34164 25906 34192 26998
rect 34440 26994 34468 27270
rect 34624 26994 34652 27338
rect 34716 27062 34744 27406
rect 34704 27056 34756 27062
rect 34704 26998 34756 27004
rect 34244 26988 34296 26994
rect 34244 26930 34296 26936
rect 34428 26988 34480 26994
rect 34428 26930 34480 26936
rect 34612 26988 34664 26994
rect 34612 26930 34664 26936
rect 34256 26314 34284 26930
rect 34624 26586 34652 26930
rect 34612 26580 34664 26586
rect 34612 26522 34664 26528
rect 34704 26580 34756 26586
rect 34704 26522 34756 26528
rect 34520 26376 34572 26382
rect 34520 26318 34572 26324
rect 34244 26308 34296 26314
rect 34244 26250 34296 26256
rect 34532 25906 34560 26318
rect 34624 25974 34652 26522
rect 34716 26042 34744 26522
rect 34704 26036 34756 26042
rect 34704 25978 34756 25984
rect 34612 25968 34664 25974
rect 34612 25910 34664 25916
rect 34152 25900 34204 25906
rect 34152 25842 34204 25848
rect 34520 25900 34572 25906
rect 34520 25842 34572 25848
rect 33876 25288 33928 25294
rect 33876 25230 33928 25236
rect 34060 25288 34112 25294
rect 34060 25230 34112 25236
rect 34072 23730 34100 25230
rect 34060 23724 34112 23730
rect 34060 23666 34112 23672
rect 34152 23724 34204 23730
rect 34152 23666 34204 23672
rect 33968 23656 34020 23662
rect 33968 23598 34020 23604
rect 33876 23588 33928 23594
rect 33876 23530 33928 23536
rect 33888 23118 33916 23530
rect 33876 23112 33928 23118
rect 33876 23054 33928 23060
rect 33980 22982 34008 23598
rect 34164 23322 34192 23666
rect 34152 23316 34204 23322
rect 34152 23258 34204 23264
rect 34428 23112 34480 23118
rect 34428 23054 34480 23060
rect 33968 22976 34020 22982
rect 33968 22918 34020 22924
rect 33980 22574 34008 22918
rect 34336 22636 34388 22642
rect 34336 22578 34388 22584
rect 34440 22624 34468 23054
rect 34612 22636 34664 22642
rect 34440 22596 34612 22624
rect 33968 22568 34020 22574
rect 33968 22510 34020 22516
rect 33784 22500 33836 22506
rect 33784 22442 33836 22448
rect 33508 22432 33560 22438
rect 33508 22374 33560 22380
rect 33796 22166 33824 22442
rect 33980 22234 34008 22510
rect 33968 22228 34020 22234
rect 33968 22170 34020 22176
rect 33784 22160 33836 22166
rect 33784 22102 33836 22108
rect 34348 21962 34376 22578
rect 34336 21956 34388 21962
rect 34336 21898 34388 21904
rect 34348 21690 34376 21898
rect 34440 21894 34468 22596
rect 34612 22578 34664 22584
rect 34808 22506 34836 27934
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 35348 26784 35400 26790
rect 35348 26726 35400 26732
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 35360 26518 35388 26726
rect 35348 26512 35400 26518
rect 35348 26454 35400 26460
rect 35360 25906 35388 26454
rect 35348 25900 35400 25906
rect 35348 25842 35400 25848
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 35532 23656 35584 23662
rect 35532 23598 35584 23604
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 35544 22574 35572 23598
rect 35532 22568 35584 22574
rect 35532 22510 35584 22516
rect 34796 22500 34848 22506
rect 34796 22442 34848 22448
rect 34704 22432 34756 22438
rect 34704 22374 34756 22380
rect 34716 22030 34744 22374
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 35544 22030 35572 22510
rect 34704 22024 34756 22030
rect 34704 21966 34756 21972
rect 35532 22024 35584 22030
rect 35532 21966 35584 21972
rect 34428 21888 34480 21894
rect 34428 21830 34480 21836
rect 34796 21888 34848 21894
rect 34796 21830 34848 21836
rect 34336 21684 34388 21690
rect 34336 21626 34388 21632
rect 34808 21622 34836 21830
rect 34796 21616 34848 21622
rect 34796 21558 34848 21564
rect 35348 21480 35400 21486
rect 35348 21422 35400 21428
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 33140 21140 33192 21146
rect 33140 21082 33192 21088
rect 33416 20868 33468 20874
rect 33416 20810 33468 20816
rect 33048 20800 33100 20806
rect 33048 20742 33100 20748
rect 33324 20460 33376 20466
rect 33324 20402 33376 20408
rect 32956 19916 33008 19922
rect 32956 19858 33008 19864
rect 32680 19848 32732 19854
rect 32680 19790 32732 19796
rect 32968 19446 32996 19858
rect 32956 19440 33008 19446
rect 32956 19382 33008 19388
rect 33336 19378 33364 20402
rect 33428 20398 33456 20810
rect 35256 20800 35308 20806
rect 35256 20742 35308 20748
rect 33416 20392 33468 20398
rect 33416 20334 33468 20340
rect 35268 20330 35296 20742
rect 35360 20534 35388 21422
rect 35440 21344 35492 21350
rect 35440 21286 35492 21292
rect 35452 21010 35480 21286
rect 35440 21004 35492 21010
rect 35440 20946 35492 20952
rect 35348 20528 35400 20534
rect 35348 20470 35400 20476
rect 35256 20324 35308 20330
rect 35256 20266 35308 20272
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 35360 19922 35388 20470
rect 35348 19916 35400 19922
rect 35348 19858 35400 19864
rect 33324 19372 33376 19378
rect 33324 19314 33376 19320
rect 31576 19168 31628 19174
rect 31576 19110 31628 19116
rect 31300 18760 31352 18766
rect 31300 18702 31352 18708
rect 31024 15496 31076 15502
rect 31024 15438 31076 15444
rect 31208 15496 31260 15502
rect 31208 15438 31260 15444
rect 30840 15088 30892 15094
rect 30840 15030 30892 15036
rect 30656 14816 30708 14822
rect 30656 14758 30708 14764
rect 30012 14612 30064 14618
rect 30012 14554 30064 14560
rect 30196 14612 30248 14618
rect 30196 14554 30248 14560
rect 29920 14476 29972 14482
rect 29920 14418 29972 14424
rect 30196 14476 30248 14482
rect 30196 14418 30248 14424
rect 30104 14408 30156 14414
rect 30104 14350 30156 14356
rect 30116 14074 30144 14350
rect 30104 14068 30156 14074
rect 30104 14010 30156 14016
rect 29736 14000 29788 14006
rect 29736 13942 29788 13948
rect 30208 13938 30236 14418
rect 30196 13932 30248 13938
rect 30196 13874 30248 13880
rect 29276 13864 29328 13870
rect 29276 13806 29328 13812
rect 29828 12844 29880 12850
rect 29828 12786 29880 12792
rect 28816 12640 28868 12646
rect 28816 12582 28868 12588
rect 27988 12232 28040 12238
rect 27988 12174 28040 12180
rect 28448 12232 28500 12238
rect 28448 12174 28500 12180
rect 28000 11218 28028 12174
rect 28460 11762 28488 12174
rect 28828 11830 28856 12582
rect 29840 11898 29868 12786
rect 30472 12640 30524 12646
rect 30472 12582 30524 12588
rect 30484 12170 30512 12582
rect 30852 12434 30880 15030
rect 31588 14414 31616 19110
rect 32588 18624 32640 18630
rect 32588 18566 32640 18572
rect 32600 18290 32628 18566
rect 32588 18284 32640 18290
rect 32588 18226 32640 18232
rect 33140 18284 33192 18290
rect 33140 18226 33192 18232
rect 32600 17746 32628 18226
rect 33152 17882 33180 18226
rect 33232 18216 33284 18222
rect 33232 18158 33284 18164
rect 33140 17876 33192 17882
rect 33140 17818 33192 17824
rect 32588 17740 32640 17746
rect 32588 17682 32640 17688
rect 33152 17610 33180 17818
rect 33244 17678 33272 18158
rect 33336 17814 33364 19314
rect 34704 19168 34756 19174
rect 34704 19110 34756 19116
rect 34612 18828 34664 18834
rect 34612 18770 34664 18776
rect 34428 18692 34480 18698
rect 34428 18634 34480 18640
rect 34440 18358 34468 18634
rect 34428 18352 34480 18358
rect 34428 18294 34480 18300
rect 34520 18284 34572 18290
rect 34520 18226 34572 18232
rect 33324 17808 33376 17814
rect 33324 17750 33376 17756
rect 34532 17746 34560 18226
rect 34520 17740 34572 17746
rect 34520 17682 34572 17688
rect 34624 17678 34652 18770
rect 34716 18766 34744 19110
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 34980 18828 35032 18834
rect 34980 18770 35032 18776
rect 35256 18828 35308 18834
rect 35256 18770 35308 18776
rect 34704 18760 34756 18766
rect 34704 18702 34756 18708
rect 34888 18760 34940 18766
rect 34888 18702 34940 18708
rect 34900 18358 34928 18702
rect 34888 18352 34940 18358
rect 34808 18300 34888 18306
rect 34808 18294 34940 18300
rect 34704 18284 34756 18290
rect 34704 18226 34756 18232
rect 34808 18278 34928 18294
rect 34992 18290 35020 18770
rect 34980 18284 35032 18290
rect 34716 17882 34744 18226
rect 34704 17876 34756 17882
rect 34704 17818 34756 17824
rect 34808 17746 34836 18278
rect 34980 18226 35032 18232
rect 35268 18222 35296 18770
rect 35256 18216 35308 18222
rect 35256 18158 35308 18164
rect 35348 18080 35400 18086
rect 35348 18022 35400 18028
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 34796 17740 34848 17746
rect 34796 17682 34848 17688
rect 35360 17678 35388 18022
rect 33232 17672 33284 17678
rect 33232 17614 33284 17620
rect 34612 17672 34664 17678
rect 34612 17614 34664 17620
rect 34888 17672 34940 17678
rect 34888 17614 34940 17620
rect 35348 17672 35400 17678
rect 35348 17614 35400 17620
rect 33140 17604 33192 17610
rect 33140 17546 33192 17552
rect 34900 17270 34928 17614
rect 35348 17536 35400 17542
rect 35348 17478 35400 17484
rect 34888 17264 34940 17270
rect 34888 17206 34940 17212
rect 32864 17196 32916 17202
rect 32864 17138 32916 17144
rect 33048 17196 33100 17202
rect 33048 17138 33100 17144
rect 32876 16182 32904 17138
rect 33060 16726 33088 17138
rect 33784 16992 33836 16998
rect 33784 16934 33836 16940
rect 33048 16720 33100 16726
rect 33048 16662 33100 16668
rect 32956 16516 33008 16522
rect 32956 16458 33008 16464
rect 32968 16250 32996 16458
rect 32956 16244 33008 16250
rect 32956 16186 33008 16192
rect 33060 16182 33088 16662
rect 33796 16658 33824 16934
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 35360 16658 35388 17478
rect 33784 16652 33836 16658
rect 33784 16594 33836 16600
rect 34060 16652 34112 16658
rect 34060 16594 34112 16600
rect 35348 16652 35400 16658
rect 35348 16594 35400 16600
rect 33232 16448 33284 16454
rect 33232 16390 33284 16396
rect 33244 16250 33272 16390
rect 33232 16244 33284 16250
rect 33232 16186 33284 16192
rect 32864 16176 32916 16182
rect 32864 16118 32916 16124
rect 33048 16176 33100 16182
rect 33048 16118 33100 16124
rect 33796 16114 33824 16594
rect 33784 16108 33836 16114
rect 33784 16050 33836 16056
rect 32956 15496 33008 15502
rect 32956 15438 33008 15444
rect 33232 15496 33284 15502
rect 33232 15438 33284 15444
rect 32312 15360 32364 15366
rect 32312 15302 32364 15308
rect 32220 14884 32272 14890
rect 32220 14826 32272 14832
rect 31576 14408 31628 14414
rect 31576 14350 31628 14356
rect 32232 13938 32260 14826
rect 32324 13938 32352 15302
rect 32968 14890 32996 15438
rect 33140 15360 33192 15366
rect 33140 15302 33192 15308
rect 33152 15026 33180 15302
rect 33244 15094 33272 15438
rect 33600 15360 33652 15366
rect 33600 15302 33652 15308
rect 33232 15088 33284 15094
rect 33232 15030 33284 15036
rect 33140 15020 33192 15026
rect 33140 14962 33192 14968
rect 32956 14884 33008 14890
rect 32956 14826 33008 14832
rect 32404 14816 32456 14822
rect 32404 14758 32456 14764
rect 32416 14414 32444 14758
rect 32404 14408 32456 14414
rect 32404 14350 32456 14356
rect 33244 14074 33272 15030
rect 33612 15026 33640 15302
rect 34072 15026 34100 16594
rect 34888 16584 34940 16590
rect 34888 16526 34940 16532
rect 34900 16250 34928 16526
rect 34888 16244 34940 16250
rect 34888 16186 34940 16192
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 33600 15020 33652 15026
rect 33600 14962 33652 14968
rect 34060 15020 34112 15026
rect 34060 14962 34112 14968
rect 35532 14952 35584 14958
rect 35532 14894 35584 14900
rect 34428 14816 34480 14822
rect 34428 14758 34480 14764
rect 35348 14816 35400 14822
rect 35348 14758 35400 14764
rect 33508 14272 33560 14278
rect 33508 14214 33560 14220
rect 34336 14272 34388 14278
rect 34336 14214 34388 14220
rect 33232 14068 33284 14074
rect 33232 14010 33284 14016
rect 32220 13932 32272 13938
rect 32220 13874 32272 13880
rect 32312 13932 32364 13938
rect 32312 13874 32364 13880
rect 33520 13870 33548 14214
rect 34348 14074 34376 14214
rect 34440 14074 34468 14758
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 35360 14414 35388 14758
rect 35544 14482 35572 14894
rect 35532 14476 35584 14482
rect 35532 14418 35584 14424
rect 35348 14408 35400 14414
rect 35348 14350 35400 14356
rect 35544 14226 35572 14418
rect 35360 14198 35572 14226
rect 34336 14068 34388 14074
rect 34336 14010 34388 14016
rect 34428 14068 34480 14074
rect 34428 14010 34480 14016
rect 31484 13864 31536 13870
rect 31484 13806 31536 13812
rect 33508 13864 33560 13870
rect 33508 13806 33560 13812
rect 34428 13864 34480 13870
rect 34428 13806 34480 13812
rect 31496 12918 31524 13806
rect 33968 13728 34020 13734
rect 33968 13670 34020 13676
rect 33980 13326 34008 13670
rect 33968 13320 34020 13326
rect 33968 13262 34020 13268
rect 32680 13184 32732 13190
rect 32680 13126 32732 13132
rect 31116 12912 31168 12918
rect 31116 12854 31168 12860
rect 31484 12912 31536 12918
rect 31484 12854 31536 12860
rect 30760 12406 30880 12434
rect 30472 12164 30524 12170
rect 30472 12106 30524 12112
rect 30760 11898 30788 12406
rect 31128 12238 31156 12854
rect 32692 12850 32720 13126
rect 32680 12844 32732 12850
rect 32680 12786 32732 12792
rect 33508 12844 33560 12850
rect 33508 12786 33560 12792
rect 32128 12640 32180 12646
rect 32128 12582 32180 12588
rect 32140 12306 32168 12582
rect 32128 12300 32180 12306
rect 32128 12242 32180 12248
rect 32312 12300 32364 12306
rect 32312 12242 32364 12248
rect 31116 12232 31168 12238
rect 31116 12174 31168 12180
rect 31024 12096 31076 12102
rect 31024 12038 31076 12044
rect 31208 12096 31260 12102
rect 31208 12038 31260 12044
rect 32128 12096 32180 12102
rect 32128 12038 32180 12044
rect 29828 11892 29880 11898
rect 29828 11834 29880 11840
rect 30748 11892 30800 11898
rect 30748 11834 30800 11840
rect 28816 11824 28868 11830
rect 28816 11766 28868 11772
rect 31036 11762 31064 12038
rect 31220 11898 31248 12038
rect 32140 11898 32168 12038
rect 31208 11892 31260 11898
rect 31208 11834 31260 11840
rect 32128 11892 32180 11898
rect 32128 11834 32180 11840
rect 28448 11756 28500 11762
rect 28448 11698 28500 11704
rect 31024 11756 31076 11762
rect 31024 11698 31076 11704
rect 27988 11212 28040 11218
rect 27988 11154 28040 11160
rect 27620 11076 27672 11082
rect 27620 11018 27672 11024
rect 27804 11076 27856 11082
rect 27804 11018 27856 11024
rect 27344 10804 27396 10810
rect 27344 10746 27396 10752
rect 27632 9994 27660 11018
rect 28172 11008 28224 11014
rect 28172 10950 28224 10956
rect 28184 10674 28212 10950
rect 28460 10674 28488 11698
rect 31300 11688 31352 11694
rect 31300 11630 31352 11636
rect 31312 11354 31340 11630
rect 31300 11348 31352 11354
rect 31300 11290 31352 11296
rect 30196 11144 30248 11150
rect 30196 11086 30248 11092
rect 30208 10810 30236 11086
rect 32324 11082 32352 12242
rect 33324 12232 33376 12238
rect 33324 12174 33376 12180
rect 33140 12096 33192 12102
rect 33140 12038 33192 12044
rect 33152 11830 33180 12038
rect 33336 11898 33364 12174
rect 33324 11892 33376 11898
rect 33324 11834 33376 11840
rect 33140 11824 33192 11830
rect 33140 11766 33192 11772
rect 33520 11762 33548 12786
rect 34440 12782 34468 13806
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 34428 12776 34480 12782
rect 34428 12718 34480 12724
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 35360 12306 35388 14198
rect 35440 12640 35492 12646
rect 35440 12582 35492 12588
rect 35348 12300 35400 12306
rect 35348 12242 35400 12248
rect 33784 12096 33836 12102
rect 33784 12038 33836 12044
rect 33508 11756 33560 11762
rect 33508 11698 33560 11704
rect 33520 11150 33548 11698
rect 33508 11144 33560 11150
rect 33508 11086 33560 11092
rect 33796 11082 33824 12038
rect 34704 11756 34756 11762
rect 34704 11698 34756 11704
rect 34716 11354 34744 11698
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 34704 11348 34756 11354
rect 34704 11290 34756 11296
rect 35360 11150 35388 12242
rect 35452 12238 35480 12582
rect 35440 12232 35492 12238
rect 35440 12174 35492 12180
rect 35532 12096 35584 12102
rect 35532 12038 35584 12044
rect 35544 11898 35572 12038
rect 35532 11892 35584 11898
rect 35532 11834 35584 11840
rect 35348 11144 35400 11150
rect 35348 11086 35400 11092
rect 32312 11076 32364 11082
rect 32312 11018 32364 11024
rect 33784 11076 33836 11082
rect 33784 11018 33836 11024
rect 30840 11008 30892 11014
rect 30840 10950 30892 10956
rect 30196 10804 30248 10810
rect 30196 10746 30248 10752
rect 28172 10668 28224 10674
rect 28172 10610 28224 10616
rect 28448 10668 28500 10674
rect 28448 10610 28500 10616
rect 28460 10130 28488 10610
rect 28448 10124 28500 10130
rect 28448 10066 28500 10072
rect 30852 10062 30880 10950
rect 32324 10266 32352 11018
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 32312 10260 32364 10266
rect 32312 10202 32364 10208
rect 30840 10056 30892 10062
rect 30840 9998 30892 10004
rect 27620 9988 27672 9994
rect 27620 9930 27672 9936
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 26332 7744 26384 7750
rect 26332 7686 26384 7692
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 35636 6914 35664 29514
rect 35808 29504 35860 29510
rect 35808 29446 35860 29452
rect 35820 29170 35848 29446
rect 35990 29336 36046 29345
rect 35990 29271 36046 29280
rect 36004 29238 36032 29271
rect 35992 29232 36044 29238
rect 35992 29174 36044 29180
rect 35808 29164 35860 29170
rect 35808 29106 35860 29112
rect 35716 28960 35768 28966
rect 35716 28902 35768 28908
rect 36544 28960 36596 28966
rect 36544 28902 36596 28908
rect 35728 28762 35756 28902
rect 35716 28756 35768 28762
rect 35716 28698 35768 28704
rect 36556 28490 36584 28902
rect 37200 28558 37228 29582
rect 37476 28762 37504 30194
rect 37464 28756 37516 28762
rect 37464 28698 37516 28704
rect 37188 28552 37240 28558
rect 37188 28494 37240 28500
rect 36084 28484 36136 28490
rect 36084 28426 36136 28432
rect 36544 28484 36596 28490
rect 36544 28426 36596 28432
rect 36728 28484 36780 28490
rect 36728 28426 36780 28432
rect 36096 28218 36124 28426
rect 36176 28416 36228 28422
rect 36176 28358 36228 28364
rect 36084 28212 36136 28218
rect 36084 28154 36136 28160
rect 36096 27470 36124 28154
rect 36188 27878 36216 28358
rect 36740 28218 36768 28426
rect 36728 28212 36780 28218
rect 36728 28154 36780 28160
rect 36268 28076 36320 28082
rect 36268 28018 36320 28024
rect 36176 27872 36228 27878
rect 36176 27814 36228 27820
rect 36188 27470 36216 27814
rect 36280 27674 36308 28018
rect 36268 27668 36320 27674
rect 36268 27610 36320 27616
rect 36084 27464 36136 27470
rect 36084 27406 36136 27412
rect 36176 27464 36228 27470
rect 36176 27406 36228 27412
rect 35992 26308 36044 26314
rect 35992 26250 36044 26256
rect 35716 26240 35768 26246
rect 35716 26182 35768 26188
rect 35728 25906 35756 26182
rect 36004 26042 36032 26250
rect 35992 26036 36044 26042
rect 35992 25978 36044 25984
rect 35716 25900 35768 25906
rect 35716 25842 35768 25848
rect 35900 24064 35952 24070
rect 35900 24006 35952 24012
rect 35912 23254 35940 24006
rect 35900 23248 35952 23254
rect 35900 23190 35952 23196
rect 35912 22710 35940 23190
rect 35900 22704 35952 22710
rect 35952 22664 36032 22692
rect 35900 22646 35952 22652
rect 35900 22568 35952 22574
rect 35900 22510 35952 22516
rect 35808 22024 35860 22030
rect 35912 22012 35940 22510
rect 36004 22030 36032 22664
rect 36188 22094 36216 27406
rect 37200 26926 37228 28494
rect 37464 28416 37516 28422
rect 37464 28358 37516 28364
rect 37476 28082 37504 28358
rect 37464 28076 37516 28082
rect 37464 28018 37516 28024
rect 37188 26920 37240 26926
rect 37188 26862 37240 26868
rect 37200 26382 37228 26862
rect 37188 26376 37240 26382
rect 37188 26318 37240 26324
rect 37200 25838 37228 26318
rect 37372 25900 37424 25906
rect 37372 25842 37424 25848
rect 37188 25832 37240 25838
rect 37188 25774 37240 25780
rect 37200 24886 37228 25774
rect 37188 24880 37240 24886
rect 37188 24822 37240 24828
rect 37200 24206 37228 24822
rect 37188 24200 37240 24206
rect 37188 24142 37240 24148
rect 37384 23730 37412 25842
rect 37832 24200 37884 24206
rect 37832 24142 37884 24148
rect 37844 23866 37872 24142
rect 37832 23860 37884 23866
rect 37832 23802 37884 23808
rect 36360 23724 36412 23730
rect 36360 23666 36412 23672
rect 37372 23724 37424 23730
rect 37372 23666 37424 23672
rect 36372 23118 36400 23666
rect 36360 23112 36412 23118
rect 36360 23054 36412 23060
rect 37384 23050 37412 23666
rect 37844 23186 37872 23802
rect 37832 23180 37884 23186
rect 37832 23122 37884 23128
rect 37648 23112 37700 23118
rect 37648 23054 37700 23060
rect 37372 23044 37424 23050
rect 37372 22986 37424 22992
rect 37660 22642 37688 23054
rect 37648 22636 37700 22642
rect 37648 22578 37700 22584
rect 36096 22066 36216 22094
rect 35860 21984 35940 22012
rect 35992 22024 36044 22030
rect 35808 21966 35860 21972
rect 35992 21966 36044 21972
rect 36096 21690 36124 22066
rect 37660 22030 37688 22578
rect 37648 22024 37700 22030
rect 37648 21966 37700 21972
rect 36176 21888 36228 21894
rect 36176 21830 36228 21836
rect 36084 21684 36136 21690
rect 36084 21626 36136 21632
rect 36188 21554 36216 21830
rect 36176 21548 36228 21554
rect 36176 21490 36228 21496
rect 35900 21480 35952 21486
rect 35900 21422 35952 21428
rect 35912 21078 35940 21422
rect 35900 21072 35952 21078
rect 35900 21014 35952 21020
rect 37936 20602 37964 41550
rect 39868 41274 39896 41550
rect 41510 41511 41566 41520
rect 39856 41268 39908 41274
rect 39856 41210 39908 41216
rect 41524 41070 41552 41511
rect 42168 41414 42196 45070
rect 42522 44976 42578 44985
rect 42522 44911 42578 44920
rect 42536 41682 42564 44911
rect 42892 43104 42944 43110
rect 42892 43046 42944 43052
rect 42904 42770 42932 43046
rect 43824 42770 43852 45200
rect 44180 43104 44232 43110
rect 44180 43046 44232 43052
rect 42892 42764 42944 42770
rect 42892 42706 42944 42712
rect 43812 42764 43864 42770
rect 43812 42706 43864 42712
rect 42708 42628 42760 42634
rect 42708 42570 42760 42576
rect 42720 42362 42748 42570
rect 42708 42356 42760 42362
rect 42708 42298 42760 42304
rect 42616 42288 42668 42294
rect 42614 42256 42616 42265
rect 42668 42256 42670 42265
rect 42614 42191 42670 42200
rect 42800 42220 42852 42226
rect 42800 42162 42852 42168
rect 43536 42220 43588 42226
rect 43536 42162 43588 42168
rect 43904 42220 43956 42226
rect 43904 42162 43956 42168
rect 42812 42090 42840 42162
rect 42800 42084 42852 42090
rect 42800 42026 42852 42032
rect 42524 41676 42576 41682
rect 42524 41618 42576 41624
rect 41708 41386 42196 41414
rect 41512 41064 41564 41070
rect 41512 41006 41564 41012
rect 40684 40656 40736 40662
rect 40684 40598 40736 40604
rect 39948 40520 40000 40526
rect 39948 40462 40000 40468
rect 40040 40520 40092 40526
rect 40040 40462 40092 40468
rect 40500 40520 40552 40526
rect 40500 40462 40552 40468
rect 39212 40384 39264 40390
rect 39212 40326 39264 40332
rect 38936 39908 38988 39914
rect 38936 39850 38988 39856
rect 38948 39642 38976 39850
rect 39224 39642 39252 40326
rect 39488 40112 39540 40118
rect 39488 40054 39540 40060
rect 39396 39840 39448 39846
rect 39396 39782 39448 39788
rect 38936 39636 38988 39642
rect 38936 39578 38988 39584
rect 39212 39636 39264 39642
rect 39212 39578 39264 39584
rect 38948 38962 38976 39578
rect 39224 39438 39252 39578
rect 39408 39574 39436 39782
rect 39500 39642 39528 40054
rect 39960 39982 39988 40462
rect 39948 39976 40000 39982
rect 39948 39918 40000 39924
rect 39488 39636 39540 39642
rect 39488 39578 39540 39584
rect 39396 39568 39448 39574
rect 39396 39510 39448 39516
rect 39212 39432 39264 39438
rect 39212 39374 39264 39380
rect 39304 39364 39356 39370
rect 39304 39306 39356 39312
rect 39316 38962 39344 39306
rect 38844 38956 38896 38962
rect 38844 38898 38896 38904
rect 38936 38956 38988 38962
rect 38936 38898 38988 38904
rect 39304 38956 39356 38962
rect 39304 38898 39356 38904
rect 38856 38418 38884 38898
rect 39120 38888 39172 38894
rect 39120 38830 39172 38836
rect 38660 38412 38712 38418
rect 38660 38354 38712 38360
rect 38844 38412 38896 38418
rect 38844 38354 38896 38360
rect 38672 38010 38700 38354
rect 38844 38208 38896 38214
rect 38844 38150 38896 38156
rect 38660 38004 38712 38010
rect 38660 37946 38712 37952
rect 38660 36780 38712 36786
rect 38660 36722 38712 36728
rect 38476 35692 38528 35698
rect 38476 35634 38528 35640
rect 38488 35222 38516 35634
rect 38476 35216 38528 35222
rect 38476 35158 38528 35164
rect 38488 34746 38516 35158
rect 38672 35154 38700 36722
rect 38752 36304 38804 36310
rect 38752 36246 38804 36252
rect 38764 35698 38792 36246
rect 38856 36242 38884 38150
rect 39132 37330 39160 38830
rect 39120 37324 39172 37330
rect 39120 37266 39172 37272
rect 39304 37256 39356 37262
rect 39304 37198 39356 37204
rect 38936 37120 38988 37126
rect 38936 37062 38988 37068
rect 38948 36786 38976 37062
rect 38936 36780 38988 36786
rect 38936 36722 38988 36728
rect 38844 36236 38896 36242
rect 38844 36178 38896 36184
rect 38936 36168 38988 36174
rect 38936 36110 38988 36116
rect 38752 35692 38804 35698
rect 38752 35634 38804 35640
rect 38660 35148 38712 35154
rect 38660 35090 38712 35096
rect 38568 35012 38620 35018
rect 38568 34954 38620 34960
rect 38200 34740 38252 34746
rect 38200 34682 38252 34688
rect 38476 34740 38528 34746
rect 38476 34682 38528 34688
rect 38212 33590 38240 34682
rect 38580 34610 38608 34954
rect 38568 34604 38620 34610
rect 38568 34546 38620 34552
rect 38384 34536 38436 34542
rect 38384 34478 38436 34484
rect 38396 33658 38424 34478
rect 38568 34128 38620 34134
rect 38568 34070 38620 34076
rect 38384 33652 38436 33658
rect 38384 33594 38436 33600
rect 38200 33584 38252 33590
rect 38200 33526 38252 33532
rect 38396 32434 38424 33594
rect 38580 33522 38608 34070
rect 38568 33516 38620 33522
rect 38568 33458 38620 33464
rect 38672 32978 38700 35090
rect 38948 34950 38976 36110
rect 39316 35834 39344 37198
rect 39304 35828 39356 35834
rect 39304 35770 39356 35776
rect 39408 35494 39436 39510
rect 39672 39432 39724 39438
rect 39672 39374 39724 39380
rect 39684 38962 39712 39374
rect 39672 38956 39724 38962
rect 39672 38898 39724 38904
rect 39684 38282 39712 38898
rect 39856 38752 39908 38758
rect 39856 38694 39908 38700
rect 39868 38350 39896 38694
rect 39960 38418 39988 39918
rect 40052 39914 40080 40462
rect 40040 39908 40092 39914
rect 40040 39850 40092 39856
rect 40512 39438 40540 40462
rect 40592 40384 40644 40390
rect 40592 40326 40644 40332
rect 40500 39432 40552 39438
rect 40500 39374 40552 39380
rect 40604 39370 40632 40326
rect 40696 40118 40724 40598
rect 40776 40452 40828 40458
rect 40776 40394 40828 40400
rect 40684 40112 40736 40118
rect 40684 40054 40736 40060
rect 40788 39642 40816 40394
rect 40776 39636 40828 39642
rect 40776 39578 40828 39584
rect 41052 39568 41104 39574
rect 41052 39510 41104 39516
rect 40776 39500 40828 39506
rect 40776 39442 40828 39448
rect 40592 39364 40644 39370
rect 40592 39306 40644 39312
rect 40788 39302 40816 39442
rect 40776 39296 40828 39302
rect 40776 39238 40828 39244
rect 41064 38894 41092 39510
rect 40776 38888 40828 38894
rect 40776 38830 40828 38836
rect 41052 38888 41104 38894
rect 41052 38830 41104 38836
rect 40040 38820 40092 38826
rect 40040 38762 40092 38768
rect 39948 38412 40000 38418
rect 39948 38354 40000 38360
rect 39856 38344 39908 38350
rect 39856 38286 39908 38292
rect 39672 38276 39724 38282
rect 39672 38218 39724 38224
rect 39580 38208 39632 38214
rect 39580 38150 39632 38156
rect 39592 37942 39620 38150
rect 39580 37936 39632 37942
rect 39580 37878 39632 37884
rect 39960 37874 39988 38354
rect 40052 38350 40080 38762
rect 40040 38344 40092 38350
rect 40040 38286 40092 38292
rect 39948 37868 40000 37874
rect 39948 37810 40000 37816
rect 39960 37194 39988 37810
rect 39948 37188 40000 37194
rect 39948 37130 40000 37136
rect 39960 36854 39988 37130
rect 40224 37120 40276 37126
rect 40224 37062 40276 37068
rect 39948 36848 40000 36854
rect 39948 36790 40000 36796
rect 40040 36576 40092 36582
rect 40040 36518 40092 36524
rect 40052 36378 40080 36518
rect 40236 36378 40264 37062
rect 40788 36922 40816 38830
rect 41064 37874 41092 38830
rect 41708 38298 41736 41386
rect 41880 39840 41932 39846
rect 41880 39782 41932 39788
rect 41892 39438 41920 39782
rect 42706 39536 42762 39545
rect 42706 39471 42708 39480
rect 42760 39471 42762 39480
rect 42708 39442 42760 39448
rect 41880 39432 41932 39438
rect 41880 39374 41932 39380
rect 41144 38276 41196 38282
rect 41144 38218 41196 38224
rect 41524 38270 41736 38298
rect 41156 38010 41184 38218
rect 41144 38004 41196 38010
rect 41144 37946 41196 37952
rect 41052 37868 41104 37874
rect 41052 37810 41104 37816
rect 41420 37256 41472 37262
rect 41420 37198 41472 37204
rect 40776 36916 40828 36922
rect 40776 36858 40828 36864
rect 41432 36854 41460 37198
rect 41420 36848 41472 36854
rect 41420 36790 41472 36796
rect 40040 36372 40092 36378
rect 40040 36314 40092 36320
rect 40224 36372 40276 36378
rect 40224 36314 40276 36320
rect 40500 36304 40552 36310
rect 41524 36258 41552 38270
rect 41604 38208 41656 38214
rect 41604 38150 41656 38156
rect 41616 37330 41644 38150
rect 41696 37460 41748 37466
rect 41696 37402 41748 37408
rect 41604 37324 41656 37330
rect 41604 37266 41656 37272
rect 41616 36922 41644 37266
rect 41708 36922 41736 37402
rect 41892 37194 41920 39374
rect 42708 38412 42760 38418
rect 42708 38354 42760 38360
rect 42432 38208 42484 38214
rect 42720 38185 42748 38354
rect 42432 38150 42484 38156
rect 42706 38176 42762 38185
rect 42444 37874 42472 38150
rect 42706 38111 42762 38120
rect 42432 37868 42484 37874
rect 42432 37810 42484 37816
rect 42708 37800 42760 37806
rect 42708 37742 42760 37748
rect 42432 37732 42484 37738
rect 42432 37674 42484 37680
rect 42248 37664 42300 37670
rect 42248 37606 42300 37612
rect 42260 37194 42288 37606
rect 41880 37188 41932 37194
rect 41880 37130 41932 37136
rect 42248 37188 42300 37194
rect 42248 37130 42300 37136
rect 42444 36922 42472 37674
rect 42720 37466 42748 37742
rect 42708 37460 42760 37466
rect 42708 37402 42760 37408
rect 41604 36916 41656 36922
rect 41604 36858 41656 36864
rect 41696 36916 41748 36922
rect 41696 36858 41748 36864
rect 42432 36916 42484 36922
rect 42432 36858 42484 36864
rect 41708 36582 41736 36858
rect 41972 36848 42024 36854
rect 41972 36790 42024 36796
rect 42614 36816 42670 36825
rect 41984 36718 42012 36790
rect 42614 36751 42670 36760
rect 41972 36712 42024 36718
rect 41972 36654 42024 36660
rect 41696 36576 41748 36582
rect 41696 36518 41748 36524
rect 40500 36246 40552 36252
rect 40040 36168 40092 36174
rect 40040 36110 40092 36116
rect 39856 36032 39908 36038
rect 39856 35974 39908 35980
rect 39764 35624 39816 35630
rect 39764 35566 39816 35572
rect 39672 35556 39724 35562
rect 39672 35498 39724 35504
rect 39396 35488 39448 35494
rect 39396 35430 39448 35436
rect 39684 35222 39712 35498
rect 39672 35216 39724 35222
rect 39672 35158 39724 35164
rect 38936 34944 38988 34950
rect 38936 34886 38988 34892
rect 38948 34610 38976 34886
rect 39776 34610 39804 35566
rect 39868 35290 39896 35974
rect 40052 35834 40080 36110
rect 40040 35828 40092 35834
rect 40040 35770 40092 35776
rect 39856 35284 39908 35290
rect 39856 35226 39908 35232
rect 39948 35148 40000 35154
rect 39948 35090 40000 35096
rect 38936 34604 38988 34610
rect 38936 34546 38988 34552
rect 39764 34604 39816 34610
rect 39764 34546 39816 34552
rect 38752 34400 38804 34406
rect 38752 34342 38804 34348
rect 38764 33930 38792 34342
rect 38844 33992 38896 33998
rect 38844 33934 38896 33940
rect 38752 33924 38804 33930
rect 38752 33866 38804 33872
rect 38856 33590 38884 33934
rect 38844 33584 38896 33590
rect 38844 33526 38896 33532
rect 38948 33386 38976 34546
rect 39120 33856 39172 33862
rect 39120 33798 39172 33804
rect 38936 33380 38988 33386
rect 38936 33322 38988 33328
rect 38660 32972 38712 32978
rect 38660 32914 38712 32920
rect 38948 32570 38976 33322
rect 39132 32910 39160 33798
rect 39776 33522 39804 34546
rect 39960 34066 39988 35090
rect 40052 34542 40080 35770
rect 40512 35698 40540 36246
rect 41432 36230 41552 36258
rect 40868 36168 40920 36174
rect 40868 36110 40920 36116
rect 40684 36032 40736 36038
rect 40684 35974 40736 35980
rect 40500 35692 40552 35698
rect 40500 35634 40552 35640
rect 40696 35018 40724 35974
rect 40880 35834 40908 36110
rect 40868 35828 40920 35834
rect 40868 35770 40920 35776
rect 41432 35714 41460 36230
rect 41512 36168 41564 36174
rect 41512 36110 41564 36116
rect 41340 35686 41460 35714
rect 40684 35012 40736 35018
rect 40684 34954 40736 34960
rect 40132 34604 40184 34610
rect 40132 34546 40184 34552
rect 40040 34536 40092 34542
rect 40040 34478 40092 34484
rect 39948 34060 40000 34066
rect 39948 34002 40000 34008
rect 40052 33862 40080 34478
rect 40040 33856 40092 33862
rect 40040 33798 40092 33804
rect 40052 33590 40080 33798
rect 40144 33658 40172 34546
rect 41236 34536 41288 34542
rect 41236 34478 41288 34484
rect 41340 34490 41368 35686
rect 41524 34746 41552 36110
rect 41604 36032 41656 36038
rect 41604 35974 41656 35980
rect 41616 35086 41644 35974
rect 41708 35834 41736 36518
rect 41696 35828 41748 35834
rect 41696 35770 41748 35776
rect 41708 35290 41736 35770
rect 41984 35698 42012 36654
rect 42064 36644 42116 36650
rect 42064 36586 42116 36592
rect 42076 36174 42104 36586
rect 42064 36168 42116 36174
rect 42064 36110 42116 36116
rect 42076 35834 42104 36110
rect 42064 35828 42116 35834
rect 42064 35770 42116 35776
rect 41972 35692 42024 35698
rect 41972 35634 42024 35640
rect 41696 35284 41748 35290
rect 41696 35226 41748 35232
rect 41604 35080 41656 35086
rect 41604 35022 41656 35028
rect 41512 34740 41564 34746
rect 41512 34682 41564 34688
rect 41708 34610 41736 35226
rect 41696 34604 41748 34610
rect 41696 34546 41748 34552
rect 40224 34400 40276 34406
rect 40224 34342 40276 34348
rect 40236 33998 40264 34342
rect 41248 34202 41276 34478
rect 41340 34462 41460 34490
rect 41984 34474 42012 35634
rect 41236 34196 41288 34202
rect 41236 34138 41288 34144
rect 40224 33992 40276 33998
rect 40224 33934 40276 33940
rect 40132 33652 40184 33658
rect 40132 33594 40184 33600
rect 40040 33584 40092 33590
rect 40040 33526 40092 33532
rect 39764 33516 39816 33522
rect 39764 33458 39816 33464
rect 39120 32904 39172 32910
rect 39120 32846 39172 32852
rect 39948 32768 40000 32774
rect 39948 32710 40000 32716
rect 38936 32564 38988 32570
rect 38936 32506 38988 32512
rect 39960 32434 39988 32710
rect 38384 32428 38436 32434
rect 38384 32370 38436 32376
rect 39948 32428 40000 32434
rect 39948 32370 40000 32376
rect 41432 26450 41460 34462
rect 41972 34468 42024 34474
rect 41972 34410 42024 34416
rect 42340 34400 42392 34406
rect 42340 34342 42392 34348
rect 42352 34066 42380 34342
rect 42340 34060 42392 34066
rect 42340 34002 42392 34008
rect 42340 32904 42392 32910
rect 42340 32846 42392 32852
rect 42352 32434 42380 32846
rect 42340 32428 42392 32434
rect 42340 32370 42392 32376
rect 41420 26444 41472 26450
rect 41420 26386 41472 26392
rect 41604 26376 41656 26382
rect 41604 26318 41656 26324
rect 41616 26042 41644 26318
rect 41788 26308 41840 26314
rect 41788 26250 41840 26256
rect 41604 26036 41656 26042
rect 41604 25978 41656 25984
rect 41418 25936 41474 25945
rect 38936 25900 38988 25906
rect 41418 25871 41474 25880
rect 41696 25900 41748 25906
rect 38936 25842 38988 25848
rect 38948 25498 38976 25842
rect 38936 25492 38988 25498
rect 38936 25434 38988 25440
rect 41432 25362 41460 25871
rect 41696 25842 41748 25848
rect 41420 25356 41472 25362
rect 41420 25298 41472 25304
rect 39304 25288 39356 25294
rect 39304 25230 39356 25236
rect 39316 24954 39344 25230
rect 40868 25220 40920 25226
rect 40868 25162 40920 25168
rect 39304 24948 39356 24954
rect 39304 24890 39356 24896
rect 38568 24812 38620 24818
rect 38568 24754 38620 24760
rect 40040 24812 40092 24818
rect 40040 24754 40092 24760
rect 38016 24200 38068 24206
rect 38016 24142 38068 24148
rect 38028 23322 38056 24142
rect 38580 23866 38608 24754
rect 39948 24744 40000 24750
rect 39948 24686 40000 24692
rect 38752 24132 38804 24138
rect 38752 24074 38804 24080
rect 38568 23860 38620 23866
rect 38568 23802 38620 23808
rect 38764 23662 38792 24074
rect 39028 23724 39080 23730
rect 39028 23666 39080 23672
rect 38752 23656 38804 23662
rect 38752 23598 38804 23604
rect 38844 23656 38896 23662
rect 38844 23598 38896 23604
rect 38016 23316 38068 23322
rect 38016 23258 38068 23264
rect 38764 23118 38792 23598
rect 38856 23118 38884 23598
rect 39040 23118 39068 23666
rect 39960 23186 39988 24686
rect 39948 23180 40000 23186
rect 39948 23122 40000 23128
rect 38752 23112 38804 23118
rect 38752 23054 38804 23060
rect 38844 23112 38896 23118
rect 38844 23054 38896 23060
rect 39028 23112 39080 23118
rect 39028 23054 39080 23060
rect 38200 22976 38252 22982
rect 38200 22918 38252 22924
rect 38212 22642 38240 22918
rect 38200 22636 38252 22642
rect 38200 22578 38252 22584
rect 38764 22506 38792 23054
rect 39040 22710 39068 23054
rect 40052 22778 40080 24754
rect 40880 24206 40908 25162
rect 41512 24608 41564 24614
rect 41512 24550 41564 24556
rect 41524 24274 41552 24550
rect 41708 24410 41736 25842
rect 41800 24750 41828 26250
rect 42340 25288 42392 25294
rect 42340 25230 42392 25236
rect 41788 24744 41840 24750
rect 41788 24686 41840 24692
rect 41696 24404 41748 24410
rect 41696 24346 41748 24352
rect 41512 24268 41564 24274
rect 41512 24210 41564 24216
rect 40868 24200 40920 24206
rect 40868 24142 40920 24148
rect 41604 24200 41656 24206
rect 41604 24142 41656 24148
rect 41696 24200 41748 24206
rect 41696 24142 41748 24148
rect 41616 23730 41644 24142
rect 41604 23724 41656 23730
rect 41604 23666 41656 23672
rect 40040 22772 40092 22778
rect 40040 22714 40092 22720
rect 38844 22704 38896 22710
rect 38844 22646 38896 22652
rect 39028 22704 39080 22710
rect 39028 22646 39080 22652
rect 38856 22574 38884 22646
rect 41616 22642 41644 23666
rect 39120 22636 39172 22642
rect 39120 22578 39172 22584
rect 41604 22636 41656 22642
rect 41604 22578 41656 22584
rect 38844 22568 38896 22574
rect 38844 22510 38896 22516
rect 38752 22500 38804 22506
rect 38752 22442 38804 22448
rect 38108 22432 38160 22438
rect 38108 22374 38160 22380
rect 37924 20596 37976 20602
rect 37924 20538 37976 20544
rect 38120 20466 38148 22374
rect 38764 22166 38792 22442
rect 38752 22160 38804 22166
rect 38752 22102 38804 22108
rect 38764 21962 38792 22102
rect 38856 22030 38884 22510
rect 39132 22030 39160 22578
rect 38844 22024 38896 22030
rect 38844 21966 38896 21972
rect 39120 22024 39172 22030
rect 39120 21966 39172 21972
rect 40408 22024 40460 22030
rect 40408 21966 40460 21972
rect 41420 22024 41472 22030
rect 41420 21966 41472 21972
rect 38752 21956 38804 21962
rect 38752 21898 38804 21904
rect 38200 21888 38252 21894
rect 38200 21830 38252 21836
rect 38212 21554 38240 21830
rect 38200 21548 38252 21554
rect 38200 21490 38252 21496
rect 38752 21480 38804 21486
rect 38752 21422 38804 21428
rect 38764 20942 38792 21422
rect 38856 21146 38884 21966
rect 39132 21690 39160 21966
rect 40132 21956 40184 21962
rect 40132 21898 40184 21904
rect 39764 21888 39816 21894
rect 39764 21830 39816 21836
rect 39120 21684 39172 21690
rect 39120 21626 39172 21632
rect 38844 21140 38896 21146
rect 38844 21082 38896 21088
rect 38752 20936 38804 20942
rect 38752 20878 38804 20884
rect 39776 20466 39804 21830
rect 40144 21690 40172 21898
rect 40132 21684 40184 21690
rect 40132 21626 40184 21632
rect 40132 20868 40184 20874
rect 40132 20810 40184 20816
rect 38108 20460 38160 20466
rect 38108 20402 38160 20408
rect 39764 20460 39816 20466
rect 39764 20402 39816 20408
rect 39304 20256 39356 20262
rect 39304 20198 39356 20204
rect 39316 19922 39344 20198
rect 39304 19916 39356 19922
rect 39304 19858 39356 19864
rect 40144 19854 40172 20810
rect 40420 20534 40448 21966
rect 41432 21865 41460 21966
rect 41418 21856 41474 21865
rect 41418 21791 41474 21800
rect 41052 21004 41104 21010
rect 41052 20946 41104 20952
rect 41064 20602 41092 20946
rect 41328 20800 41380 20806
rect 41328 20742 41380 20748
rect 41052 20596 41104 20602
rect 41052 20538 41104 20544
rect 40408 20528 40460 20534
rect 40408 20470 40460 20476
rect 40132 19848 40184 19854
rect 40132 19790 40184 19796
rect 36912 19712 36964 19718
rect 36912 19654 36964 19660
rect 38936 19712 38988 19718
rect 38936 19654 38988 19660
rect 36924 18766 36952 19654
rect 38948 19378 38976 19654
rect 38936 19372 38988 19378
rect 38936 19314 38988 19320
rect 38752 19168 38804 19174
rect 38752 19110 38804 19116
rect 36912 18760 36964 18766
rect 36912 18702 36964 18708
rect 35716 18624 35768 18630
rect 35716 18566 35768 18572
rect 37464 18624 37516 18630
rect 37464 18566 37516 18572
rect 38384 18624 38436 18630
rect 38384 18566 38436 18572
rect 35728 18358 35756 18566
rect 35716 18352 35768 18358
rect 35716 18294 35768 18300
rect 35728 17882 35756 18294
rect 37476 18290 37504 18566
rect 38396 18358 38424 18566
rect 38384 18352 38436 18358
rect 38384 18294 38436 18300
rect 35808 18284 35860 18290
rect 35808 18226 35860 18232
rect 35992 18284 36044 18290
rect 35992 18226 36044 18232
rect 37464 18284 37516 18290
rect 37464 18226 37516 18232
rect 35716 17876 35768 17882
rect 35716 17818 35768 17824
rect 35820 17678 35848 18226
rect 36004 17882 36032 18226
rect 38764 18222 38792 19110
rect 38752 18216 38804 18222
rect 38752 18158 38804 18164
rect 39948 18216 40000 18222
rect 39948 18158 40000 18164
rect 37280 18080 37332 18086
rect 37280 18022 37332 18028
rect 37464 18080 37516 18086
rect 37464 18022 37516 18028
rect 35992 17876 36044 17882
rect 35992 17818 36044 17824
rect 35808 17672 35860 17678
rect 35808 17614 35860 17620
rect 37004 17672 37056 17678
rect 37004 17614 37056 17620
rect 35716 17536 35768 17542
rect 35716 17478 35768 17484
rect 35728 17270 35756 17478
rect 35716 17264 35768 17270
rect 35716 17206 35768 17212
rect 35820 17082 35848 17614
rect 37016 17202 37044 17614
rect 37004 17196 37056 17202
rect 37004 17138 37056 17144
rect 35820 17066 35940 17082
rect 35820 17060 35952 17066
rect 35820 17054 35900 17060
rect 35900 17002 35952 17008
rect 37016 16590 37044 17138
rect 37004 16584 37056 16590
rect 37004 16526 37056 16532
rect 37292 16538 37320 18022
rect 37476 17202 37504 18022
rect 38108 17740 38160 17746
rect 38108 17682 38160 17688
rect 37464 17196 37516 17202
rect 37464 17138 37516 17144
rect 37476 16658 37504 17138
rect 37464 16652 37516 16658
rect 37464 16594 37516 16600
rect 37924 16584 37976 16590
rect 35808 16516 35860 16522
rect 37292 16510 37412 16538
rect 37924 16526 37976 16532
rect 35808 16458 35860 16464
rect 35820 16114 35848 16458
rect 37280 16448 37332 16454
rect 37280 16390 37332 16396
rect 35808 16108 35860 16114
rect 35808 16050 35860 16056
rect 35820 15502 35848 16050
rect 36268 16040 36320 16046
rect 36268 15982 36320 15988
rect 36084 15632 36136 15638
rect 36084 15574 36136 15580
rect 35808 15496 35860 15502
rect 35808 15438 35860 15444
rect 35820 13938 35848 15438
rect 36096 15094 36124 15574
rect 36084 15088 36136 15094
rect 36084 15030 36136 15036
rect 36280 15026 36308 15982
rect 37292 15434 37320 16390
rect 37384 16182 37412 16510
rect 37372 16176 37424 16182
rect 37372 16118 37424 16124
rect 37384 15570 37412 16118
rect 37936 15910 37964 16526
rect 38120 16114 38148 17682
rect 38936 16992 38988 16998
rect 38936 16934 38988 16940
rect 38108 16108 38160 16114
rect 38108 16050 38160 16056
rect 37464 15904 37516 15910
rect 37464 15846 37516 15852
rect 37924 15904 37976 15910
rect 37924 15846 37976 15852
rect 37372 15564 37424 15570
rect 37372 15506 37424 15512
rect 37280 15428 37332 15434
rect 37280 15370 37332 15376
rect 36820 15360 36872 15366
rect 36820 15302 36872 15308
rect 36832 15026 36860 15302
rect 37292 15094 37320 15370
rect 37384 15366 37412 15506
rect 37372 15360 37424 15366
rect 37372 15302 37424 15308
rect 37280 15088 37332 15094
rect 37280 15030 37332 15036
rect 35992 15020 36044 15026
rect 35992 14962 36044 14968
rect 36268 15020 36320 15026
rect 36268 14962 36320 14968
rect 36452 15020 36504 15026
rect 36452 14962 36504 14968
rect 36820 15020 36872 15026
rect 36820 14962 36872 14968
rect 36004 14618 36032 14962
rect 35992 14612 36044 14618
rect 35992 14554 36044 14560
rect 36464 14550 36492 14962
rect 36544 14884 36596 14890
rect 36544 14826 36596 14832
rect 36556 14618 36584 14826
rect 36544 14612 36596 14618
rect 36544 14554 36596 14560
rect 36452 14544 36504 14550
rect 36452 14486 36504 14492
rect 35808 13932 35860 13938
rect 35808 13874 35860 13880
rect 36464 13870 36492 14486
rect 36832 14482 36860 14962
rect 37384 14958 37412 15302
rect 37476 15026 37504 15846
rect 37740 15496 37792 15502
rect 37740 15438 37792 15444
rect 37464 15020 37516 15026
rect 37464 14962 37516 14968
rect 37372 14952 37424 14958
rect 37372 14894 37424 14900
rect 37464 14884 37516 14890
rect 37464 14826 37516 14832
rect 37648 14884 37700 14890
rect 37648 14826 37700 14832
rect 37280 14816 37332 14822
rect 37280 14758 37332 14764
rect 36820 14476 36872 14482
rect 36820 14418 36872 14424
rect 37292 14414 37320 14758
rect 37476 14634 37504 14826
rect 37476 14606 37596 14634
rect 37464 14476 37516 14482
rect 37464 14418 37516 14424
rect 37280 14408 37332 14414
rect 37280 14350 37332 14356
rect 36544 14272 36596 14278
rect 36544 14214 36596 14220
rect 36556 14074 36584 14214
rect 36544 14068 36596 14074
rect 36544 14010 36596 14016
rect 37096 14000 37148 14006
rect 37096 13942 37148 13948
rect 37108 13870 37136 13942
rect 37372 13932 37424 13938
rect 37372 13874 37424 13880
rect 36452 13864 36504 13870
rect 36452 13806 36504 13812
rect 37096 13864 37148 13870
rect 37096 13806 37148 13812
rect 36084 13184 36136 13190
rect 36084 13126 36136 13132
rect 36096 12986 36124 13126
rect 36084 12980 36136 12986
rect 36084 12922 36136 12928
rect 36544 12844 36596 12850
rect 36544 12786 36596 12792
rect 35716 12776 35768 12782
rect 35716 12718 35768 12724
rect 35728 11898 35756 12718
rect 35900 12096 35952 12102
rect 35900 12038 35952 12044
rect 36268 12096 36320 12102
rect 36268 12038 36320 12044
rect 35716 11892 35768 11898
rect 35716 11834 35768 11840
rect 35728 11626 35756 11834
rect 35912 11830 35940 12038
rect 35900 11824 35952 11830
rect 35900 11766 35952 11772
rect 36176 11688 36228 11694
rect 36176 11630 36228 11636
rect 35716 11620 35768 11626
rect 35716 11562 35768 11568
rect 36188 11218 36216 11630
rect 36280 11626 36308 12038
rect 36556 11898 36584 12786
rect 36544 11892 36596 11898
rect 36544 11834 36596 11840
rect 37108 11830 37136 13806
rect 37280 13728 37332 13734
rect 37280 13670 37332 13676
rect 36636 11824 36688 11830
rect 36636 11766 36688 11772
rect 37096 11824 37148 11830
rect 37292 11778 37320 13670
rect 37384 13326 37412 13874
rect 37476 13734 37504 14418
rect 37568 13870 37596 14606
rect 37556 13864 37608 13870
rect 37556 13806 37608 13812
rect 37464 13728 37516 13734
rect 37464 13670 37516 13676
rect 37372 13320 37424 13326
rect 37372 13262 37424 13268
rect 37568 11830 37596 13806
rect 37660 13326 37688 14826
rect 37752 14482 37780 15438
rect 37936 14958 37964 15846
rect 37924 14952 37976 14958
rect 37924 14894 37976 14900
rect 37740 14476 37792 14482
rect 37740 14418 37792 14424
rect 37752 14006 37780 14418
rect 38016 14408 38068 14414
rect 38016 14350 38068 14356
rect 38028 14249 38056 14350
rect 38014 14240 38070 14249
rect 38014 14175 38070 14184
rect 37740 14000 37792 14006
rect 37740 13942 37792 13948
rect 38016 13388 38068 13394
rect 38016 13330 38068 13336
rect 37648 13320 37700 13326
rect 37648 13262 37700 13268
rect 37832 13320 37884 13326
rect 37832 13262 37884 13268
rect 37660 12238 37688 13262
rect 37844 12986 37872 13262
rect 37832 12980 37884 12986
rect 37832 12922 37884 12928
rect 37648 12232 37700 12238
rect 37648 12174 37700 12180
rect 37096 11766 37148 11772
rect 36268 11620 36320 11626
rect 36268 11562 36320 11568
rect 36176 11212 36228 11218
rect 36176 11154 36228 11160
rect 36648 11082 36676 11766
rect 37200 11762 37320 11778
rect 37556 11824 37608 11830
rect 37556 11766 37608 11772
rect 37188 11756 37320 11762
rect 37240 11750 37320 11756
rect 37188 11698 37240 11704
rect 37372 11688 37424 11694
rect 37372 11630 37424 11636
rect 37384 11150 37412 11630
rect 37372 11144 37424 11150
rect 37372 11086 37424 11092
rect 37660 11082 37688 12174
rect 37844 11558 37872 12922
rect 38028 12850 38056 13330
rect 38120 13274 38148 16050
rect 38948 15502 38976 16934
rect 38936 15496 38988 15502
rect 38988 15444 39160 15450
rect 38936 15438 39160 15444
rect 38948 15422 39160 15438
rect 39028 15360 39080 15366
rect 39028 15302 39080 15308
rect 38936 15020 38988 15026
rect 38936 14962 38988 14968
rect 38384 14952 38436 14958
rect 38384 14894 38436 14900
rect 38292 14816 38344 14822
rect 38292 14758 38344 14764
rect 38200 14544 38252 14550
rect 38200 14486 38252 14492
rect 38212 14074 38240 14486
rect 38200 14068 38252 14074
rect 38200 14010 38252 14016
rect 38304 13734 38332 14758
rect 38396 14074 38424 14894
rect 38948 14822 38976 14962
rect 38936 14816 38988 14822
rect 38936 14758 38988 14764
rect 39040 14482 39068 15302
rect 39028 14476 39080 14482
rect 39028 14418 39080 14424
rect 38568 14408 38620 14414
rect 38488 14368 38568 14396
rect 38384 14068 38436 14074
rect 38384 14010 38436 14016
rect 38488 14006 38516 14368
rect 38568 14350 38620 14356
rect 38936 14340 38988 14346
rect 38936 14282 38988 14288
rect 38568 14272 38620 14278
rect 38566 14240 38568 14249
rect 38620 14240 38622 14249
rect 38566 14175 38622 14184
rect 38568 14068 38620 14074
rect 38568 14010 38620 14016
rect 38476 14000 38528 14006
rect 38476 13942 38528 13948
rect 38292 13728 38344 13734
rect 38292 13670 38344 13676
rect 38304 13546 38332 13670
rect 38304 13530 38424 13546
rect 38292 13524 38424 13530
rect 38344 13518 38424 13524
rect 38292 13466 38344 13472
rect 38120 13258 38240 13274
rect 38120 13252 38252 13258
rect 38120 13246 38200 13252
rect 38200 13194 38252 13200
rect 38108 13184 38160 13190
rect 38108 13126 38160 13132
rect 38016 12844 38068 12850
rect 38016 12786 38068 12792
rect 38120 11830 38148 13126
rect 38200 12844 38252 12850
rect 38200 12786 38252 12792
rect 38108 11824 38160 11830
rect 38108 11766 38160 11772
rect 38212 11762 38240 12786
rect 38396 12434 38424 13518
rect 38580 13410 38608 14010
rect 38844 14000 38896 14006
rect 38844 13942 38896 13948
rect 38580 13382 38700 13410
rect 38672 13258 38700 13382
rect 38568 13252 38620 13258
rect 38568 13194 38620 13200
rect 38660 13252 38712 13258
rect 38660 13194 38712 13200
rect 38580 12782 38608 13194
rect 38672 12918 38700 13194
rect 38660 12912 38712 12918
rect 38660 12854 38712 12860
rect 38568 12776 38620 12782
rect 38568 12718 38620 12724
rect 38304 12406 38424 12434
rect 38304 12306 38332 12406
rect 38292 12300 38344 12306
rect 38292 12242 38344 12248
rect 38856 12170 38884 13942
rect 38948 13530 38976 14282
rect 39132 13802 39160 15422
rect 39120 13796 39172 13802
rect 39120 13738 39172 13744
rect 38936 13524 38988 13530
rect 38936 13466 38988 13472
rect 38948 12374 38976 13466
rect 39132 13326 39160 13738
rect 39120 13320 39172 13326
rect 39120 13262 39172 13268
rect 38936 12368 38988 12374
rect 38936 12310 38988 12316
rect 38844 12164 38896 12170
rect 38844 12106 38896 12112
rect 38292 12096 38344 12102
rect 38292 12038 38344 12044
rect 38304 11762 38332 12038
rect 38200 11756 38252 11762
rect 38200 11698 38252 11704
rect 38292 11756 38344 11762
rect 38292 11698 38344 11704
rect 37832 11552 37884 11558
rect 37832 11494 37884 11500
rect 36636 11076 36688 11082
rect 36636 11018 36688 11024
rect 37648 11076 37700 11082
rect 37648 11018 37700 11024
rect 35544 6886 35664 6914
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 18696 4140 18748 4146
rect 18696 4082 18748 4088
rect 16120 3596 16172 3602
rect 16120 3538 16172 3544
rect 15936 2644 15988 2650
rect 15936 2586 15988 2592
rect 12440 2576 12492 2582
rect 12440 2518 12492 2524
rect 11888 2508 11940 2514
rect 11888 2450 11940 2456
rect 12256 2508 12308 2514
rect 12256 2450 12308 2456
rect 12268 800 12296 2450
rect 16132 800 16160 3538
rect 16856 3528 16908 3534
rect 16856 3470 16908 3476
rect 16868 2514 16896 3470
rect 18708 3126 18736 4082
rect 20812 3936 20864 3942
rect 20812 3878 20864 3884
rect 24216 3936 24268 3942
rect 24216 3878 24268 3884
rect 20824 3602 20852 3878
rect 20812 3596 20864 3602
rect 20812 3538 20864 3544
rect 21272 3596 21324 3602
rect 21272 3538 21324 3544
rect 18788 3528 18840 3534
rect 18788 3470 18840 3476
rect 18696 3120 18748 3126
rect 18696 3062 18748 3068
rect 18800 3058 18828 3470
rect 18972 3392 19024 3398
rect 18972 3334 19024 3340
rect 18984 3126 19012 3334
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 18972 3120 19024 3126
rect 18972 3062 19024 3068
rect 18788 3052 18840 3058
rect 18788 2994 18840 3000
rect 19340 2984 19392 2990
rect 19340 2926 19392 2932
rect 17040 2848 17092 2854
rect 17040 2790 17092 2796
rect 17052 2514 17080 2790
rect 16856 2508 16908 2514
rect 16856 2450 16908 2456
rect 17040 2508 17092 2514
rect 17040 2450 17092 2456
rect 17408 2508 17460 2514
rect 17408 2450 17460 2456
rect 17420 800 17448 2450
rect 19352 800 19380 2926
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 21284 800 21312 3538
rect 22100 3528 22152 3534
rect 22100 3470 22152 3476
rect 22112 3058 22140 3470
rect 23756 3392 23808 3398
rect 23756 3334 23808 3340
rect 22100 3052 22152 3058
rect 22100 2994 22152 3000
rect 22284 2984 22336 2990
rect 22284 2926 22336 2932
rect 23204 2984 23256 2990
rect 23204 2926 23256 2932
rect 22296 2650 22324 2926
rect 23020 2916 23072 2922
rect 23020 2858 23072 2864
rect 22284 2644 22336 2650
rect 22284 2586 22336 2592
rect 23032 2582 23060 2858
rect 23020 2576 23072 2582
rect 23020 2518 23072 2524
rect 23216 800 23244 2926
rect 23768 2378 23796 3334
rect 24228 2514 24256 3878
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 24766 3632 24822 3641
rect 35544 3602 35572 6886
rect 38016 4684 38068 4690
rect 38016 4626 38068 4632
rect 37372 4616 37424 4622
rect 37372 4558 37424 4564
rect 37384 4146 37412 4558
rect 37556 4548 37608 4554
rect 37556 4490 37608 4496
rect 36544 4140 36596 4146
rect 36544 4082 36596 4088
rect 37372 4140 37424 4146
rect 37372 4082 37424 4088
rect 36452 4004 36504 4010
rect 36452 3946 36504 3952
rect 36464 3602 36492 3946
rect 36556 3670 36584 4082
rect 37464 4004 37516 4010
rect 37464 3946 37516 3952
rect 37280 3936 37332 3942
rect 37280 3878 37332 3884
rect 36544 3664 36596 3670
rect 36544 3606 36596 3612
rect 24766 3567 24822 3576
rect 35532 3596 35584 3602
rect 24780 3534 24808 3567
rect 35532 3538 35584 3544
rect 36084 3596 36136 3602
rect 36084 3538 36136 3544
rect 36452 3596 36504 3602
rect 36452 3538 36504 3544
rect 24768 3528 24820 3534
rect 24768 3470 24820 3476
rect 29184 3528 29236 3534
rect 29184 3470 29236 3476
rect 35624 3528 35676 3534
rect 35624 3470 35676 3476
rect 24400 3460 24452 3466
rect 24400 3402 24452 3408
rect 24412 3058 24440 3402
rect 24584 3392 24636 3398
rect 24584 3334 24636 3340
rect 24596 3126 24624 3334
rect 24584 3120 24636 3126
rect 24584 3062 24636 3068
rect 29196 3058 29224 3470
rect 29368 3392 29420 3398
rect 29368 3334 29420 3340
rect 29380 3126 29408 3334
rect 29368 3120 29420 3126
rect 29368 3062 29420 3068
rect 35636 3058 35664 3470
rect 24400 3052 24452 3058
rect 24400 2994 24452 3000
rect 29184 3052 29236 3058
rect 29184 2994 29236 3000
rect 35624 3052 35676 3058
rect 35624 2994 35676 3000
rect 25136 2984 25188 2990
rect 25136 2926 25188 2932
rect 29644 2984 29696 2990
rect 29644 2926 29696 2932
rect 24216 2508 24268 2514
rect 24216 2450 24268 2456
rect 24584 2508 24636 2514
rect 24584 2450 24636 2456
rect 23756 2372 23808 2378
rect 23756 2314 23808 2320
rect 24596 1306 24624 2450
rect 24504 1278 24624 1306
rect 24504 800 24532 1278
rect 25148 800 25176 2926
rect 29656 800 29684 2926
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 36096 800 36124 3538
rect 36544 3392 36596 3398
rect 36544 3334 36596 3340
rect 36556 3058 36584 3334
rect 36544 3052 36596 3058
rect 36544 2994 36596 3000
rect 37292 2514 37320 3878
rect 37372 3460 37424 3466
rect 37372 3402 37424 3408
rect 37280 2508 37332 2514
rect 37280 2450 37332 2456
rect 37384 800 37412 3402
rect 37476 2514 37504 3946
rect 37568 3194 37596 4490
rect 37556 3188 37608 3194
rect 37556 3130 37608 3136
rect 37464 2508 37516 2514
rect 37464 2450 37516 2456
rect 38028 800 38056 4626
rect 38200 4072 38252 4078
rect 38200 4014 38252 4020
rect 38844 4072 38896 4078
rect 38844 4014 38896 4020
rect 38212 3534 38240 4014
rect 38292 4004 38344 4010
rect 38292 3946 38344 3952
rect 38304 3738 38332 3946
rect 38856 3738 38884 4014
rect 38292 3732 38344 3738
rect 38292 3674 38344 3680
rect 38844 3732 38896 3738
rect 38844 3674 38896 3680
rect 38200 3528 38252 3534
rect 38200 3470 38252 3476
rect 39960 3466 39988 18158
rect 40144 16522 40172 19790
rect 41340 19378 41368 20742
rect 41420 20052 41472 20058
rect 41420 19994 41472 20000
rect 41432 19378 41460 19994
rect 41616 19922 41644 22578
rect 41708 22234 41736 24142
rect 42352 23866 42380 25230
rect 42524 25220 42576 25226
rect 42524 25162 42576 25168
rect 42432 24812 42484 24818
rect 42432 24754 42484 24760
rect 42444 24206 42472 24754
rect 42536 24410 42564 25162
rect 42524 24404 42576 24410
rect 42524 24346 42576 24352
rect 42432 24200 42484 24206
rect 42432 24142 42484 24148
rect 42340 23860 42392 23866
rect 42340 23802 42392 23808
rect 41788 23724 41840 23730
rect 41788 23666 41840 23672
rect 41800 23322 41828 23666
rect 42340 23520 42392 23526
rect 42340 23462 42392 23468
rect 42524 23520 42576 23526
rect 42524 23462 42576 23468
rect 41788 23316 41840 23322
rect 41788 23258 41840 23264
rect 41696 22228 41748 22234
rect 41696 22170 41748 22176
rect 41708 21554 41736 22170
rect 42352 22098 42380 23462
rect 42432 22568 42484 22574
rect 42432 22510 42484 22516
rect 42444 22234 42472 22510
rect 42432 22228 42484 22234
rect 42432 22170 42484 22176
rect 42536 22098 42564 23462
rect 42628 22098 42656 36751
rect 42708 36236 42760 36242
rect 42708 36178 42760 36184
rect 42720 36145 42748 36178
rect 42706 36136 42762 36145
rect 42706 36071 42762 36080
rect 42706 35456 42762 35465
rect 42706 35391 42762 35400
rect 42720 35154 42748 35391
rect 42708 35148 42760 35154
rect 42708 35090 42760 35096
rect 42706 30016 42762 30025
rect 42706 29951 42762 29960
rect 42720 29714 42748 29951
rect 42708 29708 42760 29714
rect 42708 29650 42760 29656
rect 42708 27532 42760 27538
rect 42708 27474 42760 27480
rect 42720 27305 42748 27474
rect 42706 27296 42762 27305
rect 42706 27231 42762 27240
rect 42706 25256 42762 25265
rect 42706 25191 42762 25200
rect 42720 24274 42748 25191
rect 42708 24268 42760 24274
rect 42708 24210 42760 24216
rect 42812 23866 42840 42026
rect 43352 42016 43404 42022
rect 43352 41958 43404 41964
rect 42892 41744 42944 41750
rect 42892 41686 42944 41692
rect 42904 41414 42932 41686
rect 43260 41472 43312 41478
rect 43260 41414 43312 41420
rect 42904 41386 43024 41414
rect 42892 37800 42944 37806
rect 42892 37742 42944 37748
rect 42904 36718 42932 37742
rect 42892 36712 42944 36718
rect 42892 36654 42944 36660
rect 42892 33312 42944 33318
rect 42892 33254 42944 33260
rect 42904 32978 42932 33254
rect 42892 32972 42944 32978
rect 42892 32914 42944 32920
rect 42996 26234 43024 41386
rect 43272 40594 43300 41414
rect 43364 40594 43392 41958
rect 43444 41064 43496 41070
rect 43444 41006 43496 41012
rect 43260 40588 43312 40594
rect 43260 40530 43312 40536
rect 43352 40588 43404 40594
rect 43352 40530 43404 40536
rect 43456 40474 43484 41006
rect 43364 40446 43484 40474
rect 43168 38956 43220 38962
rect 43168 38898 43220 38904
rect 43076 33516 43128 33522
rect 43076 33458 43128 33464
rect 42904 26206 43024 26234
rect 42800 23860 42852 23866
rect 42800 23802 42852 23808
rect 42800 23724 42852 23730
rect 42800 23666 42852 23672
rect 42706 23216 42762 23225
rect 42706 23151 42708 23160
rect 42760 23151 42762 23160
rect 42708 23122 42760 23128
rect 42812 22778 42840 23666
rect 42800 22772 42852 22778
rect 42800 22714 42852 22720
rect 42340 22092 42392 22098
rect 42340 22034 42392 22040
rect 42524 22092 42576 22098
rect 42524 22034 42576 22040
rect 42616 22092 42668 22098
rect 42616 22034 42668 22040
rect 41696 21548 41748 21554
rect 41696 21490 41748 21496
rect 42064 21344 42116 21350
rect 42064 21286 42116 21292
rect 42616 21344 42668 21350
rect 42616 21286 42668 21292
rect 42076 19922 42104 21286
rect 42628 21010 42656 21286
rect 42616 21004 42668 21010
rect 42616 20946 42668 20952
rect 41604 19916 41656 19922
rect 41604 19858 41656 19864
rect 42064 19916 42116 19922
rect 42064 19858 42116 19864
rect 41512 19848 41564 19854
rect 41512 19790 41564 19796
rect 42614 19816 42670 19825
rect 41524 19514 41552 19790
rect 42614 19751 42670 19760
rect 41512 19508 41564 19514
rect 41512 19450 41564 19456
rect 41328 19372 41380 19378
rect 41328 19314 41380 19320
rect 41420 19372 41472 19378
rect 41420 19314 41472 19320
rect 42628 17814 42656 19751
rect 42706 19136 42762 19145
rect 42706 19071 42762 19080
rect 42720 18834 42748 19071
rect 42708 18828 42760 18834
rect 42708 18770 42760 18776
rect 42616 17808 42668 17814
rect 42616 17750 42668 17756
rect 42338 17096 42394 17105
rect 42338 17031 42394 17040
rect 42352 16590 42380 17031
rect 42340 16584 42392 16590
rect 42340 16526 42392 16532
rect 40132 16516 40184 16522
rect 40132 16458 40184 16464
rect 42708 15904 42760 15910
rect 42708 15846 42760 15852
rect 42614 15736 42670 15745
rect 42614 15671 42670 15680
rect 42628 15570 42656 15671
rect 42616 15564 42668 15570
rect 42616 15506 42668 15512
rect 42720 14482 42748 15846
rect 42708 14476 42760 14482
rect 42708 14418 42760 14424
rect 42800 13728 42852 13734
rect 42800 13670 42852 13676
rect 42812 13394 42840 13670
rect 42800 13388 42852 13394
rect 42800 13330 42852 13336
rect 41418 13016 41474 13025
rect 41418 12951 41474 12960
rect 41432 12782 41460 12951
rect 41420 12776 41472 12782
rect 41420 12718 41472 12724
rect 42708 12300 42760 12306
rect 42708 12242 42760 12248
rect 42720 11665 42748 12242
rect 42904 11762 42932 26206
rect 43088 22642 43116 33458
rect 43076 22636 43128 22642
rect 43076 22578 43128 22584
rect 43076 20868 43128 20874
rect 43076 20810 43128 20816
rect 43088 20602 43116 20810
rect 43076 20596 43128 20602
rect 43076 20538 43128 20544
rect 43076 19916 43128 19922
rect 43076 19858 43128 19864
rect 42984 19372 43036 19378
rect 42984 19314 43036 19320
rect 42996 17746 43024 19314
rect 42984 17740 43036 17746
rect 42984 17682 43036 17688
rect 42984 17604 43036 17610
rect 42984 17546 43036 17552
rect 42996 17202 43024 17546
rect 42984 17196 43036 17202
rect 42984 17138 43036 17144
rect 42892 11756 42944 11762
rect 42892 11698 42944 11704
rect 42706 11656 42762 11665
rect 42706 11591 42762 11600
rect 42524 9376 42576 9382
rect 42524 9318 42576 9324
rect 42536 9042 42564 9318
rect 42524 9036 42576 9042
rect 42524 8978 42576 8984
rect 42340 8968 42392 8974
rect 42340 8910 42392 8916
rect 42352 8498 42380 8910
rect 42340 8492 42392 8498
rect 42340 8434 42392 8440
rect 42708 6860 42760 6866
rect 42708 6802 42760 6808
rect 42720 6225 42748 6802
rect 42706 6216 42762 6225
rect 42706 6151 42762 6160
rect 42708 5772 42760 5778
rect 42708 5714 42760 5720
rect 42524 5024 42576 5030
rect 42524 4966 42576 4972
rect 42536 4690 42564 4966
rect 42524 4684 42576 4690
rect 42524 4626 42576 4632
rect 41328 4072 41380 4078
rect 41328 4014 41380 4020
rect 40040 3528 40092 3534
rect 40040 3470 40092 3476
rect 39948 3460 40000 3466
rect 39948 3402 40000 3408
rect 40052 3058 40080 3470
rect 40224 3392 40276 3398
rect 40224 3334 40276 3340
rect 40040 3052 40092 3058
rect 40040 2994 40092 3000
rect 40236 2990 40264 3334
rect 40224 2984 40276 2990
rect 40224 2926 40276 2932
rect 41236 2984 41288 2990
rect 41236 2926 41288 2932
rect 38660 2508 38712 2514
rect 38660 2450 38712 2456
rect 38672 800 38700 2450
rect 41248 800 41276 2926
rect 41340 2666 41368 4014
rect 41880 3936 41932 3942
rect 41880 3878 41932 3884
rect 42432 3936 42484 3942
rect 42432 3878 42484 3884
rect 41892 3602 41920 3878
rect 42444 3670 42472 3878
rect 42432 3664 42484 3670
rect 42432 3606 42484 3612
rect 41880 3596 41932 3602
rect 41880 3538 41932 3544
rect 42524 3596 42576 3602
rect 42524 3538 42576 3544
rect 41340 2638 41460 2666
rect 41328 2508 41380 2514
rect 41328 2450 41380 2456
rect 41340 1170 41368 2450
rect 41432 2145 41460 2638
rect 41418 2136 41474 2145
rect 41418 2071 41474 2080
rect 41340 1142 41460 1170
rect -10 0 102 800
rect 634 0 746 800
rect 1278 0 1390 800
rect 1922 0 2034 800
rect 3210 0 3322 800
rect 3854 0 3966 800
rect 4498 0 4610 800
rect 5786 0 5898 800
rect 6430 0 6542 800
rect 7074 0 7186 800
rect 8362 0 8474 800
rect 9006 0 9118 800
rect 9650 0 9762 800
rect 10938 0 11050 800
rect 11582 0 11694 800
rect 12226 0 12338 800
rect 13514 0 13626 800
rect 14158 0 14270 800
rect 14802 0 14914 800
rect 16090 0 16202 800
rect 16734 0 16846 800
rect 17378 0 17490 800
rect 18666 0 18778 800
rect 19310 0 19422 800
rect 19954 0 20066 800
rect 21242 0 21354 800
rect 21886 0 21998 800
rect 22530 0 22642 800
rect 23174 0 23286 800
rect 24462 0 24574 800
rect 25106 0 25218 800
rect 25750 0 25862 800
rect 27038 0 27150 800
rect 27682 0 27794 800
rect 28326 0 28438 800
rect 29614 0 29726 800
rect 30258 0 30370 800
rect 30902 0 31014 800
rect 32190 0 32302 800
rect 32834 0 32946 800
rect 33478 0 33590 800
rect 34766 0 34878 800
rect 35410 0 35522 800
rect 36054 0 36166 800
rect 37342 0 37454 800
rect 37986 0 38098 800
rect 38630 0 38742 800
rect 39918 0 40030 800
rect 40562 0 40674 800
rect 41206 0 41318 800
rect 41432 82 41460 1142
rect 42536 800 42564 3538
rect 42720 921 42748 5714
rect 42800 5228 42852 5234
rect 42800 5170 42852 5176
rect 42812 3738 42840 5170
rect 42996 4146 43024 17138
rect 43088 16574 43116 19858
rect 43180 17610 43208 38898
rect 43260 37936 43312 37942
rect 43260 37878 43312 37884
rect 43272 36922 43300 37878
rect 43260 36916 43312 36922
rect 43260 36858 43312 36864
rect 43260 35692 43312 35698
rect 43260 35634 43312 35640
rect 43272 35601 43300 35634
rect 43258 35592 43314 35601
rect 43258 35527 43314 35536
rect 43272 35494 43300 35527
rect 43260 35488 43312 35494
rect 43260 35430 43312 35436
rect 43364 30258 43392 40446
rect 43444 39364 43496 39370
rect 43444 39306 43496 39312
rect 43456 39098 43484 39306
rect 43444 39092 43496 39098
rect 43444 39034 43496 39040
rect 43548 35578 43576 42162
rect 43916 41750 43944 42162
rect 43996 42016 44048 42022
rect 43996 41958 44048 41964
rect 43904 41744 43956 41750
rect 43904 41686 43956 41692
rect 44008 41682 44036 41958
rect 44192 41682 44220 43046
rect 43996 41676 44048 41682
rect 43996 41618 44048 41624
rect 44180 41676 44232 41682
rect 44180 41618 44232 41624
rect 44468 41478 44496 45200
rect 44456 41472 44508 41478
rect 44456 41414 44508 41420
rect 44180 40928 44232 40934
rect 44180 40870 44232 40876
rect 44192 40594 44220 40870
rect 44180 40588 44232 40594
rect 44180 40530 44232 40536
rect 44180 39840 44232 39846
rect 44180 39782 44232 39788
rect 44192 39506 44220 39782
rect 44180 39500 44232 39506
rect 44180 39442 44232 39448
rect 44180 38752 44232 38758
rect 44180 38694 44232 38700
rect 44192 38418 44220 38694
rect 44180 38412 44232 38418
rect 44180 38354 44232 38360
rect 43628 38276 43680 38282
rect 43628 38218 43680 38224
rect 43640 38010 43668 38218
rect 43628 38004 43680 38010
rect 43628 37946 43680 37952
rect 43720 37868 43772 37874
rect 43720 37810 43772 37816
rect 43732 37670 43760 37810
rect 43720 37664 43772 37670
rect 43720 37606 43772 37612
rect 43456 35550 43576 35578
rect 43456 33522 43484 35550
rect 43628 35012 43680 35018
rect 43628 34954 43680 34960
rect 43640 34746 43668 34954
rect 43628 34740 43680 34746
rect 43628 34682 43680 34688
rect 43732 34626 43760 37606
rect 43812 37120 43864 37126
rect 43812 37062 43864 37068
rect 43824 36786 43852 37062
rect 43812 36780 43864 36786
rect 43812 36722 43864 36728
rect 44180 36576 44232 36582
rect 44180 36518 44232 36524
rect 44192 36242 44220 36518
rect 44180 36236 44232 36242
rect 44180 36178 44232 36184
rect 43996 36100 44048 36106
rect 43996 36042 44048 36048
rect 44008 35834 44036 36042
rect 43996 35828 44048 35834
rect 43996 35770 44048 35776
rect 44180 35488 44232 35494
rect 44180 35430 44232 35436
rect 44192 35154 44220 35430
rect 44180 35148 44232 35154
rect 44180 35090 44232 35096
rect 43640 34610 43760 34626
rect 43628 34604 43760 34610
rect 43680 34598 43760 34604
rect 43628 34546 43680 34552
rect 43536 33924 43588 33930
rect 43536 33866 43588 33872
rect 43548 33658 43576 33866
rect 43536 33652 43588 33658
rect 43536 33594 43588 33600
rect 43444 33516 43496 33522
rect 43444 33458 43496 33464
rect 43352 30252 43404 30258
rect 43352 30194 43404 30200
rect 43364 29850 43392 30194
rect 43352 29844 43404 29850
rect 43352 29786 43404 29792
rect 43456 28558 43484 33458
rect 43444 28552 43496 28558
rect 43444 28494 43496 28500
rect 43640 26234 43668 34546
rect 44086 34096 44142 34105
rect 44086 34031 44088 34040
rect 44140 34031 44142 34040
rect 44088 34002 44140 34008
rect 44086 33416 44142 33425
rect 44086 33351 44142 33360
rect 44100 32978 44128 33351
rect 44088 32972 44140 32978
rect 44088 32914 44140 32920
rect 44086 30696 44142 30705
rect 43720 30660 43772 30666
rect 44086 30631 44088 30640
rect 43720 30602 43772 30608
rect 44140 30631 44142 30640
rect 44088 30602 44140 30608
rect 43732 29306 43760 30602
rect 43996 30048 44048 30054
rect 43996 29990 44048 29996
rect 44180 30048 44232 30054
rect 44180 29990 44232 29996
rect 44008 29714 44036 29990
rect 44192 29714 44220 29990
rect 43996 29708 44048 29714
rect 43996 29650 44048 29656
rect 44180 29708 44232 29714
rect 44180 29650 44232 29656
rect 43720 29300 43772 29306
rect 43720 29242 43772 29248
rect 43996 28416 44048 28422
rect 43996 28358 44048 28364
rect 44008 27538 44036 28358
rect 44180 27872 44232 27878
rect 44180 27814 44232 27820
rect 44192 27538 44220 27814
rect 43996 27532 44048 27538
rect 43996 27474 44048 27480
rect 44180 27532 44232 27538
rect 44180 27474 44232 27480
rect 43904 26376 43956 26382
rect 43904 26318 43956 26324
rect 43548 26206 43668 26234
rect 43260 24812 43312 24818
rect 43260 24754 43312 24760
rect 43272 23730 43300 24754
rect 43352 24608 43404 24614
rect 43352 24550 43404 24556
rect 43364 24274 43392 24550
rect 43352 24268 43404 24274
rect 43352 24210 43404 24216
rect 43352 23860 43404 23866
rect 43352 23802 43404 23808
rect 43260 23724 43312 23730
rect 43260 23666 43312 23672
rect 43272 18902 43300 23666
rect 43260 18896 43312 18902
rect 43260 18838 43312 18844
rect 43364 18290 43392 23802
rect 43444 23044 43496 23050
rect 43444 22986 43496 22992
rect 43456 22778 43484 22986
rect 43444 22772 43496 22778
rect 43444 22714 43496 22720
rect 43444 18692 43496 18698
rect 43444 18634 43496 18640
rect 43456 18426 43484 18634
rect 43444 18420 43496 18426
rect 43444 18362 43496 18368
rect 43352 18284 43404 18290
rect 43352 18226 43404 18232
rect 43168 17604 43220 17610
rect 43168 17546 43220 17552
rect 43088 16546 43208 16574
rect 42984 4140 43036 4146
rect 42984 4082 43036 4088
rect 42890 4040 42946 4049
rect 42890 3975 42946 3984
rect 42800 3732 42852 3738
rect 42800 3674 42852 3680
rect 42904 3466 42932 3975
rect 42892 3460 42944 3466
rect 42892 3402 42944 3408
rect 42904 3058 42932 3402
rect 42984 3188 43036 3194
rect 42984 3130 43036 3136
rect 42892 3052 42944 3058
rect 42892 2994 42944 3000
rect 42996 2650 43024 3130
rect 42984 2644 43036 2650
rect 42984 2586 43036 2592
rect 42706 912 42762 921
rect 42706 847 42762 856
rect 43180 800 43208 16546
rect 43260 16108 43312 16114
rect 43260 16050 43312 16056
rect 43272 6914 43300 16050
rect 43364 10674 43392 18226
rect 43548 16574 43576 26206
rect 43916 25362 43944 26318
rect 44180 25696 44232 25702
rect 44180 25638 44232 25644
rect 43904 25356 43956 25362
rect 43904 25298 43956 25304
rect 44088 25356 44140 25362
rect 44088 25298 44140 25304
rect 43996 25152 44048 25158
rect 43996 25094 44048 25100
rect 44008 24818 44036 25094
rect 43720 24812 43772 24818
rect 43720 24754 43772 24760
rect 43996 24812 44048 24818
rect 43996 24754 44048 24760
rect 43628 20256 43680 20262
rect 43628 20198 43680 20204
rect 43640 17882 43668 20198
rect 43732 19446 43760 24754
rect 44100 24585 44128 25298
rect 44086 24576 44142 24585
rect 44086 24511 44142 24520
rect 44192 24274 44220 25638
rect 44180 24268 44232 24274
rect 44180 24210 44232 24216
rect 44180 23520 44232 23526
rect 44180 23462 44232 23468
rect 44192 23186 44220 23462
rect 44180 23180 44232 23186
rect 44180 23122 44232 23128
rect 44086 21176 44142 21185
rect 44086 21111 44142 21120
rect 44100 21010 44128 21111
rect 44088 21004 44140 21010
rect 44088 20946 44140 20952
rect 43720 19440 43772 19446
rect 43720 19382 43772 19388
rect 43628 17876 43680 17882
rect 43628 17818 43680 17824
rect 43548 16546 43668 16574
rect 43444 15904 43496 15910
rect 43444 15846 43496 15852
rect 43456 14346 43484 15846
rect 43444 14340 43496 14346
rect 43444 14282 43496 14288
rect 43536 13728 43588 13734
rect 43536 13670 43588 13676
rect 43548 13258 43576 13670
rect 43536 13252 43588 13258
rect 43536 13194 43588 13200
rect 43444 12164 43496 12170
rect 43444 12106 43496 12112
rect 43456 11898 43484 12106
rect 43444 11892 43496 11898
rect 43444 11834 43496 11840
rect 43352 10668 43404 10674
rect 43352 10610 43404 10616
rect 43640 7410 43668 16546
rect 43732 13938 43760 19382
rect 44180 19168 44232 19174
rect 44180 19110 44232 19116
rect 44192 18834 44220 19110
rect 44180 18828 44232 18834
rect 44180 18770 44232 18776
rect 43996 16992 44048 16998
rect 43996 16934 44048 16940
rect 44180 16992 44232 16998
rect 44180 16934 44232 16940
rect 44008 16658 44036 16934
rect 44192 16658 44220 16934
rect 43996 16652 44048 16658
rect 43996 16594 44048 16600
rect 44180 16652 44232 16658
rect 44180 16594 44232 16600
rect 44086 16416 44142 16425
rect 44086 16351 44142 16360
rect 43996 15428 44048 15434
rect 43996 15370 44048 15376
rect 44008 15162 44036 15370
rect 43996 15156 44048 15162
rect 43996 15098 44048 15104
rect 43904 15020 43956 15026
rect 43904 14962 43956 14968
rect 43916 14618 43944 14962
rect 43904 14612 43956 14618
rect 43904 14554 43956 14560
rect 43720 13932 43772 13938
rect 43720 13874 43772 13880
rect 43732 12850 43760 13874
rect 43720 12844 43772 12850
rect 43720 12786 43772 12792
rect 43720 11212 43772 11218
rect 43720 11154 43772 11160
rect 43732 10985 43760 11154
rect 43718 10976 43774 10985
rect 43718 10911 43774 10920
rect 43628 7404 43680 7410
rect 43628 7346 43680 7352
rect 43272 6886 43392 6914
rect 43364 4146 43392 6886
rect 43628 5024 43680 5030
rect 43628 4966 43680 4972
rect 43640 4758 43668 4966
rect 43628 4752 43680 4758
rect 43628 4694 43680 4700
rect 43352 4140 43404 4146
rect 43352 4082 43404 4088
rect 43364 2582 43392 4082
rect 43444 3936 43496 3942
rect 43444 3878 43496 3884
rect 43536 3936 43588 3942
rect 43536 3878 43588 3884
rect 43352 2576 43404 2582
rect 43352 2518 43404 2524
rect 43456 2514 43484 3878
rect 43444 2508 43496 2514
rect 43444 2450 43496 2456
rect 43548 2446 43576 3878
rect 43916 3534 43944 14554
rect 44100 14482 44128 16351
rect 44180 15904 44232 15910
rect 44180 15846 44232 15852
rect 44192 15570 44220 15846
rect 44180 15564 44232 15570
rect 44180 15506 44232 15512
rect 44088 14476 44140 14482
rect 44088 14418 44140 14424
rect 44086 13696 44142 13705
rect 44086 13631 44142 13640
rect 44100 13394 44128 13631
rect 44088 13388 44140 13394
rect 44088 13330 44140 13336
rect 44180 12232 44232 12238
rect 44180 12174 44232 12180
rect 44192 11762 44220 12174
rect 44180 11756 44232 11762
rect 44180 11698 44232 11704
rect 44180 11144 44232 11150
rect 44180 11086 44232 11092
rect 43996 11076 44048 11082
rect 43996 11018 44048 11024
rect 44008 10810 44036 11018
rect 43996 10804 44048 10810
rect 43996 10746 44048 10752
rect 44192 10674 44220 11086
rect 44180 10668 44232 10674
rect 44180 10610 44232 10616
rect 45100 8900 45152 8906
rect 45100 8842 45152 8848
rect 44180 7880 44232 7886
rect 44180 7822 44232 7828
rect 44192 7585 44220 7822
rect 44178 7576 44234 7585
rect 44178 7511 44234 7520
rect 43996 7200 44048 7206
rect 43996 7142 44048 7148
rect 44008 6866 44036 7142
rect 43996 6860 44048 6866
rect 43996 6802 44048 6808
rect 44180 6792 44232 6798
rect 44180 6734 44232 6740
rect 44192 6322 44220 6734
rect 44180 6316 44232 6322
rect 44180 6258 44232 6264
rect 44180 5704 44232 5710
rect 44180 5646 44232 5652
rect 43996 5636 44048 5642
rect 43996 5578 44048 5584
rect 44008 3738 44036 5578
rect 44086 4856 44142 4865
rect 44086 4791 44142 4800
rect 44100 4690 44128 4791
rect 44088 4684 44140 4690
rect 44088 4626 44140 4632
rect 43996 3732 44048 3738
rect 43996 3674 44048 3680
rect 43904 3528 43956 3534
rect 43904 3470 43956 3476
rect 44192 3058 44220 5646
rect 44180 3052 44232 3058
rect 44180 2994 44232 3000
rect 43812 2848 43864 2854
rect 43812 2790 43864 2796
rect 43536 2440 43588 2446
rect 43536 2382 43588 2388
rect 43824 800 43852 2790
rect 45112 800 45140 8842
rect 41510 96 41566 105
rect 41432 54 41510 82
rect 41510 31 41566 40
rect 42494 0 42606 800
rect 43138 0 43250 800
rect 43782 0 43894 800
rect 45070 0 45182 800
rect 45714 0 45826 800
<< via2 >>
rect 1858 42880 1914 42936
rect 2870 44920 2926 44976
rect 2962 43560 3018 43616
rect 2870 42200 2926 42256
rect 1398 37440 1454 37496
rect 1398 23180 1454 23216
rect 1398 23160 1400 23180
rect 1400 23160 1452 23180
rect 1452 23160 1454 23180
rect 1398 10240 1454 10296
rect 2778 40160 2834 40216
rect 2778 29960 2834 30016
rect 2962 22516 2964 22536
rect 2964 22516 3016 22536
rect 3016 22516 3018 22536
rect 2962 22480 3018 22516
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 3330 38120 3386 38176
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 2778 20440 2834 20496
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 2962 18400 3018 18456
rect 2778 17076 2780 17096
rect 2780 17076 2832 17096
rect 2832 17076 2834 17096
rect 2778 17040 2834 17076
rect 2778 15680 2834 15736
rect 2778 14320 2834 14376
rect 2778 12960 2834 13016
rect 2870 9560 2926 9616
rect 2778 8880 2834 8936
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 3974 6840 4030 6896
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 2778 6196 2780 6216
rect 2780 6196 2832 6216
rect 2832 6196 2834 6216
rect 2778 6160 2834 6196
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 2778 4800 2834 4856
rect 2778 4120 2834 4176
rect 1398 3476 1400 3496
rect 1400 3476 1452 3496
rect 1452 3476 1454 3496
rect 1398 3440 1454 3476
rect 2778 1400 2834 1456
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 5906 40432 5962 40488
rect 3422 2080 3478 2136
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 8206 3576 8262 3632
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19338 37848 19394 37904
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19522 37868 19578 37904
rect 19522 37848 19524 37868
rect 19524 37848 19576 37868
rect 19576 37848 19578 37868
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 20626 27512 20682 27568
rect 24122 40432 24178 40488
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 25318 31084 25320 31104
rect 25320 31084 25372 31104
rect 25372 31084 25374 31104
rect 25318 31048 25374 31084
rect 25870 24676 25926 24712
rect 25870 24656 25872 24676
rect 25872 24656 25924 24676
rect 25924 24656 25926 24676
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 41786 43560 41842 43616
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 31114 24692 31116 24712
rect 31116 24692 31168 24712
rect 31168 24692 31170 24712
rect 31114 24656 31170 24692
rect 33322 29280 33378 29336
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 35990 29280 36046 29336
rect 41510 41520 41566 41576
rect 42522 44920 42578 44976
rect 42614 42236 42616 42256
rect 42616 42236 42668 42256
rect 42668 42236 42670 42256
rect 42614 42200 42670 42236
rect 42706 39500 42762 39536
rect 42706 39480 42708 39500
rect 42708 39480 42760 39500
rect 42760 39480 42762 39500
rect 42706 38120 42762 38176
rect 42614 36760 42670 36816
rect 41418 25880 41474 25936
rect 41418 21800 41474 21856
rect 38014 14184 38070 14240
rect 38566 14220 38568 14240
rect 38568 14220 38620 14240
rect 38620 14220 38622 14240
rect 38566 14184 38622 14220
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 24766 3576 24822 3632
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 42706 36080 42762 36136
rect 42706 35400 42762 35456
rect 42706 29960 42762 30016
rect 42706 27240 42762 27296
rect 42706 25200 42762 25256
rect 42706 23180 42762 23216
rect 42706 23160 42708 23180
rect 42708 23160 42760 23180
rect 42760 23160 42762 23180
rect 42614 19760 42670 19816
rect 42706 19080 42762 19136
rect 42338 17040 42394 17096
rect 42614 15680 42670 15736
rect 41418 12960 41474 13016
rect 42706 11600 42762 11656
rect 42706 6160 42762 6216
rect 41418 2080 41474 2136
rect 43258 35536 43314 35592
rect 44086 34060 44142 34096
rect 44086 34040 44088 34060
rect 44088 34040 44140 34060
rect 44140 34040 44142 34060
rect 44086 33360 44142 33416
rect 44086 30660 44142 30696
rect 44086 30640 44088 30660
rect 44088 30640 44140 30660
rect 44140 30640 44142 30660
rect 42890 3984 42946 4040
rect 42706 856 42762 912
rect 44086 24520 44142 24576
rect 44086 21120 44142 21176
rect 44086 16360 44142 16416
rect 43718 10920 43774 10976
rect 44086 13640 44142 13696
rect 44178 7520 44234 7576
rect 44086 4800 44142 4856
rect 41510 40 41566 96
<< metal3 >>
rect 0 45508 800 45748
rect 0 44978 800 45068
rect 2865 44978 2931 44981
rect 0 44976 2931 44978
rect 0 44920 2870 44976
rect 2926 44920 2931 44976
rect 0 44918 2931 44920
rect 0 44828 800 44918
rect 2865 44915 2931 44918
rect 42517 44978 42583 44981
rect 45200 44978 46000 45068
rect 42517 44976 46000 44978
rect 42517 44920 42522 44976
rect 42578 44920 46000 44976
rect 42517 44918 46000 44920
rect 42517 44915 42583 44918
rect 45200 44828 46000 44918
rect 45200 44148 46000 44388
rect 0 43618 800 43708
rect 2957 43618 3023 43621
rect 0 43616 3023 43618
rect 0 43560 2962 43616
rect 3018 43560 3023 43616
rect 0 43558 3023 43560
rect 0 43468 800 43558
rect 2957 43555 3023 43558
rect 41781 43618 41847 43621
rect 45200 43618 46000 43708
rect 41781 43616 46000 43618
rect 41781 43560 41786 43616
rect 41842 43560 46000 43616
rect 41781 43558 46000 43560
rect 41781 43555 41847 43558
rect 19568 43552 19888 43553
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 43487 19888 43488
rect 45200 43468 46000 43558
rect 0 42938 800 43028
rect 4208 43008 4528 43009
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 42943 4528 42944
rect 34928 43008 35248 43009
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 42943 35248 42944
rect 1853 42938 1919 42941
rect 0 42936 1919 42938
rect 0 42880 1858 42936
rect 1914 42880 1919 42936
rect 0 42878 1919 42880
rect 0 42788 800 42878
rect 1853 42875 1919 42878
rect 19568 42464 19888 42465
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 42399 19888 42400
rect 0 42258 800 42348
rect 2865 42258 2931 42261
rect 0 42256 2931 42258
rect 0 42200 2870 42256
rect 2926 42200 2931 42256
rect 0 42198 2931 42200
rect 0 42108 800 42198
rect 2865 42195 2931 42198
rect 42609 42258 42675 42261
rect 45200 42258 46000 42348
rect 42609 42256 46000 42258
rect 42609 42200 42614 42256
rect 42670 42200 46000 42256
rect 42609 42198 46000 42200
rect 42609 42195 42675 42198
rect 45200 42108 46000 42198
rect 4208 41920 4528 41921
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 41855 4528 41856
rect 34928 41920 35248 41921
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 41855 35248 41856
rect 41505 41578 41571 41581
rect 45200 41578 46000 41668
rect 41505 41576 46000 41578
rect 41505 41520 41510 41576
rect 41566 41520 46000 41576
rect 41505 41518 46000 41520
rect 41505 41515 41571 41518
rect 45200 41428 46000 41518
rect 19568 41376 19888 41377
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 41311 19888 41312
rect 0 40748 800 40988
rect 4208 40832 4528 40833
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 40767 4528 40768
rect 34928 40832 35248 40833
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 40767 35248 40768
rect 45200 40748 46000 40988
rect 5901 40490 5967 40493
rect 24117 40490 24183 40493
rect 5901 40488 24183 40490
rect 5901 40432 5906 40488
rect 5962 40432 24122 40488
rect 24178 40432 24183 40488
rect 5901 40430 24183 40432
rect 5901 40427 5967 40430
rect 24117 40427 24183 40430
rect 0 40218 800 40308
rect 19568 40288 19888 40289
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 40223 19888 40224
rect 2773 40218 2839 40221
rect 0 40216 2839 40218
rect 0 40160 2778 40216
rect 2834 40160 2839 40216
rect 0 40158 2839 40160
rect 0 40068 800 40158
rect 2773 40155 2839 40158
rect 4208 39744 4528 39745
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 39679 4528 39680
rect 34928 39744 35248 39745
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 39679 35248 39680
rect 0 39388 800 39628
rect 42701 39538 42767 39541
rect 45200 39538 46000 39628
rect 42701 39536 46000 39538
rect 42701 39480 42706 39536
rect 42762 39480 46000 39536
rect 42701 39478 46000 39480
rect 42701 39475 42767 39478
rect 45200 39388 46000 39478
rect 19568 39200 19888 39201
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 39135 19888 39136
rect 45200 38708 46000 38948
rect 4208 38656 4528 38657
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 38591 4528 38592
rect 34928 38656 35248 38657
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 38591 35248 38592
rect 0 38178 800 38268
rect 3325 38178 3391 38181
rect 0 38176 3391 38178
rect 0 38120 3330 38176
rect 3386 38120 3391 38176
rect 0 38118 3391 38120
rect 0 38028 800 38118
rect 3325 38115 3391 38118
rect 42701 38178 42767 38181
rect 45200 38178 46000 38268
rect 42701 38176 46000 38178
rect 42701 38120 42706 38176
rect 42762 38120 46000 38176
rect 42701 38118 46000 38120
rect 42701 38115 42767 38118
rect 19568 38112 19888 38113
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 38047 19888 38048
rect 45200 38028 46000 38118
rect 19333 37906 19399 37909
rect 19517 37906 19583 37909
rect 19333 37904 19583 37906
rect 19333 37848 19338 37904
rect 19394 37848 19522 37904
rect 19578 37848 19583 37904
rect 19333 37846 19583 37848
rect 19333 37843 19399 37846
rect 19517 37843 19583 37846
rect 0 37498 800 37588
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 1393 37498 1459 37501
rect 0 37496 1459 37498
rect 0 37440 1398 37496
rect 1454 37440 1459 37496
rect 0 37438 1459 37440
rect 0 37348 800 37438
rect 1393 37435 1459 37438
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 0 36668 800 36908
rect 42609 36818 42675 36821
rect 45200 36818 46000 36908
rect 42609 36816 46000 36818
rect 42609 36760 42614 36816
rect 42670 36760 46000 36816
rect 42609 36758 46000 36760
rect 42609 36755 42675 36758
rect 45200 36668 46000 36758
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 42701 36138 42767 36141
rect 45200 36138 46000 36228
rect 42701 36136 46000 36138
rect 42701 36080 42706 36136
rect 42762 36080 46000 36136
rect 42701 36078 46000 36080
rect 42701 36075 42767 36078
rect 45200 35988 46000 36078
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 0 35308 800 35548
rect 43110 35532 43116 35596
rect 43180 35594 43186 35596
rect 43253 35594 43319 35597
rect 43180 35592 43319 35594
rect 43180 35536 43258 35592
rect 43314 35536 43319 35592
rect 43180 35534 43319 35536
rect 43180 35532 43186 35534
rect 43253 35531 43319 35534
rect 42701 35458 42767 35461
rect 45200 35458 46000 35548
rect 42701 35456 46000 35458
rect 42701 35400 42706 35456
rect 42762 35400 46000 35456
rect 42701 35398 46000 35400
rect 42701 35395 42767 35398
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 45200 35308 46000 35398
rect 0 34628 800 34868
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 0 33948 800 34188
rect 44081 34098 44147 34101
rect 45200 34098 46000 34188
rect 44081 34096 46000 34098
rect 44081 34040 44086 34096
rect 44142 34040 46000 34096
rect 44081 34038 46000 34040
rect 44081 34035 44147 34038
rect 45200 33948 46000 34038
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 44081 33418 44147 33421
rect 45200 33418 46000 33508
rect 44081 33416 46000 33418
rect 44081 33360 44086 33416
rect 44142 33360 46000 33416
rect 44081 33358 46000 33360
rect 44081 33355 44147 33358
rect 45200 33268 46000 33358
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 0 32588 800 32828
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 45200 32588 46000 32828
rect 0 31908 800 32148
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 0 31228 800 31468
rect 45200 31228 46000 31468
rect 24894 31044 24900 31108
rect 24964 31106 24970 31108
rect 25313 31106 25379 31109
rect 24964 31104 25379 31106
rect 24964 31048 25318 31104
rect 25374 31048 25379 31104
rect 24964 31046 25379 31048
rect 24964 31044 24970 31046
rect 25313 31043 25379 31046
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 44081 30698 44147 30701
rect 45200 30698 46000 30788
rect 44081 30696 46000 30698
rect 44081 30640 44086 30696
rect 44142 30640 46000 30696
rect 44081 30638 46000 30640
rect 44081 30635 44147 30638
rect 45200 30548 46000 30638
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 0 30018 800 30108
rect 2773 30018 2839 30021
rect 0 30016 2839 30018
rect 0 29960 2778 30016
rect 2834 29960 2839 30016
rect 0 29958 2839 29960
rect 0 29868 800 29958
rect 2773 29955 2839 29958
rect 42701 30018 42767 30021
rect 45200 30018 46000 30108
rect 42701 30016 46000 30018
rect 42701 29960 42706 30016
rect 42762 29960 46000 30016
rect 42701 29958 46000 29960
rect 42701 29955 42767 29958
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 45200 29868 46000 29958
rect 0 29188 800 29428
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 33317 29338 33383 29341
rect 35985 29338 36051 29341
rect 33317 29336 36051 29338
rect 33317 29280 33322 29336
rect 33378 29280 35990 29336
rect 36046 29280 36051 29336
rect 33317 29278 36051 29280
rect 33317 29275 33383 29278
rect 35985 29275 36051 29278
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 0 28508 800 28748
rect 45200 28508 46000 28748
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 45200 27828 46000 28068
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 20621 27570 20687 27573
rect 24894 27570 24900 27572
rect 20621 27568 24900 27570
rect 20621 27512 20626 27568
rect 20682 27512 24900 27568
rect 20621 27510 24900 27512
rect 20621 27507 20687 27510
rect 24894 27508 24900 27510
rect 24964 27508 24970 27572
rect 0 27148 800 27388
rect 42701 27298 42767 27301
rect 45200 27298 46000 27388
rect 42701 27296 46000 27298
rect 42701 27240 42706 27296
rect 42762 27240 46000 27296
rect 42701 27238 46000 27240
rect 42701 27235 42767 27238
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 45200 27148 46000 27238
rect 0 26468 800 26708
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 0 25788 800 26028
rect 41413 25938 41479 25941
rect 45200 25938 46000 26028
rect 41413 25936 46000 25938
rect 41413 25880 41418 25936
rect 41474 25880 46000 25936
rect 41413 25878 46000 25880
rect 41413 25875 41479 25878
rect 45200 25788 46000 25878
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 42701 25258 42767 25261
rect 45200 25258 46000 25348
rect 42701 25256 46000 25258
rect 42701 25200 42706 25256
rect 42762 25200 46000 25256
rect 42701 25198 46000 25200
rect 42701 25195 42767 25198
rect 45200 25108 46000 25198
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 25865 24714 25931 24717
rect 31109 24714 31175 24717
rect 25865 24712 31175 24714
rect 0 24428 800 24668
rect 25865 24656 25870 24712
rect 25926 24656 31114 24712
rect 31170 24656 31175 24712
rect 25865 24654 31175 24656
rect 25865 24651 25931 24654
rect 31109 24651 31175 24654
rect 44081 24578 44147 24581
rect 45200 24578 46000 24668
rect 44081 24576 46000 24578
rect 44081 24520 44086 24576
rect 44142 24520 46000 24576
rect 44081 24518 46000 24520
rect 44081 24515 44147 24518
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 45200 24428 46000 24518
rect 0 23748 800 23988
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 0 23218 800 23308
rect 1393 23218 1459 23221
rect 0 23216 1459 23218
rect 0 23160 1398 23216
rect 1454 23160 1459 23216
rect 0 23158 1459 23160
rect 0 23068 800 23158
rect 1393 23155 1459 23158
rect 42701 23218 42767 23221
rect 45200 23218 46000 23308
rect 42701 23216 46000 23218
rect 42701 23160 42706 23216
rect 42762 23160 46000 23216
rect 42701 23158 46000 23160
rect 42701 23155 42767 23158
rect 45200 23068 46000 23158
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 0 22538 800 22628
rect 2957 22538 3023 22541
rect 0 22536 3023 22538
rect 0 22480 2962 22536
rect 3018 22480 3023 22536
rect 0 22478 3023 22480
rect 0 22388 800 22478
rect 2957 22475 3023 22478
rect 45200 22388 46000 22628
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 41413 21858 41479 21861
rect 45200 21858 46000 21948
rect 41413 21856 46000 21858
rect 41413 21800 41418 21856
rect 41474 21800 46000 21856
rect 41413 21798 46000 21800
rect 41413 21795 41479 21798
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 45200 21708 46000 21798
rect 0 21028 800 21268
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 44081 21178 44147 21181
rect 45200 21178 46000 21268
rect 44081 21176 46000 21178
rect 44081 21120 44086 21176
rect 44142 21120 46000 21176
rect 44081 21118 46000 21120
rect 44081 21115 44147 21118
rect 45200 21028 46000 21118
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 0 20498 800 20588
rect 2773 20498 2839 20501
rect 0 20496 2839 20498
rect 0 20440 2778 20496
rect 2834 20440 2839 20496
rect 0 20438 2839 20440
rect 0 20348 800 20438
rect 2773 20435 2839 20438
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 0 19668 800 19908
rect 42609 19818 42675 19821
rect 45200 19818 46000 19908
rect 42609 19816 46000 19818
rect 42609 19760 42614 19816
rect 42670 19760 46000 19816
rect 42609 19758 46000 19760
rect 42609 19755 42675 19758
rect 45200 19668 46000 19758
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 42701 19138 42767 19141
rect 45200 19138 46000 19228
rect 42701 19136 46000 19138
rect 42701 19080 42706 19136
rect 42762 19080 46000 19136
rect 42701 19078 46000 19080
rect 42701 19075 42767 19078
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 45200 18988 46000 19078
rect 0 18458 800 18548
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 2957 18458 3023 18461
rect 0 18456 3023 18458
rect 0 18400 2962 18456
rect 3018 18400 3023 18456
rect 0 18398 3023 18400
rect 0 18308 800 18398
rect 2957 18395 3023 18398
rect 45200 18308 46000 18548
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 0 17628 800 17868
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 0 17098 800 17188
rect 2773 17098 2839 17101
rect 0 17096 2839 17098
rect 0 17040 2778 17096
rect 2834 17040 2839 17096
rect 0 17038 2839 17040
rect 0 16948 800 17038
rect 2773 17035 2839 17038
rect 42333 17098 42399 17101
rect 45200 17098 46000 17188
rect 42333 17096 46000 17098
rect 42333 17040 42338 17096
rect 42394 17040 46000 17096
rect 42333 17038 46000 17040
rect 42333 17035 42399 17038
rect 45200 16948 46000 17038
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 44081 16418 44147 16421
rect 45200 16418 46000 16508
rect 44081 16416 46000 16418
rect 44081 16360 44086 16416
rect 44142 16360 46000 16416
rect 44081 16358 46000 16360
rect 44081 16355 44147 16358
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 45200 16268 46000 16358
rect 0 15738 800 15828
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 2773 15738 2839 15741
rect 0 15736 2839 15738
rect 0 15680 2778 15736
rect 2834 15680 2839 15736
rect 0 15678 2839 15680
rect 0 15588 800 15678
rect 2773 15675 2839 15678
rect 42609 15738 42675 15741
rect 45200 15738 46000 15828
rect 42609 15736 46000 15738
rect 42609 15680 42614 15736
rect 42670 15680 46000 15736
rect 42609 15678 46000 15680
rect 42609 15675 42675 15678
rect 45200 15588 46000 15678
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 0 14908 800 15148
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 0 14378 800 14468
rect 2773 14378 2839 14381
rect 0 14376 2839 14378
rect 0 14320 2778 14376
rect 2834 14320 2839 14376
rect 0 14318 2839 14320
rect 0 14228 800 14318
rect 2773 14315 2839 14318
rect 38009 14242 38075 14245
rect 38561 14242 38627 14245
rect 38009 14240 38627 14242
rect 38009 14184 38014 14240
rect 38070 14184 38566 14240
rect 38622 14184 38627 14240
rect 45200 14228 46000 14468
rect 38009 14182 38627 14184
rect 38009 14179 38075 14182
rect 38561 14179 38627 14182
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 44081 13698 44147 13701
rect 45200 13698 46000 13788
rect 44081 13696 46000 13698
rect 44081 13640 44086 13696
rect 44142 13640 46000 13696
rect 44081 13638 46000 13640
rect 44081 13635 44147 13638
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 45200 13548 46000 13638
rect 0 13018 800 13108
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 2773 13018 2839 13021
rect 0 13016 2839 13018
rect 0 12960 2778 13016
rect 2834 12960 2839 13016
rect 0 12958 2839 12960
rect 0 12868 800 12958
rect 2773 12955 2839 12958
rect 41413 13018 41479 13021
rect 45200 13018 46000 13108
rect 41413 13016 46000 13018
rect 41413 12960 41418 13016
rect 41474 12960 46000 13016
rect 41413 12958 46000 12960
rect 41413 12955 41479 12958
rect 45200 12868 46000 12958
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 0 12188 800 12428
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 0 11508 800 11748
rect 42701 11658 42767 11661
rect 45200 11658 46000 11748
rect 42701 11656 46000 11658
rect 42701 11600 42706 11656
rect 42762 11600 46000 11656
rect 42701 11598 46000 11600
rect 42701 11595 42767 11598
rect 45200 11508 46000 11598
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 43713 10978 43779 10981
rect 45200 10978 46000 11068
rect 43713 10976 46000 10978
rect 43713 10920 43718 10976
rect 43774 10920 46000 10976
rect 43713 10918 46000 10920
rect 43713 10915 43779 10918
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 45200 10828 46000 10918
rect 0 10298 800 10388
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 1393 10298 1459 10301
rect 0 10296 1459 10298
rect 0 10240 1398 10296
rect 1454 10240 1459 10296
rect 0 10238 1459 10240
rect 0 10148 800 10238
rect 1393 10235 1459 10238
rect 45200 10148 46000 10388
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 0 9618 800 9708
rect 2865 9618 2931 9621
rect 0 9616 2931 9618
rect 0 9560 2870 9616
rect 2926 9560 2931 9616
rect 0 9558 2931 9560
rect 0 9468 800 9558
rect 2865 9555 2931 9558
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 0 8938 800 9028
rect 2773 8938 2839 8941
rect 0 8936 2839 8938
rect 0 8880 2778 8936
rect 2834 8880 2839 8936
rect 0 8878 2839 8880
rect 0 8788 800 8878
rect 2773 8875 2839 8878
rect 45200 8788 46000 9028
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 45200 8108 46000 8348
rect 0 7428 800 7668
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 44173 7578 44239 7581
rect 45200 7578 46000 7668
rect 44173 7576 46000 7578
rect 44173 7520 44178 7576
rect 44234 7520 46000 7576
rect 44173 7518 46000 7520
rect 44173 7515 44239 7518
rect 45200 7428 46000 7518
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 0 6898 800 6988
rect 3969 6898 4035 6901
rect 0 6896 4035 6898
rect 0 6840 3974 6896
rect 4030 6840 4035 6896
rect 0 6838 4035 6840
rect 0 6748 800 6838
rect 3969 6835 4035 6838
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 0 6218 800 6308
rect 2773 6218 2839 6221
rect 0 6216 2839 6218
rect 0 6160 2778 6216
rect 2834 6160 2839 6216
rect 0 6158 2839 6160
rect 0 6068 800 6158
rect 2773 6155 2839 6158
rect 42701 6218 42767 6221
rect 45200 6218 46000 6308
rect 42701 6216 46000 6218
rect 42701 6160 42706 6216
rect 42762 6160 46000 6216
rect 42701 6158 46000 6160
rect 42701 6155 42767 6158
rect 45200 6068 46000 6158
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 45200 5388 46000 5628
rect 0 4858 800 4948
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 2773 4858 2839 4861
rect 0 4856 2839 4858
rect 0 4800 2778 4856
rect 2834 4800 2839 4856
rect 0 4798 2839 4800
rect 0 4708 800 4798
rect 2773 4795 2839 4798
rect 44081 4858 44147 4861
rect 45200 4858 46000 4948
rect 44081 4856 46000 4858
rect 44081 4800 44086 4856
rect 44142 4800 46000 4856
rect 44081 4798 46000 4800
rect 44081 4795 44147 4798
rect 45200 4708 46000 4798
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 0 4178 800 4268
rect 2773 4178 2839 4181
rect 0 4176 2839 4178
rect 0 4120 2778 4176
rect 2834 4120 2839 4176
rect 0 4118 2839 4120
rect 0 4028 800 4118
rect 2773 4115 2839 4118
rect 42885 4042 42951 4045
rect 43110 4042 43116 4044
rect 42885 4040 43116 4042
rect 42885 3984 42890 4040
rect 42946 3984 43116 4040
rect 42885 3982 43116 3984
rect 42885 3979 42951 3982
rect 43110 3980 43116 3982
rect 43180 3980 43186 4044
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 8201 3634 8267 3637
rect 24761 3634 24827 3637
rect 8201 3632 24827 3634
rect 0 3498 800 3588
rect 8201 3576 8206 3632
rect 8262 3576 24766 3632
rect 24822 3576 24827 3632
rect 8201 3574 24827 3576
rect 8201 3571 8267 3574
rect 24761 3571 24827 3574
rect 1393 3498 1459 3501
rect 0 3496 1459 3498
rect 0 3440 1398 3496
rect 1454 3440 1459 3496
rect 0 3438 1459 3440
rect 0 3348 800 3438
rect 1393 3435 1459 3438
rect 45200 3348 46000 3588
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 45200 2668 46000 2908
rect 0 2138 800 2228
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 3417 2138 3483 2141
rect 0 2136 3483 2138
rect 0 2080 3422 2136
rect 3478 2080 3483 2136
rect 0 2078 3483 2080
rect 0 1988 800 2078
rect 3417 2075 3483 2078
rect 41413 2138 41479 2141
rect 45200 2138 46000 2228
rect 41413 2136 46000 2138
rect 41413 2080 41418 2136
rect 41474 2080 46000 2136
rect 41413 2078 46000 2080
rect 41413 2075 41479 2078
rect 45200 1988 46000 2078
rect 0 1458 800 1548
rect 2773 1458 2839 1461
rect 0 1456 2839 1458
rect 0 1400 2778 1456
rect 2834 1400 2839 1456
rect 0 1398 2839 1400
rect 0 1308 800 1398
rect 2773 1395 2839 1398
rect 42701 914 42767 917
rect 42701 912 42810 914
rect 0 628 800 868
rect 42701 856 42706 912
rect 42762 856 42810 912
rect 42701 851 42810 856
rect 42750 778 42810 851
rect 45200 778 46000 868
rect 42750 718 46000 778
rect 45200 628 46000 718
rect 41505 98 41571 101
rect 45200 98 46000 188
rect 41505 96 46000 98
rect 41505 40 41510 96
rect 41566 40 46000 96
rect 41505 38 46000 40
rect 41505 35 41571 38
rect 45200 -52 46000 38
<< via3 >>
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 43116 35532 43180 35596
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 24900 31044 24964 31108
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 24900 27508 24964 27572
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 43116 3980 43180 4044
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 43008 4528 43568
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 43552 19888 43568
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 34928 43008 35248 43568
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 43115 35596 43181 35597
rect 43115 35532 43116 35596
rect 43180 35532 43181 35596
rect 43115 35531 43181 35532
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 24899 31108 24965 31109
rect 24899 31044 24900 31108
rect 24964 31044 24965 31108
rect 24899 31043 24965 31044
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 24902 27573 24962 31043
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 24899 27572 24965 27573
rect 24899 27508 24900 27572
rect 24964 27508 24965 27572
rect 24899 27507 24965 27508
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 43118 4045 43178 35531
rect 43115 4044 43181 4045
rect 43115 3980 43116 4044
rect 43180 3980 43181 4044
rect 43115 3979 43181 3980
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__decap_4  FILLER_0_24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5704 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78
timestamp 1644511149
transform 1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_97
timestamp 1644511149
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 1644511149
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_153
timestamp 1644511149
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1644511149
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_192
timestamp 1644511149
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_209
timestamp 1644511149
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1644511149
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_225 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_233
timestamp 1644511149
transform 1 0 22540 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_239
timestamp 1644511149
transform 1 0 23092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_274
timestamp 1644511149
transform 1 0 26312 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_293
timestamp 1644511149
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1644511149
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_309
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_321
timestamp 1644511149
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1644511149
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_349
timestamp 1644511149
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1644511149
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_377
timestamp 1644511149
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1644511149
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_414
timestamp 1644511149
transform 1 0 39192 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_421
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_444
timestamp 1644511149
transform 1 0 41952 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_449
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_458
timestamp 1644511149
transform 1 0 43240 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_470
timestamp 1644511149
transform 1 0 44344 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_7
timestamp 1644511149
transform 1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_14
timestamp 1644511149
transform 1 0 2392 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_18
timestamp 1644511149
transform 1 0 2760 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_22
timestamp 1644511149
transform 1 0 3128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_47
timestamp 1644511149
transform 1 0 5428 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1644511149
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_60
timestamp 1644511149
transform 1 0 6624 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_66
timestamp 1644511149
transform 1 0 7176 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_88
timestamp 1644511149
transform 1 0 9200 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_100
timestamp 1644511149
transform 1 0 10304 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_134
timestamp 1644511149
transform 1 0 13432 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_146
timestamp 1644511149
transform 1 0 14536 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1644511149
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1644511149
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_175
timestamp 1644511149
transform 1 0 17204 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_187
timestamp 1644511149
transform 1 0 18308 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_191
timestamp 1644511149
transform 1 0 18676 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_213
timestamp 1644511149
transform 1 0 20700 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_221
timestamp 1644511149
transform 1 0 21436 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_249
timestamp 1644511149
transform 1 0 24012 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_274
timestamp 1644511149
transform 1 0 26312 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_293
timestamp 1644511149
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_326
timestamp 1644511149
transform 1 0 31096 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_334
timestamp 1644511149
transform 1 0 31832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_349
timestamp 1644511149
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_361
timestamp 1644511149
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_373
timestamp 1644511149
transform 1 0 35420 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_379
timestamp 1644511149
transform 1 0 35972 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_388
timestamp 1644511149
transform 1 0 36800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_393
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_397
timestamp 1644511149
transform 1 0 37628 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_419
timestamp 1644511149
transform 1 0 39652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_444
timestamp 1644511149
transform 1 0 41952 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_449
timestamp 1644511149
transform 1 0 42412 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_456
timestamp 1644511149
transform 1 0 43056 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_465
timestamp 1644511149
transform 1 0 43884 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1644511149
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_29
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_38
timestamp 1644511149
transform 1 0 4600 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_67
timestamp 1644511149
transform 1 0 7268 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_75
timestamp 1644511149
transform 1 0 8004 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_79
timestamp 1644511149
transform 1 0 8372 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1644511149
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_109
timestamp 1644511149
transform 1 0 11132 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_117
timestamp 1644511149
transform 1 0 11868 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_122
timestamp 1644511149
transform 1 0 12328 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_129
timestamp 1644511149
transform 1 0 12972 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_137
timestamp 1644511149
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_153
timestamp 1644511149
transform 1 0 15180 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_177
timestamp 1644511149
transform 1 0 17388 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_184
timestamp 1644511149
transform 1 0 18032 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_188
timestamp 1644511149
transform 1 0 18400 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1644511149
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_200
timestamp 1644511149
transform 1 0 19504 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_204
timestamp 1644511149
transform 1 0 19872 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_208
timestamp 1644511149
transform 1 0 20240 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_233
timestamp 1644511149
transform 1 0 22540 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_240
timestamp 1644511149
transform 1 0 23184 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_244
timestamp 1644511149
transform 1 0 23552 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_248
timestamp 1644511149
transform 1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_258
timestamp 1644511149
transform 1 0 24840 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_265
timestamp 1644511149
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_277
timestamp 1644511149
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_289
timestamp 1644511149
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_304
timestamp 1644511149
transform 1 0 29072 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_312
timestamp 1644511149
transform 1 0 29808 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_324
timestamp 1644511149
transform 1 0 30912 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_336
timestamp 1644511149
transform 1 0 32016 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_348
timestamp 1644511149
transform 1 0 33120 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_360
timestamp 1644511149
transform 1 0 34224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_373
timestamp 1644511149
transform 1 0 35420 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_396
timestamp 1644511149
transform 1 0 37536 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_402
timestamp 1644511149
transform 1 0 38088 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_406
timestamp 1644511149
transform 1 0 38456 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1644511149
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1644511149
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_421
timestamp 1644511149
transform 1 0 39836 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_426
timestamp 1644511149
transform 1 0 40296 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_433
timestamp 1644511149
transform 1 0 40940 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_462
timestamp 1644511149
transform 1 0 43608 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_469
timestamp 1644511149
transform 1 0 44252 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_7
timestamp 1644511149
transform 1 0 1748 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_11
timestamp 1644511149
transform 1 0 2116 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_36
timestamp 1644511149
transform 1 0 4416 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_44
timestamp 1644511149
transform 1 0 5152 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_49
timestamp 1644511149
transform 1 0 5612 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1644511149
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_60
timestamp 1644511149
transform 1 0 6624 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_71
timestamp 1644511149
transform 1 0 7636 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_83
timestamp 1644511149
transform 1 0 8740 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_92
timestamp 1644511149
transform 1 0 9568 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_104
timestamp 1644511149
transform 1 0 10672 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_119
timestamp 1644511149
transform 1 0 12052 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_126
timestamp 1644511149
transform 1 0 12696 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_138
timestamp 1644511149
transform 1 0 13800 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_150
timestamp 1644511149
transform 1 0 14904 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_156
timestamp 1644511149
transform 1 0 15456 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_160
timestamp 1644511149
transform 1 0 15824 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_181
timestamp 1644511149
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_193
timestamp 1644511149
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_205
timestamp 1644511149
transform 1 0 19964 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_213
timestamp 1644511149
transform 1 0 20700 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1644511149
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1644511149
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_237
timestamp 1644511149
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_252
timestamp 1644511149
transform 1 0 24288 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_264
timestamp 1644511149
transform 1 0 25392 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_276
timestamp 1644511149
transform 1 0 26496 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_305
timestamp 1644511149
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_317
timestamp 1644511149
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1644511149
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1644511149
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_349
timestamp 1644511149
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_361
timestamp 1644511149
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_373
timestamp 1644511149
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_388
timestamp 1644511149
transform 1 0 36800 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_396
timestamp 1644511149
transform 1 0 37536 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_403
timestamp 1644511149
transform 1 0 38180 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_409
timestamp 1644511149
transform 1 0 38732 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_431
timestamp 1644511149
transform 1 0 40756 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_439
timestamp 1644511149
transform 1 0 41492 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_444
timestamp 1644511149
transform 1 0 41952 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_452
timestamp 1644511149
transform 1 0 42688 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_458
timestamp 1644511149
transform 1 0 43240 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_462
timestamp 1644511149
transform 1 0 43608 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_469
timestamp 1644511149
transform 1 0 44252 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_10
timestamp 1644511149
transform 1 0 2024 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_17
timestamp 1644511149
transform 1 0 2668 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1644511149
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_60
timestamp 1644511149
transform 1 0 6624 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_72
timestamp 1644511149
transform 1 0 7728 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_97
timestamp 1644511149
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_109
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_121
timestamp 1644511149
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1644511149
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1644511149
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1644511149
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_209
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_221
timestamp 1644511149
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_233
timestamp 1644511149
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1644511149
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1644511149
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_277
timestamp 1644511149
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_289
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1644511149
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1644511149
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_345
timestamp 1644511149
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1644511149
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_389
timestamp 1644511149
transform 1 0 36892 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_393
timestamp 1644511149
transform 1 0 37260 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_415
timestamp 1644511149
transform 1 0 39284 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1644511149
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_421
timestamp 1644511149
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_433
timestamp 1644511149
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_445
timestamp 1644511149
transform 1 0 42044 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_469
timestamp 1644511149
transform 1 0 44252 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_30
timestamp 1644511149
transform 1 0 3864 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_37
timestamp 1644511149
transform 1 0 4508 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_44
timestamp 1644511149
transform 1 0 5152 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_193
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_205
timestamp 1644511149
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1644511149
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_249
timestamp 1644511149
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_261
timestamp 1644511149
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1644511149
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_373
timestamp 1644511149
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1644511149
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_405
timestamp 1644511149
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_417
timestamp 1644511149
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_429
timestamp 1644511149
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1644511149
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1644511149
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_449
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_456
timestamp 1644511149
transform 1 0 43056 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_5_465
timestamp 1644511149
transform 1 0 43884 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_6
timestamp 1644511149
transform 1 0 1656 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_13
timestamp 1644511149
transform 1 0 2300 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_17
timestamp 1644511149
transform 1 0 2668 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_21
timestamp 1644511149
transform 1 0 3036 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_32
timestamp 1644511149
transform 1 0 4048 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_39
timestamp 1644511149
transform 1 0 4692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_51
timestamp 1644511149
transform 1 0 5796 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_63
timestamp 1644511149
transform 1 0 6900 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_75
timestamp 1644511149
transform 1 0 8004 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_401
timestamp 1644511149
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1644511149
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1644511149
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_421
timestamp 1644511149
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_433
timestamp 1644511149
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_445
timestamp 1644511149
transform 1 0 42044 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_469
timestamp 1644511149
transform 1 0 44252 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1644511149
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1644511149
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_417
timestamp 1644511149
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_429
timestamp 1644511149
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1644511149
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1644511149
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_449
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_461
timestamp 1644511149
transform 1 0 43516 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_465
timestamp 1644511149
transform 1 0 43884 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_10
timestamp 1644511149
transform 1 0 2024 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_22
timestamp 1644511149
transform 1 0 3128 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_50
timestamp 1644511149
transform 1 0 5704 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_62
timestamp 1644511149
transform 1 0 6808 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_74
timestamp 1644511149
transform 1 0 7912 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1644511149
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_389
timestamp 1644511149
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_401
timestamp 1644511149
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1644511149
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1644511149
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_421
timestamp 1644511149
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_433
timestamp 1644511149
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_445
timestamp 1644511149
transform 1 0 42044 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_469
timestamp 1644511149
transform 1 0 44252 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_23
timestamp 1644511149
transform 1 0 3220 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_28
timestamp 1644511149
transform 1 0 3680 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_35
timestamp 1644511149
transform 1 0 4324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_47
timestamp 1644511149
transform 1 0 5428 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_193
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_205
timestamp 1644511149
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1644511149
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_317
timestamp 1644511149
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1644511149
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_361
timestamp 1644511149
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1644511149
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_417
timestamp 1644511149
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_429
timestamp 1644511149
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1644511149
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1644511149
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_449
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_464
timestamp 1644511149
transform 1 0 43792 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_472
timestamp 1644511149
transform 1 0 44528 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1644511149
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_209
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_221
timestamp 1644511149
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_233
timestamp 1644511149
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1644511149
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1644511149
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_345
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1644511149
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_401
timestamp 1644511149
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1644511149
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1644511149
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_433
timestamp 1644511149
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_445
timestamp 1644511149
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_457
timestamp 1644511149
transform 1 0 43148 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_469
timestamp 1644511149
transform 1 0 44252 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_30
timestamp 1644511149
transform 1 0 3864 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_42
timestamp 1644511149
transform 1 0 4968 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1644511149
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_205
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_213
timestamp 1644511149
transform 1 0 20700 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_219
timestamp 1644511149
transform 1 0 21252 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_233
timestamp 1644511149
transform 1 0 22540 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_251
timestamp 1644511149
transform 1 0 24196 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_263
timestamp 1644511149
transform 1 0 25300 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_275
timestamp 1644511149
transform 1 0 26404 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1644511149
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_373
timestamp 1644511149
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1644511149
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1644511149
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_417
timestamp 1644511149
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_429
timestamp 1644511149
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1644511149
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1644511149
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_449
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_461
timestamp 1644511149
transform 1 0 43516 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_465
timestamp 1644511149
transform 1 0 43884 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_10
timestamp 1644511149
transform 1 0 2024 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_17
timestamp 1644511149
transform 1 0 2668 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_25
timestamp 1644511149
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_177
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_205
timestamp 1644511149
transform 1 0 19964 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_213
timestamp 1644511149
transform 1 0 20700 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_231
timestamp 1644511149
transform 1 0 22356 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_241
timestamp 1644511149
transform 1 0 23276 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_249
timestamp 1644511149
transform 1 0 24012 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_277
timestamp 1644511149
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_289
timestamp 1644511149
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1644511149
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1644511149
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1644511149
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_433
timestamp 1644511149
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_445
timestamp 1644511149
transform 1 0 42044 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_469
timestamp 1644511149
transform 1 0 44252 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_30
timestamp 1644511149
transform 1 0 3864 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_42
timestamp 1644511149
transform 1 0 4968 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1644511149
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_177
timestamp 1644511149
transform 1 0 17388 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_182
timestamp 1644511149
transform 1 0 17848 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_190
timestamp 1644511149
transform 1 0 18584 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_214
timestamp 1644511149
transform 1 0 20792 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1644511149
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_241
timestamp 1644511149
transform 1 0 23276 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_248
timestamp 1644511149
transform 1 0 23920 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_256
timestamp 1644511149
transform 1 0 24656 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_260
timestamp 1644511149
transform 1 0 25024 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_267
timestamp 1644511149
transform 1 0 25668 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1644511149
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_305
timestamp 1644511149
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_317
timestamp 1644511149
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1644511149
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1644511149
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_417
timestamp 1644511149
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_429
timestamp 1644511149
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1644511149
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1644511149
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_449
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_456
timestamp 1644511149
transform 1 0 43056 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_468
timestamp 1644511149
transform 1 0 44160 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_472
timestamp 1644511149
transform 1 0 44528 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp 1644511149
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1644511149
transform 1 0 4048 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1644511149
transform 1 0 5152 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1644511149
transform 1 0 6256 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1644511149
transform 1 0 7360 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_80
timestamp 1644511149
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_173
timestamp 1644511149
transform 1 0 17020 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_192
timestamp 1644511149
transform 1 0 18768 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_205
timestamp 1644511149
transform 1 0 19964 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_217
timestamp 1644511149
transform 1 0 21068 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_225
timestamp 1644511149
transform 1 0 21804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_242
timestamp 1644511149
transform 1 0 23368 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1644511149
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_258
timestamp 1644511149
transform 1 0 24840 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_278
timestamp 1644511149
transform 1 0 26680 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_303
timestamp 1644511149
transform 1 0 28980 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1644511149
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_345
timestamp 1644511149
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1644511149
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1644511149
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1644511149
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_421
timestamp 1644511149
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_433
timestamp 1644511149
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_445
timestamp 1644511149
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_457
timestamp 1644511149
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_469
timestamp 1644511149
transform 1 0 44252 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_10
timestamp 1644511149
transform 1 0 2024 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_17
timestamp 1644511149
transform 1 0 2668 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_29
timestamp 1644511149
transform 1 0 3772 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_41
timestamp 1644511149
transform 1 0 4876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp 1644511149
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1644511149
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_177
timestamp 1644511149
transform 1 0 17388 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_182
timestamp 1644511149
transform 1 0 17848 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_186
timestamp 1644511149
transform 1 0 18216 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_192
timestamp 1644511149
transform 1 0 18768 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_204
timestamp 1644511149
transform 1 0 19872 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1644511149
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_246
timestamp 1644511149
transform 1 0 23736 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_255
timestamp 1644511149
transform 1 0 24564 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_259
timestamp 1644511149
transform 1 0 24932 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_276
timestamp 1644511149
transform 1 0 26496 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_297
timestamp 1644511149
transform 1 0 28428 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_317
timestamp 1644511149
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1644511149
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1644511149
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1644511149
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_417
timestamp 1644511149
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_429
timestamp 1644511149
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1644511149
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1644511149
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_449
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_457
timestamp 1644511149
transform 1 0 43148 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_462
timestamp 1644511149
transform 1 0 43608 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_469
timestamp 1644511149
transform 1 0 44252 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_7
timestamp 1644511149
transform 1 0 1748 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_11
timestamp 1644511149
transform 1 0 2116 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_23
timestamp 1644511149
transform 1 0 3220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_183
timestamp 1644511149
transform 1 0 17940 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1644511149
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_204
timestamp 1644511149
transform 1 0 19872 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_224
timestamp 1644511149
transform 1 0 21712 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_236
timestamp 1644511149
transform 1 0 22816 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_240
timestamp 1644511149
transform 1 0 23184 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_246
timestamp 1644511149
transform 1 0 23736 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_258
timestamp 1644511149
transform 1 0 24840 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_262
timestamp 1644511149
transform 1 0 25208 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_279
timestamp 1644511149
transform 1 0 26772 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_289
timestamp 1644511149
transform 1 0 27692 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_298
timestamp 1644511149
transform 1 0 28520 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_306
timestamp 1644511149
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_315
timestamp 1644511149
transform 1 0 30084 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_324
timestamp 1644511149
transform 1 0 30912 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_332
timestamp 1644511149
transform 1 0 31648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_340
timestamp 1644511149
transform 1 0 32384 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_360
timestamp 1644511149
transform 1 0 34224 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_379
timestamp 1644511149
transform 1 0 35972 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_388
timestamp 1644511149
transform 1 0 36800 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_400
timestamp 1644511149
transform 1 0 37904 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_412
timestamp 1644511149
transform 1 0 39008 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_421
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_433
timestamp 1644511149
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_445
timestamp 1644511149
transform 1 0 42044 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_469
timestamp 1644511149
transform 1 0 44252 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1644511149
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_188
timestamp 1644511149
transform 1 0 18400 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_202
timestamp 1644511149
transform 1 0 19688 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_213
timestamp 1644511149
transform 1 0 20700 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_221
timestamp 1644511149
transform 1 0 21436 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_237
timestamp 1644511149
transform 1 0 22908 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_245
timestamp 1644511149
transform 1 0 23644 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_256
timestamp 1644511149
transform 1 0 24656 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_263
timestamp 1644511149
transform 1 0 25300 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_270
timestamp 1644511149
transform 1 0 25944 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_278
timestamp 1644511149
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_313
timestamp 1644511149
transform 1 0 29900 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_321
timestamp 1644511149
transform 1 0 30636 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_332
timestamp 1644511149
transform 1 0 31648 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_353
timestamp 1644511149
transform 1 0 33580 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_370
timestamp 1644511149
transform 1 0 35144 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_382
timestamp 1644511149
transform 1 0 36248 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_390
timestamp 1644511149
transform 1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_397
timestamp 1644511149
transform 1 0 37628 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_417
timestamp 1644511149
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_429
timestamp 1644511149
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1644511149
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1644511149
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_449
timestamp 1644511149
transform 1 0 42412 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_457
timestamp 1644511149
transform 1 0 43148 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_462
timestamp 1644511149
transform 1 0 43608 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_469
timestamp 1644511149
transform 1 0 44252 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_14
timestamp 1644511149
transform 1 0 2392 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1644511149
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_165
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_177
timestamp 1644511149
transform 1 0 17388 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1644511149
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1644511149
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_203
timestamp 1644511149
transform 1 0 19780 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_214
timestamp 1644511149
transform 1 0 20792 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_238
timestamp 1644511149
transform 1 0 23000 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_244
timestamp 1644511149
transform 1 0 23552 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_248
timestamp 1644511149
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_260
timestamp 1644511149
transform 1 0 25024 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_280
timestamp 1644511149
transform 1 0 26864 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1644511149
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_326
timestamp 1644511149
transform 1 0 31096 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_332
timestamp 1644511149
transform 1 0 31648 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_342
timestamp 1644511149
transform 1 0 32568 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_351
timestamp 1644511149
transform 1 0 33396 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_358
timestamp 1644511149
transform 1 0 34040 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_374
timestamp 1644511149
transform 1 0 35512 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_387
timestamp 1644511149
transform 1 0 36708 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_393
timestamp 1644511149
transform 1 0 37260 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_403
timestamp 1644511149
transform 1 0 38180 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_410
timestamp 1644511149
transform 1 0 38824 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_418
timestamp 1644511149
transform 1 0 39560 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_421
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_433
timestamp 1644511149
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_445
timestamp 1644511149
transform 1 0 42044 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_469
timestamp 1644511149
transform 1 0 44252 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1644511149
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1644511149
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1644511149
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_87
timestamp 1644511149
transform 1 0 9108 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_91
timestamp 1644511149
transform 1 0 9476 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_103
timestamp 1644511149
transform 1 0 10580 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1644511149
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_181
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_192
timestamp 1644511149
transform 1 0 18768 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_205
timestamp 1644511149
transform 1 0 19964 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_213
timestamp 1644511149
transform 1 0 20700 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_220
timestamp 1644511149
transform 1 0 21344 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_231
timestamp 1644511149
transform 1 0 22356 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_238
timestamp 1644511149
transform 1 0 23000 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_244
timestamp 1644511149
transform 1 0 23552 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_249
timestamp 1644511149
transform 1 0 24012 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_269
timestamp 1644511149
transform 1 0 25852 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_277
timestamp 1644511149
transform 1 0 26588 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_286
timestamp 1644511149
transform 1 0 27416 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_295
timestamp 1644511149
transform 1 0 28244 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_302
timestamp 1644511149
transform 1 0 28888 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_310
timestamp 1644511149
transform 1 0 29624 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_320
timestamp 1644511149
transform 1 0 30544 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_328
timestamp 1644511149
transform 1 0 31280 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_353
timestamp 1644511149
transform 1 0 33580 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_365
timestamp 1644511149
transform 1 0 34684 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_381
timestamp 1644511149
transform 1 0 36156 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_389
timestamp 1644511149
transform 1 0 36892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_397
timestamp 1644511149
transform 1 0 37628 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_408
timestamp 1644511149
transform 1 0 38640 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_415
timestamp 1644511149
transform 1 0 39284 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_444
timestamp 1644511149
transform 1 0 41952 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_449
timestamp 1644511149
transform 1 0 42412 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_456
timestamp 1644511149
transform 1 0 43056 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_463
timestamp 1644511149
transform 1 0 43700 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_471
timestamp 1644511149
transform 1 0 44436 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_10
timestamp 1644511149
transform 1 0 2024 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_22
timestamp 1644511149
transform 1 0 3128 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_165
timestamp 1644511149
transform 1 0 16284 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_172
timestamp 1644511149
transform 1 0 16928 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_180
timestamp 1644511149
transform 1 0 17664 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_190
timestamp 1644511149
transform 1 0 18584 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_201
timestamp 1644511149
transform 1 0 19596 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_212
timestamp 1644511149
transform 1 0 20608 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_216
timestamp 1644511149
transform 1 0 20976 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_221
timestamp 1644511149
transform 1 0 21436 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_229
timestamp 1644511149
transform 1 0 22172 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1644511149
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1644511149
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_269
timestamp 1644511149
transform 1 0 25852 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_281
timestamp 1644511149
transform 1 0 26956 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_293
timestamp 1644511149
transform 1 0 28060 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_305
timestamp 1644511149
transform 1 0 29164 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_321
timestamp 1644511149
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_333
timestamp 1644511149
transform 1 0 31740 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_344
timestamp 1644511149
transform 1 0 32752 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_356
timestamp 1644511149
transform 1 0 33856 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_381
timestamp 1644511149
transform 1 0 36156 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_389
timestamp 1644511149
transform 1 0 36892 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_403
timestamp 1644511149
transform 1 0 38180 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_412
timestamp 1644511149
transform 1 0 39008 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_421
timestamp 1644511149
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_433
timestamp 1644511149
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_445
timestamp 1644511149
transform 1 0 42044 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_469
timestamp 1644511149
transform 1 0 44252 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_9
timestamp 1644511149
transform 1 0 1932 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_31
timestamp 1644511149
transform 1 0 3956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_43
timestamp 1644511149
transform 1 0 5060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_141
timestamp 1644511149
transform 1 0 14076 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_153
timestamp 1644511149
transform 1 0 15180 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_165
timestamp 1644511149
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_185
timestamp 1644511149
transform 1 0 18124 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_199
timestamp 1644511149
transform 1 0 19412 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_210
timestamp 1644511149
transform 1 0 20424 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_220
timestamp 1644511149
transform 1 0 21344 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_245
timestamp 1644511149
transform 1 0 23644 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_257
timestamp 1644511149
transform 1 0 24748 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_269
timestamp 1644511149
transform 1 0 25852 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_275
timestamp 1644511149
transform 1 0 26404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1644511149
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_291
timestamp 1644511149
transform 1 0 27876 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_311
timestamp 1644511149
transform 1 0 29716 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_331
timestamp 1644511149
transform 1 0 31556 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1644511149
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_341
timestamp 1644511149
transform 1 0 32476 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_353
timestamp 1644511149
transform 1 0 33580 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_366
timestamp 1644511149
transform 1 0 34776 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_374
timestamp 1644511149
transform 1 0 35512 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_386
timestamp 1644511149
transform 1 0 36616 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_398
timestamp 1644511149
transform 1 0 37720 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_406
timestamp 1644511149
transform 1 0 38456 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_414
timestamp 1644511149
transform 1 0 39192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_421
timestamp 1644511149
transform 1 0 39836 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_433
timestamp 1644511149
transform 1 0 40940 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_445
timestamp 1644511149
transform 1 0 42044 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_449
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_456
timestamp 1644511149
transform 1 0 43056 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_463
timestamp 1644511149
transform 1 0 43700 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_471
timestamp 1644511149
transform 1 0 44436 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_14
timestamp 1644511149
transform 1 0 2392 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_18
timestamp 1644511149
transform 1 0 2760 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_22
timestamp 1644511149
transform 1 0 3128 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_162
timestamp 1644511149
transform 1 0 16008 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_174
timestamp 1644511149
transform 1 0 17112 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_188
timestamp 1644511149
transform 1 0 18400 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_217
timestamp 1644511149
transform 1 0 21068 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_228
timestamp 1644511149
transform 1 0 22080 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_237
timestamp 1644511149
transform 1 0 22908 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_246
timestamp 1644511149
transform 1 0 23736 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_265
timestamp 1644511149
transform 1 0 25484 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_273
timestamp 1644511149
transform 1 0 26220 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_287
timestamp 1644511149
transform 1 0 27508 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_299
timestamp 1644511149
transform 1 0 28612 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_317
timestamp 1644511149
transform 1 0 30268 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_325
timestamp 1644511149
transform 1 0 31004 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_333
timestamp 1644511149
transform 1 0 31740 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_339
timestamp 1644511149
transform 1 0 32292 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_353
timestamp 1644511149
transform 1 0 33580 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_360
timestamp 1644511149
transform 1 0 34224 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_390
timestamp 1644511149
transform 1 0 36984 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_402
timestamp 1644511149
transform 1 0 38088 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_409
timestamp 1644511149
transform 1 0 38732 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_417
timestamp 1644511149
transform 1 0 39468 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_421
timestamp 1644511149
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_433
timestamp 1644511149
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_445
timestamp 1644511149
transform 1 0 42044 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_469
timestamp 1644511149
transform 1 0 44252 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1644511149
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1644511149
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1644511149
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1644511149
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_136
timestamp 1644511149
transform 1 0 13616 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_148
timestamp 1644511149
transform 1 0 14720 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_160
timestamp 1644511149
transform 1 0 15824 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_177
timestamp 1644511149
transform 1 0 17388 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_183
timestamp 1644511149
transform 1 0 17940 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_192
timestamp 1644511149
transform 1 0 18768 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_196
timestamp 1644511149
transform 1 0 19136 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_203
timestamp 1644511149
transform 1 0 19780 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_211
timestamp 1644511149
transform 1 0 20516 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1644511149
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1644511149
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_235
timestamp 1644511149
transform 1 0 22724 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_243
timestamp 1644511149
transform 1 0 23460 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_251
timestamp 1644511149
transform 1 0 24196 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_267
timestamp 1644511149
transform 1 0 25668 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_276
timestamp 1644511149
transform 1 0 26496 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_288
timestamp 1644511149
transform 1 0 27600 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_292
timestamp 1644511149
transform 1 0 27968 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_296
timestamp 1644511149
transform 1 0 28336 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_316
timestamp 1644511149
transform 1 0 30176 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_327
timestamp 1644511149
transform 1 0 31188 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1644511149
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_344
timestamp 1644511149
transform 1 0 32752 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_376
timestamp 1644511149
transform 1 0 35696 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_388
timestamp 1644511149
transform 1 0 36800 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_406
timestamp 1644511149
transform 1 0 38456 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_418
timestamp 1644511149
transform 1 0 39560 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_430
timestamp 1644511149
transform 1 0 40664 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_442
timestamp 1644511149
transform 1 0 41768 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_449
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_457
timestamp 1644511149
transform 1 0 43148 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_462
timestamp 1644511149
transform 1 0 43608 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_470
timestamp 1644511149
transform 1 0 44344 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_14
timestamp 1644511149
transform 1 0 2392 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1644511149
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_121
timestamp 1644511149
transform 1 0 12236 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_129
timestamp 1644511149
transform 1 0 12972 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1644511149
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_153
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_170
timestamp 1644511149
transform 1 0 16744 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_177
timestamp 1644511149
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1644511149
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1644511149
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_205
timestamp 1644511149
transform 1 0 19964 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_212
timestamp 1644511149
transform 1 0 20608 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_216
timestamp 1644511149
transform 1 0 20976 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_223
timestamp 1644511149
transform 1 0 21620 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_234
timestamp 1644511149
transform 1 0 22632 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_242
timestamp 1644511149
transform 1 0 23368 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1644511149
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_269
timestamp 1644511149
transform 1 0 25852 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_275
timestamp 1644511149
transform 1 0 26404 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_292
timestamp 1644511149
transform 1 0 27968 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_304
timestamp 1644511149
transform 1 0 29072 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_313
timestamp 1644511149
transform 1 0 29900 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_321
timestamp 1644511149
transform 1 0 30636 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_340
timestamp 1644511149
transform 1 0 32384 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_349
timestamp 1644511149
transform 1 0 33212 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_356
timestamp 1644511149
transform 1 0 33856 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_384
timestamp 1644511149
transform 1 0 36432 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_393
timestamp 1644511149
transform 1 0 37260 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_407
timestamp 1644511149
transform 1 0 38548 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_414
timestamp 1644511149
transform 1 0 39192 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_421
timestamp 1644511149
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_433
timestamp 1644511149
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_445
timestamp 1644511149
transform 1 0 42044 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_469
timestamp 1644511149
transform 1 0 44252 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1644511149
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1644511149
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1644511149
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_149
timestamp 1644511149
transform 1 0 14812 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_164
timestamp 1644511149
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_177
timestamp 1644511149
transform 1 0 17388 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_186
timestamp 1644511149
transform 1 0 18216 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_202
timestamp 1644511149
transform 1 0 19688 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_206
timestamp 1644511149
transform 1 0 20056 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_213
timestamp 1644511149
transform 1 0 20700 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_221
timestamp 1644511149
transform 1 0 21436 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_231
timestamp 1644511149
transform 1 0 22356 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_244
timestamp 1644511149
transform 1 0 23552 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_264
timestamp 1644511149
transform 1 0 25392 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_276
timestamp 1644511149
transform 1 0 26496 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_284
timestamp 1644511149
transform 1 0 27232 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_291
timestamp 1644511149
transform 1 0 27876 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_297
timestamp 1644511149
transform 1 0 28428 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_314
timestamp 1644511149
transform 1 0 29992 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_326
timestamp 1644511149
transform 1 0 31096 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_334
timestamp 1644511149
transform 1 0 31832 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_350
timestamp 1644511149
transform 1 0 33304 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_357
timestamp 1644511149
transform 1 0 33948 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_369
timestamp 1644511149
transform 1 0 35052 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_381
timestamp 1644511149
transform 1 0 36156 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_388
timestamp 1644511149
transform 1 0 36800 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_403
timestamp 1644511149
transform 1 0 38180 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_415
timestamp 1644511149
transform 1 0 39284 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_427
timestamp 1644511149
transform 1 0 40388 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_439
timestamp 1644511149
transform 1 0 41492 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1644511149
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_449
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_455
timestamp 1644511149
transform 1 0 42964 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_462
timestamp 1644511149
transform 1 0 43608 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_469
timestamp 1644511149
transform 1 0 44252 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_8
timestamp 1644511149
transform 1 0 1840 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1644511149
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_121
timestamp 1644511149
transform 1 0 12236 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_129
timestamp 1644511149
transform 1 0 12972 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_135
timestamp 1644511149
transform 1 0 13524 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1644511149
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_160
timestamp 1644511149
transform 1 0 15824 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_172
timestamp 1644511149
transform 1 0 16928 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1644511149
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_207
timestamp 1644511149
transform 1 0 20148 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_217
timestamp 1644511149
transform 1 0 21068 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_225
timestamp 1644511149
transform 1 0 21804 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_233
timestamp 1644511149
transform 1 0 22540 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_242
timestamp 1644511149
transform 1 0 23368 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1644511149
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_259
timestamp 1644511149
transform 1 0 24932 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_271
timestamp 1644511149
transform 1 0 26036 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_283
timestamp 1644511149
transform 1 0 27140 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_295
timestamp 1644511149
transform 1 0 28244 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1644511149
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_321
timestamp 1644511149
transform 1 0 30636 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_341
timestamp 1644511149
transform 1 0 32476 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_349
timestamp 1644511149
transform 1 0 33212 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_359
timestamp 1644511149
transform 1 0 34132 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_378
timestamp 1644511149
transform 1 0 35880 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_386
timestamp 1644511149
transform 1 0 36616 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_393
timestamp 1644511149
transform 1 0 37260 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_407
timestamp 1644511149
transform 1 0 38548 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1644511149
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_421
timestamp 1644511149
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_433
timestamp 1644511149
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_445
timestamp 1644511149
transform 1 0 42044 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_469
timestamp 1644511149
transform 1 0 44252 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_28
timestamp 1644511149
transform 1 0 3680 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_40
timestamp 1644511149
transform 1 0 4784 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_52
timestamp 1644511149
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_125
timestamp 1644511149
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_137
timestamp 1644511149
transform 1 0 13708 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_145
timestamp 1644511149
transform 1 0 14444 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_150
timestamp 1644511149
transform 1 0 14904 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_162
timestamp 1644511149
transform 1 0 16008 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_176
timestamp 1644511149
transform 1 0 17296 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_186
timestamp 1644511149
transform 1 0 18216 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_204
timestamp 1644511149
transform 1 0 19872 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_213
timestamp 1644511149
transform 1 0 20700 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_221
timestamp 1644511149
transform 1 0 21436 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_228
timestamp 1644511149
transform 1 0 22080 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_240
timestamp 1644511149
transform 1 0 23184 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_259
timestamp 1644511149
transform 1 0 24932 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_267
timestamp 1644511149
transform 1 0 25668 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_274
timestamp 1644511149
transform 1 0 26312 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_288
timestamp 1644511149
transform 1 0 27600 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_296
timestamp 1644511149
transform 1 0 28336 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_314
timestamp 1644511149
transform 1 0 29992 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_322
timestamp 1644511149
transform 1 0 30728 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1644511149
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_348
timestamp 1644511149
transform 1 0 33120 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_360
timestamp 1644511149
transform 1 0 34224 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_372
timestamp 1644511149
transform 1 0 35328 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_376
timestamp 1644511149
transform 1 0 35696 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_383
timestamp 1644511149
transform 1 0 36340 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1644511149
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_398
timestamp 1644511149
transform 1 0 37720 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_410
timestamp 1644511149
transform 1 0 38824 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_422
timestamp 1644511149
transform 1 0 39928 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_434
timestamp 1644511149
transform 1 0 41032 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_446
timestamp 1644511149
transform 1 0 42136 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_449
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_457
timestamp 1644511149
transform 1 0 43148 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_462
timestamp 1644511149
transform 1 0 43608 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_469
timestamp 1644511149
transform 1 0 44252 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_7
timestamp 1644511149
transform 1 0 1748 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_11
timestamp 1644511149
transform 1 0 2116 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_17
timestamp 1644511149
transform 1 0 2668 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_21
timestamp 1644511149
transform 1 0 3036 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_121
timestamp 1644511149
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1644511149
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_157
timestamp 1644511149
transform 1 0 15548 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_171
timestamp 1644511149
transform 1 0 16836 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_184
timestamp 1644511149
transform 1 0 18032 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_203
timestamp 1644511149
transform 1 0 19780 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_211
timestamp 1644511149
transform 1 0 20516 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_230
timestamp 1644511149
transform 1 0 22264 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_242
timestamp 1644511149
transform 1 0 23368 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1644511149
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_265
timestamp 1644511149
transform 1 0 25484 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_275
timestamp 1644511149
transform 1 0 26404 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_285
timestamp 1644511149
transform 1 0 27324 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_294
timestamp 1644511149
transform 1 0 28152 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1644511149
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1644511149
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_325
timestamp 1644511149
transform 1 0 31004 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_333
timestamp 1644511149
transform 1 0 31740 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_339
timestamp 1644511149
transform 1 0 32292 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_343
timestamp 1644511149
transform 1 0 32660 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_350
timestamp 1644511149
transform 1 0 33304 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_362
timestamp 1644511149
transform 1 0 34408 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_372
timestamp 1644511149
transform 1 0 35328 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_382
timestamp 1644511149
transform 1 0 36248 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_395
timestamp 1644511149
transform 1 0 37444 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_407
timestamp 1644511149
transform 1 0 38548 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1644511149
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_421
timestamp 1644511149
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_433
timestamp 1644511149
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_445
timestamp 1644511149
transform 1 0 42044 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_469
timestamp 1644511149
transform 1 0 44252 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_9
timestamp 1644511149
transform 1 0 1932 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_31
timestamp 1644511149
transform 1 0 3956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_43
timestamp 1644511149
transform 1 0 5060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_125
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_137
timestamp 1644511149
transform 1 0 13708 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_141
timestamp 1644511149
transform 1 0 14076 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_150
timestamp 1644511149
transform 1 0 14904 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_164
timestamp 1644511149
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_174
timestamp 1644511149
transform 1 0 17112 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_178
timestamp 1644511149
transform 1 0 17480 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_185
timestamp 1644511149
transform 1 0 18124 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_194
timestamp 1644511149
transform 1 0 18952 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_202
timestamp 1644511149
transform 1 0 19688 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_211
timestamp 1644511149
transform 1 0 20516 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1644511149
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_231
timestamp 1644511149
transform 1 0 22356 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_237
timestamp 1644511149
transform 1 0 22908 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_254
timestamp 1644511149
transform 1 0 24472 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_274
timestamp 1644511149
transform 1 0 26312 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_288
timestamp 1644511149
transform 1 0 27600 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_312
timestamp 1644511149
transform 1 0 29808 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_320
timestamp 1644511149
transform 1 0 30544 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_332
timestamp 1644511149
transform 1 0 31648 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_351
timestamp 1644511149
transform 1 0 33396 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_371
timestamp 1644511149
transform 1 0 35236 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_384
timestamp 1644511149
transform 1 0 36432 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_29_396
timestamp 1644511149
transform 1 0 37536 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_402
timestamp 1644511149
transform 1 0 38088 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_424
timestamp 1644511149
transform 1 0 40112 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_436
timestamp 1644511149
transform 1 0 41216 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_449
timestamp 1644511149
transform 1 0 42412 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_457
timestamp 1644511149
transform 1 0 43148 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_462
timestamp 1644511149
transform 1 0 43608 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_470
timestamp 1644511149
transform 1 0 44344 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_9
timestamp 1644511149
transform 1 0 1932 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_13
timestamp 1644511149
transform 1 0 2300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_25
timestamp 1644511149
transform 1 0 3404 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_117
timestamp 1644511149
transform 1 0 11868 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_128
timestamp 1644511149
transform 1 0 12880 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_157
timestamp 1644511149
transform 1 0 15548 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_164
timestamp 1644511149
transform 1 0 16192 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_172
timestamp 1644511149
transform 1 0 16928 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_180
timestamp 1644511149
transform 1 0 17664 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_191
timestamp 1644511149
transform 1 0 18676 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1644511149
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_209
timestamp 1644511149
transform 1 0 20332 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_227
timestamp 1644511149
transform 1 0 21988 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_235
timestamp 1644511149
transform 1 0 22724 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_241
timestamp 1644511149
transform 1 0 23276 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_249
timestamp 1644511149
transform 1 0 24012 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_265
timestamp 1644511149
transform 1 0 25484 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_273
timestamp 1644511149
transform 1 0 26220 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_277
timestamp 1644511149
transform 1 0 26588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_291
timestamp 1644511149
transform 1 0 27876 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_299
timestamp 1644511149
transform 1 0 28612 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1644511149
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_317
timestamp 1644511149
transform 1 0 30268 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_325
timestamp 1644511149
transform 1 0 31004 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_343
timestamp 1644511149
transform 1 0 32660 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_355
timestamp 1644511149
transform 1 0 33764 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1644511149
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_372
timestamp 1644511149
transform 1 0 35328 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_384
timestamp 1644511149
transform 1 0 36432 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_391
timestamp 1644511149
transform 1 0 37076 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_398
timestamp 1644511149
transform 1 0 37720 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_407
timestamp 1644511149
transform 1 0 38548 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1644511149
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_421
timestamp 1644511149
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_433
timestamp 1644511149
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_445
timestamp 1644511149
transform 1 0 42044 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_469
timestamp 1644511149
transform 1 0 44252 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1644511149
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1644511149
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1644511149
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1644511149
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1644511149
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1644511149
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_128
timestamp 1644511149
transform 1 0 12880 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_138
timestamp 1644511149
transform 1 0 13800 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_150
timestamp 1644511149
transform 1 0 14904 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_159
timestamp 1644511149
transform 1 0 15732 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1644511149
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_181
timestamp 1644511149
transform 1 0 17756 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_187
timestamp 1644511149
transform 1 0 18308 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_192
timestamp 1644511149
transform 1 0 18768 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_205
timestamp 1644511149
transform 1 0 19964 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_215
timestamp 1644511149
transform 1 0 20884 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1644511149
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_232
timestamp 1644511149
transform 1 0 22448 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_240
timestamp 1644511149
transform 1 0 23184 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_260
timestamp 1644511149
transform 1 0 25024 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_272
timestamp 1644511149
transform 1 0 26128 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_286
timestamp 1644511149
transform 1 0 27416 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_298
timestamp 1644511149
transform 1 0 28520 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_310
timestamp 1644511149
transform 1 0 29624 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_332
timestamp 1644511149
transform 1 0 31648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_337
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_349
timestamp 1644511149
transform 1 0 33212 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_366
timestamp 1644511149
transform 1 0 34776 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_378
timestamp 1644511149
transform 1 0 35880 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_390
timestamp 1644511149
transform 1 0 36984 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_405
timestamp 1644511149
transform 1 0 38364 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_412
timestamp 1644511149
transform 1 0 39008 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_424
timestamp 1644511149
transform 1 0 40112 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_436
timestamp 1644511149
transform 1 0 41216 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_440
timestamp 1644511149
transform 1 0 41584 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_449
timestamp 1644511149
transform 1 0 42412 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_453
timestamp 1644511149
transform 1 0 42780 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_457
timestamp 1644511149
transform 1 0 43148 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_461
timestamp 1644511149
transform 1 0 43516 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_465
timestamp 1644511149
transform 1 0 43884 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_12
timestamp 1644511149
transform 1 0 2208 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_24
timestamp 1644511149
transform 1 0 3312 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_109
timestamp 1644511149
transform 1 0 11132 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_117
timestamp 1644511149
transform 1 0 11868 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_131
timestamp 1644511149
transform 1 0 13156 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1644511149
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_149
timestamp 1644511149
transform 1 0 14812 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_156
timestamp 1644511149
transform 1 0 15456 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_170
timestamp 1644511149
transform 1 0 16744 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_180
timestamp 1644511149
transform 1 0 17664 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_184
timestamp 1644511149
transform 1 0 18032 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_190
timestamp 1644511149
transform 1 0 18584 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_203
timestamp 1644511149
transform 1 0 19780 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_209
timestamp 1644511149
transform 1 0 20332 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_216
timestamp 1644511149
transform 1 0 20976 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_224
timestamp 1644511149
transform 1 0 21712 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_232
timestamp 1644511149
transform 1 0 22448 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_239
timestamp 1644511149
transform 1 0 23092 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1644511149
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_265
timestamp 1644511149
transform 1 0 25484 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_287
timestamp 1644511149
transform 1 0 27508 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_299
timestamp 1644511149
transform 1 0 28612 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1644511149
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_321
timestamp 1644511149
transform 1 0 30636 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_328
timestamp 1644511149
transform 1 0 31280 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_347
timestamp 1644511149
transform 1 0 33028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_359
timestamp 1644511149
transform 1 0 34132 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1644511149
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_389
timestamp 1644511149
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_401
timestamp 1644511149
transform 1 0 37996 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_409
timestamp 1644511149
transform 1 0 38732 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_416
timestamp 1644511149
transform 1 0 39376 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_421
timestamp 1644511149
transform 1 0 39836 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_434
timestamp 1644511149
transform 1 0 41032 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_442
timestamp 1644511149
transform 1 0 41768 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_464
timestamp 1644511149
transform 1 0 43792 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_472
timestamp 1644511149
transform 1 0 44528 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_93
timestamp 1644511149
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1644511149
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1644511149
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_130
timestamp 1644511149
transform 1 0 13064 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_138
timestamp 1644511149
transform 1 0 13800 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_156
timestamp 1644511149
transform 1 0 15456 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_164
timestamp 1644511149
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_180
timestamp 1644511149
transform 1 0 17664 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_184
timestamp 1644511149
transform 1 0 18032 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_190
timestamp 1644511149
transform 1 0 18584 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_33_203
timestamp 1644511149
transform 1 0 19780 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_209
timestamp 1644511149
transform 1 0 20332 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_220
timestamp 1644511149
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_231
timestamp 1644511149
transform 1 0 22356 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_237
timestamp 1644511149
transform 1 0 22908 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_244
timestamp 1644511149
transform 1 0 23552 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_256
timestamp 1644511149
transform 1 0 24656 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_276
timestamp 1644511149
transform 1 0 26496 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_293
timestamp 1644511149
transform 1 0 28060 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_311
timestamp 1644511149
transform 1 0 29716 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_317
timestamp 1644511149
transform 1 0 30268 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_321
timestamp 1644511149
transform 1 0 30636 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_332
timestamp 1644511149
transform 1 0 31648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_340
timestamp 1644511149
transform 1 0 32384 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_352
timestamp 1644511149
transform 1 0 33488 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_372
timestamp 1644511149
transform 1 0 35328 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_384
timestamp 1644511149
transform 1 0 36432 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_415
timestamp 1644511149
transform 1 0 39284 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_435
timestamp 1644511149
transform 1 0 41124 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1644511149
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_449
timestamp 1644511149
transform 1 0 42412 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_458
timestamp 1644511149
transform 1 0 43240 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_465
timestamp 1644511149
transform 1 0 43884 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_10
timestamp 1644511149
transform 1 0 2024 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_22
timestamp 1644511149
transform 1 0 3128 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_45
timestamp 1644511149
transform 1 0 5244 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_50
timestamp 1644511149
transform 1 0 5704 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_66
timestamp 1644511149
transform 1 0 7176 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_78
timestamp 1644511149
transform 1 0 8280 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_109
timestamp 1644511149
transform 1 0 11132 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_115
timestamp 1644511149
transform 1 0 11684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_127
timestamp 1644511149
transform 1 0 12788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1644511149
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_145
timestamp 1644511149
transform 1 0 14444 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_149
timestamp 1644511149
transform 1 0 14812 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_161
timestamp 1644511149
transform 1 0 15916 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_174
timestamp 1644511149
transform 1 0 17112 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_188
timestamp 1644511149
transform 1 0 18400 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_217
timestamp 1644511149
transform 1 0 21068 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_237
timestamp 1644511149
transform 1 0 22908 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_247
timestamp 1644511149
transform 1 0 23828 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1644511149
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_256
timestamp 1644511149
transform 1 0 24656 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_268
timestamp 1644511149
transform 1 0 25760 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_274
timestamp 1644511149
transform 1 0 26312 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_285
timestamp 1644511149
transform 1 0 27324 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_293
timestamp 1644511149
transform 1 0 28060 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_300
timestamp 1644511149
transform 1 0 28704 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_318
timestamp 1644511149
transform 1 0 30360 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_330
timestamp 1644511149
transform 1 0 31464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_337
timestamp 1644511149
transform 1 0 32108 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_349
timestamp 1644511149
transform 1 0 33212 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_359
timestamp 1644511149
transform 1 0 34132 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1644511149
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_371
timestamp 1644511149
transform 1 0 35236 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_379
timestamp 1644511149
transform 1 0 35972 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_391
timestamp 1644511149
transform 1 0 37076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_403
timestamp 1644511149
transform 1 0 38180 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_412
timestamp 1644511149
transform 1 0 39008 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_34_421
timestamp 1644511149
transform 1 0 39836 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_432
timestamp 1644511149
transform 1 0 40848 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_444
timestamp 1644511149
transform 1 0 41952 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_469
timestamp 1644511149
transform 1 0 44252 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_52
timestamp 1644511149
transform 1 0 5888 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_93
timestamp 1644511149
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1644511149
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1644511149
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_137
timestamp 1644511149
transform 1 0 13708 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_145
timestamp 1644511149
transform 1 0 14444 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_164
timestamp 1644511149
transform 1 0 16192 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_181
timestamp 1644511149
transform 1 0 17756 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_190
timestamp 1644511149
transform 1 0 18584 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_198
timestamp 1644511149
transform 1 0 19320 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_206
timestamp 1644511149
transform 1 0 20056 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_212
timestamp 1644511149
transform 1 0 20608 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_218
timestamp 1644511149
transform 1 0 21160 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_228
timestamp 1644511149
transform 1 0 22080 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_248
timestamp 1644511149
transform 1 0 23920 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_268
timestamp 1644511149
transform 1 0 25760 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_290
timestamp 1644511149
transform 1 0 27784 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_303
timestamp 1644511149
transform 1 0 28980 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_311
timestamp 1644511149
transform 1 0 29716 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_319
timestamp 1644511149
transform 1 0 30452 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_326
timestamp 1644511149
transform 1 0 31096 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_334
timestamp 1644511149
transform 1 0 31832 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_337
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_349
timestamp 1644511149
transform 1 0 33212 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_353
timestamp 1644511149
transform 1 0 33580 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_370
timestamp 1644511149
transform 1 0 35144 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_378
timestamp 1644511149
transform 1 0 35880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_388
timestamp 1644511149
transform 1 0 36800 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_401
timestamp 1644511149
transform 1 0 37996 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_415
timestamp 1644511149
transform 1 0 39284 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_421
timestamp 1644511149
transform 1 0 39836 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_425
timestamp 1644511149
transform 1 0 40204 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_437
timestamp 1644511149
transform 1 0 41308 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_445
timestamp 1644511149
transform 1 0 42044 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_452
timestamp 1644511149
transform 1 0 42688 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_460
timestamp 1644511149
transform 1 0 43424 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_465
timestamp 1644511149
transform 1 0 43884 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_9
timestamp 1644511149
transform 1 0 1932 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_13
timestamp 1644511149
transform 1 0 2300 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_17
timestamp 1644511149
transform 1 0 2668 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_21
timestamp 1644511149
transform 1 0 3036 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_66
timestamp 1644511149
transform 1 0 7176 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_78
timestamp 1644511149
transform 1 0 8280 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_109
timestamp 1644511149
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_121
timestamp 1644511149
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1644511149
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1644511149
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_153
timestamp 1644511149
transform 1 0 15180 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_36_163
timestamp 1644511149
transform 1 0 16100 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_175
timestamp 1644511149
transform 1 0 17204 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_188
timestamp 1644511149
transform 1 0 18400 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_36_200
timestamp 1644511149
transform 1 0 19504 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_36_209
timestamp 1644511149
transform 1 0 20332 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_218
timestamp 1644511149
transform 1 0 21160 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_238
timestamp 1644511149
transform 1 0 23000 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1644511149
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_265
timestamp 1644511149
transform 1 0 25484 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_273
timestamp 1644511149
transform 1 0 26220 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_284
timestamp 1644511149
transform 1 0 27232 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_298
timestamp 1644511149
transform 1 0 28520 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_306
timestamp 1644511149
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_313
timestamp 1644511149
transform 1 0 29900 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_320
timestamp 1644511149
transform 1 0 30544 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_337
timestamp 1644511149
transform 1 0 32108 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_345
timestamp 1644511149
transform 1 0 32844 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_353
timestamp 1644511149
transform 1 0 33580 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_360
timestamp 1644511149
transform 1 0 34224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_368
timestamp 1644511149
transform 1 0 34960 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_374
timestamp 1644511149
transform 1 0 35512 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_382
timestamp 1644511149
transform 1 0 36248 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_394
timestamp 1644511149
transform 1 0 37352 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_403
timestamp 1644511149
transform 1 0 38180 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_409
timestamp 1644511149
transform 1 0 38732 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_416
timestamp 1644511149
transform 1 0 39376 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_421
timestamp 1644511149
transform 1 0 39836 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_443
timestamp 1644511149
transform 1 0 41860 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_447
timestamp 1644511149
transform 1 0 42228 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_469
timestamp 1644511149
transform 1 0 44252 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_30
timestamp 1644511149
transform 1 0 3864 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_42
timestamp 1644511149
transform 1 0 4968 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1644511149
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_63
timestamp 1644511149
transform 1 0 6900 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_75
timestamp 1644511149
transform 1 0 8004 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_87
timestamp 1644511149
transform 1 0 9108 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_99
timestamp 1644511149
transform 1 0 10212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_125
timestamp 1644511149
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_137
timestamp 1644511149
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_149
timestamp 1644511149
transform 1 0 14812 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_155
timestamp 1644511149
transform 1 0 15364 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_164
timestamp 1644511149
transform 1 0 16192 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_175
timestamp 1644511149
transform 1 0 17204 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_184
timestamp 1644511149
transform 1 0 18032 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_190
timestamp 1644511149
transform 1 0 18584 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_207
timestamp 1644511149
transform 1 0 20148 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_218
timestamp 1644511149
transform 1 0 21160 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_235
timestamp 1644511149
transform 1 0 22724 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_245
timestamp 1644511149
transform 1 0 23644 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_257
timestamp 1644511149
transform 1 0 24748 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1644511149
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1644511149
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_297
timestamp 1644511149
transform 1 0 28428 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_308
timestamp 1644511149
transform 1 0 29440 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_315
timestamp 1644511149
transform 1 0 30084 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_319
timestamp 1644511149
transform 1 0 30452 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_327
timestamp 1644511149
transform 1 0 31188 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1644511149
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_337
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_343
timestamp 1644511149
transform 1 0 32660 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_347
timestamp 1644511149
transform 1 0 33028 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_355
timestamp 1644511149
transform 1 0 33764 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_365
timestamp 1644511149
transform 1 0 34684 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_373
timestamp 1644511149
transform 1 0 35420 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_381
timestamp 1644511149
transform 1 0 36156 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_388
timestamp 1644511149
transform 1 0 36800 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_407
timestamp 1644511149
transform 1 0 38548 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_417
timestamp 1644511149
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_429
timestamp 1644511149
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1644511149
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1644511149
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_454
timestamp 1644511149
transform 1 0 42872 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_458
timestamp 1644511149
transform 1 0 43240 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_462
timestamp 1644511149
transform 1 0 43608 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_470
timestamp 1644511149
transform 1 0 44344 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_24
timestamp 1644511149
transform 1 0 3312 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_121
timestamp 1644511149
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1644511149
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1644511149
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_153
timestamp 1644511149
transform 1 0 15180 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_171
timestamp 1644511149
transform 1 0 16836 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_187
timestamp 1644511149
transform 1 0 18308 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1644511149
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_205
timestamp 1644511149
transform 1 0 19964 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_213
timestamp 1644511149
transform 1 0 20700 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_232
timestamp 1644511149
transform 1 0 22448 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_240
timestamp 1644511149
transform 1 0 23184 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_247
timestamp 1644511149
transform 1 0 23828 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1644511149
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_257
timestamp 1644511149
transform 1 0 24748 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_275
timestamp 1644511149
transform 1 0 26404 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_279
timestamp 1644511149
transform 1 0 26772 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_283
timestamp 1644511149
transform 1 0 27140 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_297
timestamp 1644511149
transform 1 0 28428 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_305
timestamp 1644511149
transform 1 0 29164 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_313
timestamp 1644511149
transform 1 0 29900 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_319
timestamp 1644511149
transform 1 0 30452 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_328
timestamp 1644511149
transform 1 0 31280 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_340
timestamp 1644511149
transform 1 0 32384 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_352
timestamp 1644511149
transform 1 0 33488 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1644511149
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1644511149
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_377
timestamp 1644511149
transform 1 0 35788 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_386
timestamp 1644511149
transform 1 0 36616 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_397
timestamp 1644511149
transform 1 0 37628 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_405
timestamp 1644511149
transform 1 0 38364 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_416
timestamp 1644511149
transform 1 0 39376 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_421
timestamp 1644511149
transform 1 0 39836 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_438
timestamp 1644511149
transform 1 0 41400 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_446
timestamp 1644511149
transform 1 0 42136 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_469
timestamp 1644511149
transform 1 0 44252 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_12
timestamp 1644511149
transform 1 0 2208 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_19
timestamp 1644511149
transform 1 0 2852 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_31
timestamp 1644511149
transform 1 0 3956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_43
timestamp 1644511149
transform 1 0 5060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_125
timestamp 1644511149
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_137
timestamp 1644511149
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_149
timestamp 1644511149
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_164
timestamp 1644511149
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_177
timestamp 1644511149
transform 1 0 17388 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_191
timestamp 1644511149
transform 1 0 18676 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_199
timestamp 1644511149
transform 1 0 19412 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_210
timestamp 1644511149
transform 1 0 20424 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1644511149
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1644511149
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_233
timestamp 1644511149
transform 1 0 22540 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_261
timestamp 1644511149
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1644511149
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1644511149
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_287
timestamp 1644511149
transform 1 0 27508 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_293
timestamp 1644511149
transform 1 0 28060 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_301
timestamp 1644511149
transform 1 0 28796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_309
timestamp 1644511149
transform 1 0 29532 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_317
timestamp 1644511149
transform 1 0 30268 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_321
timestamp 1644511149
transform 1 0 30636 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_332
timestamp 1644511149
transform 1 0 31648 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_340
timestamp 1644511149
transform 1 0 32384 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_348
timestamp 1644511149
transform 1 0 33120 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_354
timestamp 1644511149
transform 1 0 33672 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_374
timestamp 1644511149
transform 1 0 35512 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_388
timestamp 1644511149
transform 1 0 36800 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_398
timestamp 1644511149
transform 1 0 37720 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_412
timestamp 1644511149
transform 1 0 39008 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_424
timestamp 1644511149
transform 1 0 40112 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_435
timestamp 1644511149
transform 1 0 41124 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_444
timestamp 1644511149
transform 1 0 41952 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_452
timestamp 1644511149
transform 1 0 42688 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_459
timestamp 1644511149
transform 1 0 43332 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_466
timestamp 1644511149
transform 1 0 43976 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_472
timestamp 1644511149
transform 1 0 44528 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_109
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_121
timestamp 1644511149
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1644511149
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1644511149
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_153
timestamp 1644511149
transform 1 0 15180 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_173
timestamp 1644511149
transform 1 0 17020 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_181
timestamp 1644511149
transform 1 0 17756 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_190
timestamp 1644511149
transform 1 0 18584 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_205
timestamp 1644511149
transform 1 0 19964 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_217
timestamp 1644511149
transform 1 0 21068 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_229
timestamp 1644511149
transform 1 0 22172 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_241
timestamp 1644511149
transform 1 0 23276 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_247
timestamp 1644511149
transform 1 0 23828 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1644511149
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_263
timestamp 1644511149
transform 1 0 25300 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_274
timestamp 1644511149
transform 1 0 26312 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_282
timestamp 1644511149
transform 1 0 27048 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_292
timestamp 1644511149
transform 1 0 27968 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_296
timestamp 1644511149
transform 1 0 28336 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_302
timestamp 1644511149
transform 1 0 28888 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_40_309
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_319
timestamp 1644511149
transform 1 0 30452 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_330
timestamp 1644511149
transform 1 0 31464 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_339
timestamp 1644511149
transform 1 0 32292 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_351
timestamp 1644511149
transform 1 0 33396 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1644511149
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_377
timestamp 1644511149
transform 1 0 35788 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_395
timestamp 1644511149
transform 1 0 37444 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_404
timestamp 1644511149
transform 1 0 38272 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_416
timestamp 1644511149
transform 1 0 39376 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_421
timestamp 1644511149
transform 1 0 39836 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_429
timestamp 1644511149
transform 1 0 40572 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_435
timestamp 1644511149
transform 1 0 41124 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_444
timestamp 1644511149
transform 1 0 41952 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_469
timestamp 1644511149
transform 1 0 44252 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_93
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1644511149
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_125
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_137
timestamp 1644511149
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_149
timestamp 1644511149
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1644511149
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1644511149
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_181
timestamp 1644511149
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_193
timestamp 1644511149
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_205
timestamp 1644511149
transform 1 0 19964 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_210
timestamp 1644511149
transform 1 0 20424 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1644511149
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_233
timestamp 1644511149
transform 1 0 22540 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_243
timestamp 1644511149
transform 1 0 23460 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_255
timestamp 1644511149
transform 1 0 24564 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_259
timestamp 1644511149
transform 1 0 24932 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_270
timestamp 1644511149
transform 1 0 25944 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_278
timestamp 1644511149
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_305
timestamp 1644511149
transform 1 0 29164 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_319
timestamp 1644511149
transform 1 0 30452 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_332
timestamp 1644511149
transform 1 0 31648 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_341
timestamp 1644511149
transform 1 0 32476 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_348
timestamp 1644511149
transform 1 0 33120 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_360
timestamp 1644511149
transform 1 0 34224 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_372
timestamp 1644511149
transform 1 0 35328 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_384
timestamp 1644511149
transform 1 0 36432 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_401
timestamp 1644511149
transform 1 0 37996 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_420
timestamp 1644511149
transform 1 0 39744 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_440
timestamp 1644511149
transform 1 0 41584 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_41_452
timestamp 1644511149
transform 1 0 42688 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_461
timestamp 1644511149
transform 1 0 43516 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_468
timestamp 1644511149
transform 1 0 44160 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_472
timestamp 1644511149
transform 1 0 44528 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1644511149
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_32
timestamp 1644511149
transform 1 0 4048 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_44
timestamp 1644511149
transform 1 0 5152 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_56
timestamp 1644511149
transform 1 0 6256 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_68
timestamp 1644511149
transform 1 0 7360 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_80
timestamp 1644511149
transform 1 0 8464 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_97
timestamp 1644511149
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_109
timestamp 1644511149
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_121
timestamp 1644511149
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1644511149
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1644511149
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_153
timestamp 1644511149
transform 1 0 15180 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_173
timestamp 1644511149
transform 1 0 17020 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_181
timestamp 1644511149
transform 1 0 17756 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_188
timestamp 1644511149
transform 1 0 18400 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_210
timestamp 1644511149
transform 1 0 20424 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_221
timestamp 1644511149
transform 1 0 21436 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_227
timestamp 1644511149
transform 1 0 21988 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_231
timestamp 1644511149
transform 1 0 22356 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1644511149
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1644511149
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_263
timestamp 1644511149
transform 1 0 25300 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_277
timestamp 1644511149
transform 1 0 26588 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_289
timestamp 1644511149
transform 1 0 27692 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_304
timestamp 1644511149
transform 1 0 29072 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_314
timestamp 1644511149
transform 1 0 29992 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_323
timestamp 1644511149
transform 1 0 30820 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_334
timestamp 1644511149
transform 1 0 31832 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_342
timestamp 1644511149
transform 1 0 32568 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_360
timestamp 1644511149
transform 1 0 34224 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_377
timestamp 1644511149
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_389
timestamp 1644511149
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_401
timestamp 1644511149
transform 1 0 37996 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_409
timestamp 1644511149
transform 1 0 38732 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_416
timestamp 1644511149
transform 1 0 39376 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_421
timestamp 1644511149
transform 1 0 39836 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_444
timestamp 1644511149
transform 1 0 41952 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_469
timestamp 1644511149
transform 1 0 44252 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_23
timestamp 1644511149
transform 1 0 3220 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_45
timestamp 1644511149
transform 1 0 5244 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_53
timestamp 1644511149
transform 1 0 5980 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_125
timestamp 1644511149
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_137
timestamp 1644511149
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_149
timestamp 1644511149
transform 1 0 14812 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_157
timestamp 1644511149
transform 1 0 15548 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 1644511149
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_174
timestamp 1644511149
transform 1 0 17112 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_198
timestamp 1644511149
transform 1 0 19320 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_218
timestamp 1644511149
transform 1 0 21160 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_242
timestamp 1644511149
transform 1 0 23368 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_256
timestamp 1644511149
transform 1 0 24656 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_276
timestamp 1644511149
transform 1 0 26496 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_285
timestamp 1644511149
transform 1 0 27324 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_297
timestamp 1644511149
transform 1 0 28428 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_306
timestamp 1644511149
transform 1 0 29256 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_318
timestamp 1644511149
transform 1 0 30360 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1644511149
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1644511149
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_342
timestamp 1644511149
transform 1 0 32568 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_356
timestamp 1644511149
transform 1 0 33856 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_366
timestamp 1644511149
transform 1 0 34776 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_373
timestamp 1644511149
transform 1 0 35420 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_380
timestamp 1644511149
transform 1 0 36064 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_410
timestamp 1644511149
transform 1 0 38824 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_418
timestamp 1644511149
transform 1 0 39560 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_430
timestamp 1644511149
transform 1 0 40664 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_442
timestamp 1644511149
transform 1 0 41768 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_452
timestamp 1644511149
transform 1 0 42688 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_460
timestamp 1644511149
transform 1 0 43424 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_465
timestamp 1644511149
transform 1 0 43884 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_121
timestamp 1644511149
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1644511149
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_153
timestamp 1644511149
transform 1 0 15180 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_158
timestamp 1644511149
transform 1 0 15640 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_166
timestamp 1644511149
transform 1 0 16376 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_171
timestamp 1644511149
transform 1 0 16836 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_180
timestamp 1644511149
transform 1 0 17664 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_188
timestamp 1644511149
transform 1 0 18400 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_44_207
timestamp 1644511149
transform 1 0 20148 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_213
timestamp 1644511149
transform 1 0 20700 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_221
timestamp 1644511149
transform 1 0 21436 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_233
timestamp 1644511149
transform 1 0 22540 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_248
timestamp 1644511149
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_261
timestamp 1644511149
transform 1 0 25116 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_270
timestamp 1644511149
transform 1 0 25944 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_277
timestamp 1644511149
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_289
timestamp 1644511149
transform 1 0 27692 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_297
timestamp 1644511149
transform 1 0 28428 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1644511149
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1644511149
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_321
timestamp 1644511149
transform 1 0 30636 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_329
timestamp 1644511149
transform 1 0 31372 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_340
timestamp 1644511149
transform 1 0 32384 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_349
timestamp 1644511149
transform 1 0 33212 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_359
timestamp 1644511149
transform 1 0 34132 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1644511149
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_372
timestamp 1644511149
transform 1 0 35328 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_376
timestamp 1644511149
transform 1 0 35696 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_393
timestamp 1644511149
transform 1 0 37260 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_405
timestamp 1644511149
transform 1 0 38364 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_417
timestamp 1644511149
transform 1 0 39468 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_421
timestamp 1644511149
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_433
timestamp 1644511149
transform 1 0 40940 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_439
timestamp 1644511149
transform 1 0 41492 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_461
timestamp 1644511149
transform 1 0 43516 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_468
timestamp 1644511149
transform 1 0 44160 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_472
timestamp 1644511149
transform 1 0 44528 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1644511149
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_137
timestamp 1644511149
transform 1 0 13708 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_145
timestamp 1644511149
transform 1 0 14444 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_164
timestamp 1644511149
transform 1 0 16192 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_173
timestamp 1644511149
transform 1 0 17020 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_182
timestamp 1644511149
transform 1 0 17848 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_189
timestamp 1644511149
transform 1 0 18492 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_201
timestamp 1644511149
transform 1 0 19596 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_213
timestamp 1644511149
transform 1 0 20700 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_221
timestamp 1644511149
transform 1 0 21436 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_241
timestamp 1644511149
transform 1 0 23276 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_253
timestamp 1644511149
transform 1 0 24380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_265
timestamp 1644511149
transform 1 0 25484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_277
timestamp 1644511149
transform 1 0 26588 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_293
timestamp 1644511149
transform 1 0 28060 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_304
timestamp 1644511149
transform 1 0 29072 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_316
timestamp 1644511149
transform 1 0 30176 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_328
timestamp 1644511149
transform 1 0 31280 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_349
timestamp 1644511149
transform 1 0 33212 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_356
timestamp 1644511149
transform 1 0 33856 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_368
timestamp 1644511149
transform 1 0 34960 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_388
timestamp 1644511149
transform 1 0 36800 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_405
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_417
timestamp 1644511149
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_429
timestamp 1644511149
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1644511149
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1644511149
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_449
timestamp 1644511149
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_461
timestamp 1644511149
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_121
timestamp 1644511149
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1644511149
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1644511149
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_153
timestamp 1644511149
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_171
timestamp 1644511149
transform 1 0 16836 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_180
timestamp 1644511149
transform 1 0 17664 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_188
timestamp 1644511149
transform 1 0 18400 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_209
timestamp 1644511149
transform 1 0 20332 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_219
timestamp 1644511149
transform 1 0 21252 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_226
timestamp 1644511149
transform 1 0 21896 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_237
timestamp 1644511149
transform 1 0 22908 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_244
timestamp 1644511149
transform 1 0 23552 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_259
timestamp 1644511149
transform 1 0 24932 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_263
timestamp 1644511149
transform 1 0 25300 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_283
timestamp 1644511149
transform 1 0 27140 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_287
timestamp 1644511149
transform 1 0 27508 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_304
timestamp 1644511149
transform 1 0 29072 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_319
timestamp 1644511149
transform 1 0 30452 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_327
timestamp 1644511149
transform 1 0 31188 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_337
timestamp 1644511149
transform 1 0 32108 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_344
timestamp 1644511149
transform 1 0 32752 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_356
timestamp 1644511149
transform 1 0 33856 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_368
timestamp 1644511149
transform 1 0 34960 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_383
timestamp 1644511149
transform 1 0 36340 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_395
timestamp 1644511149
transform 1 0 37444 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_407
timestamp 1644511149
transform 1 0 38548 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1644511149
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_421
timestamp 1644511149
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_433
timestamp 1644511149
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_445
timestamp 1644511149
transform 1 0 42044 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_469
timestamp 1644511149
transform 1 0 44252 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1644511149
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_137
timestamp 1644511149
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_154
timestamp 1644511149
transform 1 0 15272 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_160
timestamp 1644511149
transform 1 0 15824 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_164
timestamp 1644511149
transform 1 0 16192 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_173
timestamp 1644511149
transform 1 0 17020 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_180
timestamp 1644511149
transform 1 0 17664 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_194
timestamp 1644511149
transform 1 0 18952 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_201
timestamp 1644511149
transform 1 0 19596 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_213
timestamp 1644511149
transform 1 0 20700 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_220
timestamp 1644511149
transform 1 0 21344 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_235
timestamp 1644511149
transform 1 0 22724 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_255
timestamp 1644511149
transform 1 0 24564 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_264
timestamp 1644511149
transform 1 0 25392 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_276
timestamp 1644511149
transform 1 0 26496 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_292
timestamp 1644511149
transform 1 0 27968 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_301
timestamp 1644511149
transform 1 0 28796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_310
timestamp 1644511149
transform 1 0 29624 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_321
timestamp 1644511149
transform 1 0 30636 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_332
timestamp 1644511149
transform 1 0 31648 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_356
timestamp 1644511149
transform 1 0 33856 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_365
timestamp 1644511149
transform 1 0 34684 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_377
timestamp 1644511149
transform 1 0 35788 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_388
timestamp 1644511149
transform 1 0 36800 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_396
timestamp 1644511149
transform 1 0 37536 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_408
timestamp 1644511149
transform 1 0 38640 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_420
timestamp 1644511149
transform 1 0 39744 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_432
timestamp 1644511149
transform 1 0 40848 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_444
timestamp 1644511149
transform 1 0 41952 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_449
timestamp 1644511149
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_461
timestamp 1644511149
transform 1 0 43516 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_465
timestamp 1644511149
transform 1 0 43884 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_109
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_121
timestamp 1644511149
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1644511149
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1644511149
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_159
timestamp 1644511149
transform 1 0 15732 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_171
timestamp 1644511149
transform 1 0 16836 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_184
timestamp 1644511149
transform 1 0 18032 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_192
timestamp 1644511149
transform 1 0 18768 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_203
timestamp 1644511149
transform 1 0 19780 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_220
timestamp 1644511149
transform 1 0 21344 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_231
timestamp 1644511149
transform 1 0 22356 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_235
timestamp 1644511149
transform 1 0 22724 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_244
timestamp 1644511149
transform 1 0 23552 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_263
timestamp 1644511149
transform 1 0 25300 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_273
timestamp 1644511149
transform 1 0 26220 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_285
timestamp 1644511149
transform 1 0 27324 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_294
timestamp 1644511149
transform 1 0 28152 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1644511149
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1644511149
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_313
timestamp 1644511149
transform 1 0 29900 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_320
timestamp 1644511149
transform 1 0 30544 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_332
timestamp 1644511149
transform 1 0 31648 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_341
timestamp 1644511149
transform 1 0 32476 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_349
timestamp 1644511149
transform 1 0 33212 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_360
timestamp 1644511149
transform 1 0 34224 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_370
timestamp 1644511149
transform 1 0 35144 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_379
timestamp 1644511149
transform 1 0 35972 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_383
timestamp 1644511149
transform 1 0 36340 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_400
timestamp 1644511149
transform 1 0 37904 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_412
timestamp 1644511149
transform 1 0 39008 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_421
timestamp 1644511149
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_433
timestamp 1644511149
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_445
timestamp 1644511149
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_457
timestamp 1644511149
transform 1 0 43148 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_463
timestamp 1644511149
transform 1 0 43700 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_471
timestamp 1644511149
transform 1 0 44436 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1644511149
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_133
timestamp 1644511149
transform 1 0 13340 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_152
timestamp 1644511149
transform 1 0 15088 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_164
timestamp 1644511149
transform 1 0 16192 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_177
timestamp 1644511149
transform 1 0 17388 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_181
timestamp 1644511149
transform 1 0 17756 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_189
timestamp 1644511149
transform 1 0 18492 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_196
timestamp 1644511149
transform 1 0 19136 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_204
timestamp 1644511149
transform 1 0 19872 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_209
timestamp 1644511149
transform 1 0 20332 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_221
timestamp 1644511149
transform 1 0 21436 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_241
timestamp 1644511149
transform 1 0 23276 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_249
timestamp 1644511149
transform 1 0 24012 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_258
timestamp 1644511149
transform 1 0 24840 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_267
timestamp 1644511149
transform 1 0 25668 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1644511149
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_293
timestamp 1644511149
transform 1 0 28060 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_49_302
timestamp 1644511149
transform 1 0 28888 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_311
timestamp 1644511149
transform 1 0 29716 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_321
timestamp 1644511149
transform 1 0 30636 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_332
timestamp 1644511149
transform 1 0 31648 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_342
timestamp 1644511149
transform 1 0 32568 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_350
timestamp 1644511149
transform 1 0 33304 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_360
timestamp 1644511149
transform 1 0 34224 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_372
timestamp 1644511149
transform 1 0 35328 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_380
timestamp 1644511149
transform 1 0 36064 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_387
timestamp 1644511149
transform 1 0 36708 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1644511149
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_405
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_417
timestamp 1644511149
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_429
timestamp 1644511149
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1644511149
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1644511149
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_449
timestamp 1644511149
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_461
timestamp 1644511149
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_14
timestamp 1644511149
transform 1 0 2392 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_26
timestamp 1644511149
transform 1 0 3496 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_146
timestamp 1644511149
transform 1 0 14536 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_158
timestamp 1644511149
transform 1 0 15640 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_162
timestamp 1644511149
transform 1 0 16008 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_171
timestamp 1644511149
transform 1 0 16836 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_50_186
timestamp 1644511149
transform 1 0 18216 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_194
timestamp 1644511149
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_204
timestamp 1644511149
transform 1 0 19872 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_214
timestamp 1644511149
transform 1 0 20792 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_226
timestamp 1644511149
transform 1 0 21896 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_238
timestamp 1644511149
transform 1 0 23000 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_250
timestamp 1644511149
transform 1 0 24104 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_265
timestamp 1644511149
transform 1 0 25484 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_283
timestamp 1644511149
transform 1 0 27140 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_296
timestamp 1644511149
transform 1 0 28336 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_303
timestamp 1644511149
transform 1 0 28980 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1644511149
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_317
timestamp 1644511149
transform 1 0 30268 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_323
timestamp 1644511149
transform 1 0 30820 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_337
timestamp 1644511149
transform 1 0 32108 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_341
timestamp 1644511149
transform 1 0 32476 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_346
timestamp 1644511149
transform 1 0 32936 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_360
timestamp 1644511149
transform 1 0 34224 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_370
timestamp 1644511149
transform 1 0 35144 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_390
timestamp 1644511149
transform 1 0 36984 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_402
timestamp 1644511149
transform 1 0 38088 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_414
timestamp 1644511149
transform 1 0 39192 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_421
timestamp 1644511149
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_433
timestamp 1644511149
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_445
timestamp 1644511149
transform 1 0 42044 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_469
timestamp 1644511149
transform 1 0 44252 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_28
timestamp 1644511149
transform 1 0 3680 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_40
timestamp 1644511149
transform 1 0 4784 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_52
timestamp 1644511149
transform 1 0 5888 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_149
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1644511149
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1644511149
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_177
timestamp 1644511149
transform 1 0 17388 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_181
timestamp 1644511149
transform 1 0 17756 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_190
timestamp 1644511149
transform 1 0 18584 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_202
timestamp 1644511149
transform 1 0 19688 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_214
timestamp 1644511149
transform 1 0 20792 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1644511149
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_233
timestamp 1644511149
transform 1 0 22540 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_245
timestamp 1644511149
transform 1 0 23644 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_249
timestamp 1644511149
transform 1 0 24012 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_257
timestamp 1644511149
transform 1 0 24748 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_265
timestamp 1644511149
transform 1 0 25484 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_269
timestamp 1644511149
transform 1 0 25852 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_275
timestamp 1644511149
transform 1 0 26404 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1644511149
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_284
timestamp 1644511149
transform 1 0 27232 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_51_306
timestamp 1644511149
transform 1 0 29256 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_320
timestamp 1644511149
transform 1 0 30544 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_332
timestamp 1644511149
transform 1 0 31648 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_340
timestamp 1644511149
transform 1 0 32384 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_360
timestamp 1644511149
transform 1 0 34224 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_374
timestamp 1644511149
transform 1 0 35512 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_51_384
timestamp 1644511149
transform 1 0 36432 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_396
timestamp 1644511149
transform 1 0 37536 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_408
timestamp 1644511149
transform 1 0 38640 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_420
timestamp 1644511149
transform 1 0 39744 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_432
timestamp 1644511149
transform 1 0 40848 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_444
timestamp 1644511149
transform 1 0 41952 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_449
timestamp 1644511149
transform 1 0 42412 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_457
timestamp 1644511149
transform 1 0 43148 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_462
timestamp 1644511149
transform 1 0 43608 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_469
timestamp 1644511149
transform 1 0 44252 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_10
timestamp 1644511149
transform 1 0 2024 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_22
timestamp 1644511149
transform 1 0 3128 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_153
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_164
timestamp 1644511149
transform 1 0 16192 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_171
timestamp 1644511149
transform 1 0 16836 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_179
timestamp 1644511149
transform 1 0 17572 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_187
timestamp 1644511149
transform 1 0 18308 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1644511149
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_200
timestamp 1644511149
transform 1 0 19504 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_216
timestamp 1644511149
transform 1 0 20976 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_228
timestamp 1644511149
transform 1 0 22080 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_234
timestamp 1644511149
transform 1 0 22632 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_242
timestamp 1644511149
transform 1 0 23368 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_248
timestamp 1644511149
transform 1 0 23920 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_260
timestamp 1644511149
transform 1 0 25024 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_270
timestamp 1644511149
transform 1 0 25944 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_278
timestamp 1644511149
transform 1 0 26680 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_289
timestamp 1644511149
transform 1 0 27692 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_298
timestamp 1644511149
transform 1 0 28520 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_306
timestamp 1644511149
transform 1 0 29256 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_327
timestamp 1644511149
transform 1 0 31188 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_339
timestamp 1644511149
transform 1 0 32292 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_343
timestamp 1644511149
transform 1 0 32660 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_360
timestamp 1644511149
transform 1 0 34224 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_377
timestamp 1644511149
transform 1 0 35788 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_395
timestamp 1644511149
transform 1 0 37444 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_407
timestamp 1644511149
transform 1 0 38548 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1644511149
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_421
timestamp 1644511149
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_433
timestamp 1644511149
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_445
timestamp 1644511149
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_457
timestamp 1644511149
transform 1 0 43148 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_469
timestamp 1644511149
transform 1 0 44252 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1644511149
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1644511149
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_39
timestamp 1644511149
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1644511149
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1644511149
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_155
timestamp 1644511149
transform 1 0 15364 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_159
timestamp 1644511149
transform 1 0 15732 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_164
timestamp 1644511149
transform 1 0 16192 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_179
timestamp 1644511149
transform 1 0 17572 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_187
timestamp 1644511149
transform 1 0 18308 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_198
timestamp 1644511149
transform 1 0 19320 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_220
timestamp 1644511149
transform 1 0 21344 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_243
timestamp 1644511149
transform 1 0 23460 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_251
timestamp 1644511149
transform 1 0 24196 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_258
timestamp 1644511149
transform 1 0 24840 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_268
timestamp 1644511149
transform 1 0 25760 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_275
timestamp 1644511149
transform 1 0 26404 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1644511149
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_287
timestamp 1644511149
transform 1 0 27508 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_296
timestamp 1644511149
transform 1 0 28336 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_308
timestamp 1644511149
transform 1 0 29440 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_312
timestamp 1644511149
transform 1 0 29808 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_323
timestamp 1644511149
transform 1 0 30820 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_332
timestamp 1644511149
transform 1 0 31648 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_340
timestamp 1644511149
transform 1 0 32384 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_352
timestamp 1644511149
transform 1 0 33488 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_364
timestamp 1644511149
transform 1 0 34592 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_372
timestamp 1644511149
transform 1 0 35328 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_384
timestamp 1644511149
transform 1 0 36432 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_405
timestamp 1644511149
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_417
timestamp 1644511149
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_429
timestamp 1644511149
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1644511149
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1644511149
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_449
timestamp 1644511149
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_461
timestamp 1644511149
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1644511149
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1644511149
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_157
timestamp 1644511149
transform 1 0 15548 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_168
timestamp 1644511149
transform 1 0 16560 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_172
timestamp 1644511149
transform 1 0 16928 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_183
timestamp 1644511149
transform 1 0 17940 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_192
timestamp 1644511149
transform 1 0 18768 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_213
timestamp 1644511149
transform 1 0 20700 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_217
timestamp 1644511149
transform 1 0 21068 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_222
timestamp 1644511149
transform 1 0 21528 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_228
timestamp 1644511149
transform 1 0 22080 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_235
timestamp 1644511149
transform 1 0 22724 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_244
timestamp 1644511149
transform 1 0 23552 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_258
timestamp 1644511149
transform 1 0 24840 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_266
timestamp 1644511149
transform 1 0 25576 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_272
timestamp 1644511149
transform 1 0 26128 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_300
timestamp 1644511149
transform 1 0 28704 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_313
timestamp 1644511149
transform 1 0 29900 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_333
timestamp 1644511149
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_345
timestamp 1644511149
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1644511149
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1644511149
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_382
timestamp 1644511149
transform 1 0 36248 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_389
timestamp 1644511149
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_401
timestamp 1644511149
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1644511149
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1644511149
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_421
timestamp 1644511149
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_433
timestamp 1644511149
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_445
timestamp 1644511149
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_457
timestamp 1644511149
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_469
timestamp 1644511149
transform 1 0 44252 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1644511149
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1644511149
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_39
timestamp 1644511149
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1644511149
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1644511149
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_164
timestamp 1644511149
transform 1 0 16192 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_174
timestamp 1644511149
transform 1 0 17112 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_190
timestamp 1644511149
transform 1 0 18584 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_202
timestamp 1644511149
transform 1 0 19688 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_214
timestamp 1644511149
transform 1 0 20792 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_220
timestamp 1644511149
transform 1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_237
timestamp 1644511149
transform 1 0 22908 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_247
timestamp 1644511149
transform 1 0 23828 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_255
timestamp 1644511149
transform 1 0 24564 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_267
timestamp 1644511149
transform 1 0 25668 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_276
timestamp 1644511149
transform 1 0 26496 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_287
timestamp 1644511149
transform 1 0 27508 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_294
timestamp 1644511149
transform 1 0 28152 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_298
timestamp 1644511149
transform 1 0 28520 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_315
timestamp 1644511149
transform 1 0 30084 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_323
timestamp 1644511149
transform 1 0 30820 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1644511149
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_349
timestamp 1644511149
transform 1 0 33212 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_367
timestamp 1644511149
transform 1 0 34868 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_375
timestamp 1644511149
transform 1 0 35604 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_382
timestamp 1644511149
transform 1 0 36248 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_390
timestamp 1644511149
transform 1 0 36984 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_396
timestamp 1644511149
transform 1 0 37536 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_408
timestamp 1644511149
transform 1 0 38640 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_426
timestamp 1644511149
transform 1 0 40296 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_438
timestamp 1644511149
transform 1 0 41400 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_446
timestamp 1644511149
transform 1 0 42136 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_449
timestamp 1644511149
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_461
timestamp 1644511149
transform 1 0 43516 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_465
timestamp 1644511149
transform 1 0 43884 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1644511149
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_160
timestamp 1644511149
transform 1 0 15824 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_172
timestamp 1644511149
transform 1 0 16928 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_180
timestamp 1644511149
transform 1 0 17664 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_187
timestamp 1644511149
transform 1 0 18308 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1644511149
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_200
timestamp 1644511149
transform 1 0 19504 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_212
timestamp 1644511149
transform 1 0 20608 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_224
timestamp 1644511149
transform 1 0 21712 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_248
timestamp 1644511149
transform 1 0 23920 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_56_272
timestamp 1644511149
transform 1 0 26128 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_278
timestamp 1644511149
transform 1 0 26680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_285
timestamp 1644511149
transform 1 0 27324 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_297
timestamp 1644511149
transform 1 0 28428 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_305
timestamp 1644511149
transform 1 0 29164 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_321
timestamp 1644511149
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_333
timestamp 1644511149
transform 1 0 31740 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_339
timestamp 1644511149
transform 1 0 32292 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_346
timestamp 1644511149
transform 1 0 32936 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_354
timestamp 1644511149
transform 1 0 33672 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_360
timestamp 1644511149
transform 1 0 34224 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_380
timestamp 1644511149
transform 1 0 36064 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_389
timestamp 1644511149
transform 1 0 36892 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_409
timestamp 1644511149
transform 1 0 38732 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_416
timestamp 1644511149
transform 1 0 39376 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_421
timestamp 1644511149
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_433
timestamp 1644511149
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_445
timestamp 1644511149
transform 1 0 42044 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_469
timestamp 1644511149
transform 1 0 44252 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1644511149
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1644511149
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1644511149
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1644511149
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_149
timestamp 1644511149
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_164
timestamp 1644511149
transform 1 0 16192 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_182
timestamp 1644511149
transform 1 0 17848 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_193
timestamp 1644511149
transform 1 0 18860 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_213
timestamp 1644511149
transform 1 0 20700 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_220
timestamp 1644511149
transform 1 0 21344 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_231
timestamp 1644511149
transform 1 0 22356 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_239
timestamp 1644511149
transform 1 0 23092 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_246
timestamp 1644511149
transform 1 0 23736 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_57_258
timestamp 1644511149
transform 1 0 24840 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_266
timestamp 1644511149
transform 1 0 25576 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_272
timestamp 1644511149
transform 1 0 26128 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_284
timestamp 1644511149
transform 1 0 27232 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_288
timestamp 1644511149
transform 1 0 27600 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_296
timestamp 1644511149
transform 1 0 28336 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_304
timestamp 1644511149
transform 1 0 29072 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_311
timestamp 1644511149
transform 1 0 29716 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_323
timestamp 1644511149
transform 1 0 30820 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_332
timestamp 1644511149
transform 1 0 31648 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_353
timestamp 1644511149
transform 1 0 33580 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_361
timestamp 1644511149
transform 1 0 34316 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_365
timestamp 1644511149
transform 1 0 34684 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_376
timestamp 1644511149
transform 1 0 35696 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_387
timestamp 1644511149
transform 1 0 36708 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1644511149
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_399
timestamp 1644511149
transform 1 0 37812 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_408
timestamp 1644511149
transform 1 0 38640 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_416
timestamp 1644511149
transform 1 0 39376 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_423
timestamp 1644511149
transform 1 0 40020 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_435
timestamp 1644511149
transform 1 0 41124 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1644511149
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_449
timestamp 1644511149
transform 1 0 42412 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_456
timestamp 1644511149
transform 1 0 43056 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_463
timestamp 1644511149
transform 1 0 43700 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_471
timestamp 1644511149
transform 1 0 44436 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1644511149
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1644511149
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_171
timestamp 1644511149
transform 1 0 16836 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_177
timestamp 1644511149
transform 1 0 17388 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_188
timestamp 1644511149
transform 1 0 18400 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_211
timestamp 1644511149
transform 1 0 20516 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_225
timestamp 1644511149
transform 1 0 21804 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_232
timestamp 1644511149
transform 1 0 22448 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_239
timestamp 1644511149
transform 1 0 23092 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1644511149
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_257
timestamp 1644511149
transform 1 0 24748 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_263
timestamp 1644511149
transform 1 0 25300 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_272
timestamp 1644511149
transform 1 0 26128 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_284
timestamp 1644511149
transform 1 0 27232 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_291
timestamp 1644511149
transform 1 0 27876 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_298
timestamp 1644511149
transform 1 0 28520 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_306
timestamp 1644511149
transform 1 0 29256 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_312
timestamp 1644511149
transform 1 0 29808 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_336
timestamp 1644511149
transform 1 0 32016 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_345
timestamp 1644511149
transform 1 0 32844 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_351
timestamp 1644511149
transform 1 0 33396 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_359
timestamp 1644511149
transform 1 0 34132 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1644511149
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_368
timestamp 1644511149
transform 1 0 34960 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_376
timestamp 1644511149
transform 1 0 35696 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_387
timestamp 1644511149
transform 1 0 36708 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_395
timestamp 1644511149
transform 1 0 37444 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_403
timestamp 1644511149
transform 1 0 38180 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_412
timestamp 1644511149
transform 1 0 39008 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_421
timestamp 1644511149
transform 1 0 39836 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_438
timestamp 1644511149
transform 1 0 41400 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_446
timestamp 1644511149
transform 1 0 42136 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_469
timestamp 1644511149
transform 1 0 44252 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1644511149
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1644511149
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1644511149
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1644511149
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1644511149
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_164
timestamp 1644511149
transform 1 0 16192 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_185
timestamp 1644511149
transform 1 0 18124 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_194
timestamp 1644511149
transform 1 0 18952 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_59_205
timestamp 1644511149
transform 1 0 19964 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_213
timestamp 1644511149
transform 1 0 20700 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_220
timestamp 1644511149
transform 1 0 21344 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_232
timestamp 1644511149
transform 1 0 22448 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_243
timestamp 1644511149
transform 1 0 23460 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_250
timestamp 1644511149
transform 1 0 24104 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_59_272
timestamp 1644511149
transform 1 0 26128 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_295
timestamp 1644511149
transform 1 0 28244 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_306
timestamp 1644511149
transform 1 0 29256 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_313
timestamp 1644511149
transform 1 0 29900 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_317
timestamp 1644511149
transform 1 0 30268 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_323
timestamp 1644511149
transform 1 0 30820 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1644511149
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_348
timestamp 1644511149
transform 1 0 33120 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_360
timestamp 1644511149
transform 1 0 34224 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_372
timestamp 1644511149
transform 1 0 35328 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_384
timestamp 1644511149
transform 1 0 36432 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_404
timestamp 1644511149
transform 1 0 38272 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_414
timestamp 1644511149
transform 1 0 39192 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_420
timestamp 1644511149
transform 1 0 39744 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_427
timestamp 1644511149
transform 1 0 40388 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_435
timestamp 1644511149
transform 1 0 41124 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_440
timestamp 1644511149
transform 1 0 41584 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_449
timestamp 1644511149
transform 1 0 42412 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_453
timestamp 1644511149
transform 1 0 42780 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_457
timestamp 1644511149
transform 1 0 43148 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_464
timestamp 1644511149
transform 1 0 43792 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_472
timestamp 1644511149
transform 1 0 44528 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1644511149
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_165
timestamp 1644511149
transform 1 0 16284 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_173
timestamp 1644511149
transform 1 0 17020 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_180
timestamp 1644511149
transform 1 0 17664 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_192
timestamp 1644511149
transform 1 0 18768 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_60_206
timestamp 1644511149
transform 1 0 20056 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_218
timestamp 1644511149
transform 1 0 21160 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_226
timestamp 1644511149
transform 1 0 21896 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_231
timestamp 1644511149
transform 1 0 22356 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_240
timestamp 1644511149
transform 1 0 23184 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_248
timestamp 1644511149
transform 1 0 23920 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_260
timestamp 1644511149
transform 1 0 25024 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_281
timestamp 1644511149
transform 1 0 26956 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_294
timestamp 1644511149
transform 1 0 28152 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_303
timestamp 1644511149
transform 1 0 28980 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1644511149
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_325
timestamp 1644511149
transform 1 0 31004 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_337
timestamp 1644511149
transform 1 0 32108 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_343
timestamp 1644511149
transform 1 0 32660 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_353
timestamp 1644511149
transform 1 0 33580 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_360
timestamp 1644511149
transform 1 0 34224 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_373
timestamp 1644511149
transform 1 0 35420 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_381
timestamp 1644511149
transform 1 0 36156 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_393
timestamp 1644511149
transform 1 0 37260 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_405
timestamp 1644511149
transform 1 0 38364 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1644511149
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1644511149
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_421
timestamp 1644511149
transform 1 0 39836 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_427
timestamp 1644511149
transform 1 0 40388 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_444
timestamp 1644511149
transform 1 0 41952 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_469
timestamp 1644511149
transform 1 0 44252 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1644511149
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1644511149
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_39
timestamp 1644511149
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1644511149
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1644511149
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_181
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_61_196
timestamp 1644511149
transform 1 0 19136 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_204
timestamp 1644511149
transform 1 0 19872 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_214
timestamp 1644511149
transform 1 0 20792 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_222
timestamp 1644511149
transform 1 0 21528 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_231
timestamp 1644511149
transform 1 0 22356 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_251
timestamp 1644511149
transform 1 0 24196 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_263
timestamp 1644511149
transform 1 0 25300 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_275
timestamp 1644511149
transform 1 0 26404 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1644511149
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_284
timestamp 1644511149
transform 1 0 27232 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_293
timestamp 1644511149
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_305
timestamp 1644511149
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_317
timestamp 1644511149
transform 1 0 30268 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_325
timestamp 1644511149
transform 1 0 31004 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_332
timestamp 1644511149
transform 1 0 31648 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_345
timestamp 1644511149
transform 1 0 32844 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_357
timestamp 1644511149
transform 1 0 33948 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_367
timestamp 1644511149
transform 1 0 34868 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_374
timestamp 1644511149
transform 1 0 35512 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_382
timestamp 1644511149
transform 1 0 36248 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_388
timestamp 1644511149
transform 1 0 36800 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_397
timestamp 1644511149
transform 1 0 37628 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_411
timestamp 1644511149
transform 1 0 38916 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_422
timestamp 1644511149
transform 1 0 39928 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_432
timestamp 1644511149
transform 1 0 40848 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_438
timestamp 1644511149
transform 1 0 41400 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_444
timestamp 1644511149
transform 1 0 41952 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_449
timestamp 1644511149
transform 1 0 42412 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_457
timestamp 1644511149
transform 1 0 43148 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_461
timestamp 1644511149
transform 1 0 43516 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_468
timestamp 1644511149
transform 1 0 44160 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_472
timestamp 1644511149
transform 1 0 44528 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1644511149
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1644511149
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_177
timestamp 1644511149
transform 1 0 17388 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_184
timestamp 1644511149
transform 1 0 18032 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_192
timestamp 1644511149
transform 1 0 18768 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_197
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_62_210
timestamp 1644511149
transform 1 0 20424 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_224
timestamp 1644511149
transform 1 0 21712 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_236
timestamp 1644511149
transform 1 0 22816 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_242
timestamp 1644511149
transform 1 0 23368 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_246
timestamp 1644511149
transform 1 0 23736 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_62_253
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_268
timestamp 1644511149
transform 1 0 25760 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_275
timestamp 1644511149
transform 1 0 26404 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_291
timestamp 1644511149
transform 1 0 27876 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_298
timestamp 1644511149
transform 1 0 28520 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_306
timestamp 1644511149
transform 1 0 29256 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_309
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_321
timestamp 1644511149
transform 1 0 30636 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_330
timestamp 1644511149
transform 1 0 31464 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_342
timestamp 1644511149
transform 1 0 32568 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_346
timestamp 1644511149
transform 1 0 32936 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_351
timestamp 1644511149
transform 1 0 33396 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_360
timestamp 1644511149
transform 1 0 34224 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_382
timestamp 1644511149
transform 1 0 36248 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_402
timestamp 1644511149
transform 1 0 38088 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_406
timestamp 1644511149
transform 1 0 38456 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_416
timestamp 1644511149
transform 1 0 39376 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_426
timestamp 1644511149
transform 1 0 40296 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_435
timestamp 1644511149
transform 1 0 41124 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_442
timestamp 1644511149
transform 1 0 41768 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_469
timestamp 1644511149
transform 1 0 44252 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_15
timestamp 1644511149
transform 1 0 2484 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_19
timestamp 1644511149
transform 1 0 2852 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_31
timestamp 1644511149
transform 1 0 3956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_43
timestamp 1644511149
transform 1 0 5060 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1644511149
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_175
timestamp 1644511149
transform 1 0 17204 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_183
timestamp 1644511149
transform 1 0 17940 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_189
timestamp 1644511149
transform 1 0 18492 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_195
timestamp 1644511149
transform 1 0 19044 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_202
timestamp 1644511149
transform 1 0 19688 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1644511149
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1644511149
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_233
timestamp 1644511149
transform 1 0 22540 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_245
timestamp 1644511149
transform 1 0 23644 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_249
timestamp 1644511149
transform 1 0 24012 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_254
timestamp 1644511149
transform 1 0 24472 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_265
timestamp 1644511149
transform 1 0 25484 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_271
timestamp 1644511149
transform 1 0 26036 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_276
timestamp 1644511149
transform 1 0 26496 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_295
timestamp 1644511149
transform 1 0 28244 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_306
timestamp 1644511149
transform 1 0 29256 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_328
timestamp 1644511149
transform 1 0 31280 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_343
timestamp 1644511149
transform 1 0 32660 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_347
timestamp 1644511149
transform 1 0 33028 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_352
timestamp 1644511149
transform 1 0 33488 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_363
timestamp 1644511149
transform 1 0 34500 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_373
timestamp 1644511149
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1644511149
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1644511149
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_397
timestamp 1644511149
transform 1 0 37628 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_424
timestamp 1644511149
transform 1 0 40112 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_436
timestamp 1644511149
transform 1 0 41216 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_444
timestamp 1644511149
transform 1 0 41952 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_454
timestamp 1644511149
transform 1 0 42872 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_462
timestamp 1644511149
transform 1 0 43608 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_469
timestamp 1644511149
transform 1 0 44252 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_24
timestamp 1644511149
transform 1 0 3312 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_177
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_64_190
timestamp 1644511149
transform 1 0 18584 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_64_207
timestamp 1644511149
transform 1 0 20148 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_215
timestamp 1644511149
transform 1 0 20884 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_219
timestamp 1644511149
transform 1 0 21252 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_231
timestamp 1644511149
transform 1 0 22356 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_239
timestamp 1644511149
transform 1 0 23092 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_248
timestamp 1644511149
transform 1 0 23920 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_265
timestamp 1644511149
transform 1 0 25484 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_275
timestamp 1644511149
transform 1 0 26404 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_283
timestamp 1644511149
transform 1 0 27140 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_292
timestamp 1644511149
transform 1 0 27968 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_303
timestamp 1644511149
transform 1 0 28980 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1644511149
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_337
timestamp 1644511149
transform 1 0 32108 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_348
timestamp 1644511149
transform 1 0 33120 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1644511149
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1644511149
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_369
timestamp 1644511149
transform 1 0 35052 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_381
timestamp 1644511149
transform 1 0 36156 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_389
timestamp 1644511149
transform 1 0 36892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_394
timestamp 1644511149
transform 1 0 37352 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_406
timestamp 1644511149
transform 1 0 38456 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_412
timestamp 1644511149
transform 1 0 39008 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_416
timestamp 1644511149
transform 1 0 39376 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_421
timestamp 1644511149
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_433
timestamp 1644511149
transform 1 0 40940 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_444
timestamp 1644511149
transform 1 0 41952 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_448
timestamp 1644511149
transform 1 0 42320 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_465
timestamp 1644511149
transform 1 0 43884 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_65_3
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_65_12
timestamp 1644511149
transform 1 0 2208 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_24
timestamp 1644511149
transform 1 0 3312 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_36
timestamp 1644511149
transform 1 0 4416 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_48
timestamp 1644511149
transform 1 0 5520 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_93
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1644511149
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_125
timestamp 1644511149
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_137
timestamp 1644511149
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_149
timestamp 1644511149
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1644511149
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1644511149
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_169
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_177
timestamp 1644511149
transform 1 0 17388 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_185
timestamp 1644511149
transform 1 0 18124 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_194
timestamp 1644511149
transform 1 0 18952 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_203
timestamp 1644511149
transform 1 0 19780 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_212
timestamp 1644511149
transform 1 0 20608 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_220
timestamp 1644511149
transform 1 0 21344 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_225
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_253
timestamp 1644511149
transform 1 0 24380 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_261
timestamp 1644511149
transform 1 0 25116 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_265
timestamp 1644511149
transform 1 0 25484 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_276
timestamp 1644511149
transform 1 0 26496 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_281
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_289
timestamp 1644511149
transform 1 0 27692 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_296
timestamp 1644511149
transform 1 0 28336 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_308
timestamp 1644511149
transform 1 0 29440 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_320
timestamp 1644511149
transform 1 0 30544 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_331
timestamp 1644511149
transform 1 0 31556 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1644511149
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_343
timestamp 1644511149
transform 1 0 32660 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_356
timestamp 1644511149
transform 1 0 33856 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_376
timestamp 1644511149
transform 1 0 35696 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_388
timestamp 1644511149
transform 1 0 36800 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_398
timestamp 1644511149
transform 1 0 37720 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_422
timestamp 1644511149
transform 1 0 39928 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_437
timestamp 1644511149
transform 1 0 41308 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_444
timestamp 1644511149
transform 1 0 41952 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_453
timestamp 1644511149
transform 1 0 42780 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_65_464
timestamp 1644511149
transform 1 0 43792 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_472
timestamp 1644511149
transform 1 0 44528 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1644511149
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1644511149
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1644511149
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_97
timestamp 1644511149
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_109
timestamp 1644511149
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_121
timestamp 1644511149
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1644511149
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1644511149
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_153
timestamp 1644511149
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_181
timestamp 1644511149
transform 1 0 17756 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_193
timestamp 1644511149
transform 1 0 18860 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_66_197
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_204
timestamp 1644511149
transform 1 0 19872 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_224
timestamp 1644511149
transform 1 0 21712 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_231
timestamp 1644511149
transform 1 0 22356 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_235
timestamp 1644511149
transform 1 0 22724 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_240
timestamp 1644511149
transform 1 0 23184 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_253
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_261
timestamp 1644511149
transform 1 0 25116 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_66_270
timestamp 1644511149
transform 1 0 25944 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_66_279
timestamp 1644511149
transform 1 0 26772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_291
timestamp 1644511149
transform 1 0 27876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_303
timestamp 1644511149
transform 1 0 28980 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1644511149
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_309
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_316
timestamp 1644511149
transform 1 0 30176 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_328
timestamp 1644511149
transform 1 0 31280 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_340
timestamp 1644511149
transform 1 0 32384 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_348
timestamp 1644511149
transform 1 0 33120 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_360
timestamp 1644511149
transform 1 0 34224 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_369
timestamp 1644511149
transform 1 0 35052 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_377
timestamp 1644511149
transform 1 0 35788 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_66_396
timestamp 1644511149
transform 1 0 37536 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_402
timestamp 1644511149
transform 1 0 38088 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_411
timestamp 1644511149
transform 1 0 38916 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1644511149
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_424
timestamp 1644511149
transform 1 0 40112 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_444
timestamp 1644511149
transform 1 0 41952 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_469
timestamp 1644511149
transform 1 0 44252 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_15
timestamp 1644511149
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_27
timestamp 1644511149
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_39
timestamp 1644511149
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1644511149
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1644511149
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_93
timestamp 1644511149
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1644511149
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1644511149
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_125
timestamp 1644511149
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_137
timestamp 1644511149
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_149
timestamp 1644511149
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1644511149
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1644511149
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_67_175
timestamp 1644511149
transform 1 0 17204 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_187
timestamp 1644511149
transform 1 0 18308 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_67_201
timestamp 1644511149
transform 1 0 19596 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_210
timestamp 1644511149
transform 1 0 20424 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_222
timestamp 1644511149
transform 1 0 21528 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_67_225
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_242
timestamp 1644511149
transform 1 0 23368 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_250
timestamp 1644511149
transform 1 0 24104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_257
timestamp 1644511149
transform 1 0 24748 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_266
timestamp 1644511149
transform 1 0 25576 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_275
timestamp 1644511149
transform 1 0 26404 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1644511149
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_287
timestamp 1644511149
transform 1 0 27508 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_294
timestamp 1644511149
transform 1 0 28152 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_306
timestamp 1644511149
transform 1 0 29256 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_324
timestamp 1644511149
transform 1 0 30912 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_331
timestamp 1644511149
transform 1 0 31556 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1644511149
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_337
timestamp 1644511149
transform 1 0 32108 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_67_353
timestamp 1644511149
transform 1 0 33580 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_357
timestamp 1644511149
transform 1 0 33948 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_361
timestamp 1644511149
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_373
timestamp 1644511149
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_388
timestamp 1644511149
transform 1 0 36800 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_399
timestamp 1644511149
transform 1 0 37812 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_407
timestamp 1644511149
transform 1 0 38548 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_414
timestamp 1644511149
transform 1 0 39192 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_425
timestamp 1644511149
transform 1 0 40204 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1644511149
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1644511149
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_449
timestamp 1644511149
transform 1 0 42412 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_457
timestamp 1644511149
transform 1 0 43148 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_462
timestamp 1644511149
transform 1 0 43608 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_469
timestamp 1644511149
transform 1 0 44252 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_15
timestamp 1644511149
transform 1 0 2484 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_68_21
timestamp 1644511149
transform 1 0 3036 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1644511149
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_32
timestamp 1644511149
transform 1 0 4048 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_68_50
timestamp 1644511149
transform 1 0 5704 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_62
timestamp 1644511149
transform 1 0 6808 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_74
timestamp 1644511149
transform 1 0 7912 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_82
timestamp 1644511149
transform 1 0 8648 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_97
timestamp 1644511149
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_109
timestamp 1644511149
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_121
timestamp 1644511149
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1644511149
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1644511149
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_153
timestamp 1644511149
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_165
timestamp 1644511149
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_177
timestamp 1644511149
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1644511149
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1644511149
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_205
timestamp 1644511149
transform 1 0 19964 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_209
timestamp 1644511149
transform 1 0 20332 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_226
timestamp 1644511149
transform 1 0 21896 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_238
timestamp 1644511149
transform 1 0 23000 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_250
timestamp 1644511149
transform 1 0 24104 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_68_257
timestamp 1644511149
transform 1 0 24748 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_271
timestamp 1644511149
transform 1 0 26036 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_283
timestamp 1644511149
transform 1 0 27140 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_303
timestamp 1644511149
transform 1 0 28980 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1644511149
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_309
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_318
timestamp 1644511149
transform 1 0 30360 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_338
timestamp 1644511149
transform 1 0 32200 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_342
timestamp 1644511149
transform 1 0 32568 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_350
timestamp 1644511149
transform 1 0 33304 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_354
timestamp 1644511149
transform 1 0 33672 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_360
timestamp 1644511149
transform 1 0 34224 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_372
timestamp 1644511149
transform 1 0 35328 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_384
timestamp 1644511149
transform 1 0 36432 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_392
timestamp 1644511149
transform 1 0 37168 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_397
timestamp 1644511149
transform 1 0 37628 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_409
timestamp 1644511149
transform 1 0 38732 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_416
timestamp 1644511149
transform 1 0 39376 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_427
timestamp 1644511149
transform 1 0 40388 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_435
timestamp 1644511149
transform 1 0 41124 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_442
timestamp 1644511149
transform 1 0 41768 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_469
timestamp 1644511149
transform 1 0 44252 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_3
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_69_30
timestamp 1644511149
transform 1 0 3864 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_36
timestamp 1644511149
transform 1 0 4416 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_49
timestamp 1644511149
transform 1 0 5612 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1644511149
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1644511149
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1644511149
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1644511149
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_93
timestamp 1644511149
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1644511149
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1644511149
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_69_113
timestamp 1644511149
transform 1 0 11500 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_128
timestamp 1644511149
transform 1 0 12880 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_140
timestamp 1644511149
transform 1 0 13984 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_152
timestamp 1644511149
transform 1 0 15088 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_164
timestamp 1644511149
transform 1 0 16192 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_169
timestamp 1644511149
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_181
timestamp 1644511149
transform 1 0 17756 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_189
timestamp 1644511149
transform 1 0 18492 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_207
timestamp 1644511149
transform 1 0 20148 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_214
timestamp 1644511149
transform 1 0 20792 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_222
timestamp 1644511149
transform 1 0 21528 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_225
timestamp 1644511149
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_237
timestamp 1644511149
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_265
timestamp 1644511149
transform 1 0 25484 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_69_277
timestamp 1644511149
transform 1 0 26588 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_297
timestamp 1644511149
transform 1 0 28428 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_69_309
timestamp 1644511149
transform 1 0 29532 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_317
timestamp 1644511149
transform 1 0 30268 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_327
timestamp 1644511149
transform 1 0 31188 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1644511149
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_342
timestamp 1644511149
transform 1 0 32568 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_353
timestamp 1644511149
transform 1 0 33580 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_361
timestamp 1644511149
transform 1 0 34316 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_379
timestamp 1644511149
transform 1 0 35972 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1644511149
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_409
timestamp 1644511149
transform 1 0 38732 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_420
timestamp 1644511149
transform 1 0 39744 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_69_444
timestamp 1644511149
transform 1 0 41952 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_449
timestamp 1644511149
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_461
timestamp 1644511149
transform 1 0 43516 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_465
timestamp 1644511149
transform 1 0 43884 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_70_3
timestamp 1644511149
transform 1 0 1380 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_9
timestamp 1644511149
transform 1 0 1932 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_13
timestamp 1644511149
transform 1 0 2300 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_20
timestamp 1644511149
transform 1 0 2944 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_29
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_34
timestamp 1644511149
transform 1 0 4232 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_58
timestamp 1644511149
transform 1 0 6440 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_71
timestamp 1644511149
transform 1 0 7636 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1644511149
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_100
timestamp 1644511149
transform 1 0 10304 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_112
timestamp 1644511149
transform 1 0 11408 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_128
timestamp 1644511149
transform 1 0 12880 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_135
timestamp 1644511149
transform 1 0 13524 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1644511149
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_141
timestamp 1644511149
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_153
timestamp 1644511149
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_165
timestamp 1644511149
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_177
timestamp 1644511149
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1644511149
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1644511149
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_197
timestamp 1644511149
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_209
timestamp 1644511149
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_221
timestamp 1644511149
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_233
timestamp 1644511149
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1644511149
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1644511149
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_253
timestamp 1644511149
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_265
timestamp 1644511149
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_277
timestamp 1644511149
transform 1 0 26588 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_285
timestamp 1644511149
transform 1 0 27324 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_291
timestamp 1644511149
transform 1 0 27876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_303
timestamp 1644511149
transform 1 0 28980 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1644511149
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_309
timestamp 1644511149
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_321
timestamp 1644511149
transform 1 0 30636 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_327
timestamp 1644511149
transform 1 0 31188 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_335
timestamp 1644511149
transform 1 0 31924 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_340
timestamp 1644511149
transform 1 0 32384 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_360
timestamp 1644511149
transform 1 0 34224 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_365
timestamp 1644511149
transform 1 0 34684 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_372
timestamp 1644511149
transform 1 0 35328 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_384
timestamp 1644511149
transform 1 0 36432 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_70_394
timestamp 1644511149
transform 1 0 37352 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_70_416
timestamp 1644511149
transform 1 0 39376 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_424
timestamp 1644511149
transform 1 0 40112 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_432
timestamp 1644511149
transform 1 0 40848 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_444
timestamp 1644511149
transform 1 0 41952 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_469
timestamp 1644511149
transform 1 0 44252 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_3
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_8
timestamp 1644511149
transform 1 0 1840 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_15
timestamp 1644511149
transform 1 0 2484 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_22
timestamp 1644511149
transform 1 0 3128 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_29
timestamp 1644511149
transform 1 0 3772 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_71_49
timestamp 1644511149
transform 1 0 5612 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1644511149
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_60
timestamp 1644511149
transform 1 0 6624 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_72
timestamp 1644511149
transform 1 0 7728 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_96
timestamp 1644511149
transform 1 0 9936 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_71_108
timestamp 1644511149
transform 1 0 11040 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_113
timestamp 1644511149
transform 1 0 11500 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_137
timestamp 1644511149
transform 1 0 13708 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_144
timestamp 1644511149
transform 1 0 14352 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_156
timestamp 1644511149
transform 1 0 15456 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_169
timestamp 1644511149
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_181
timestamp 1644511149
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_193
timestamp 1644511149
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_205
timestamp 1644511149
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1644511149
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1644511149
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_225
timestamp 1644511149
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_237
timestamp 1644511149
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_249
timestamp 1644511149
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_261
timestamp 1644511149
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1644511149
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1644511149
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_281
timestamp 1644511149
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_293
timestamp 1644511149
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_305
timestamp 1644511149
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_317
timestamp 1644511149
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1644511149
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1644511149
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_337
timestamp 1644511149
transform 1 0 32108 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_347
timestamp 1644511149
transform 1 0 33028 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_354
timestamp 1644511149
transform 1 0 33672 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_366
timestamp 1644511149
transform 1 0 34776 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_378
timestamp 1644511149
transform 1 0 35880 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_390
timestamp 1644511149
transform 1 0 36984 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_71_393
timestamp 1644511149
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_405
timestamp 1644511149
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_417
timestamp 1644511149
transform 1 0 39468 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_71_444
timestamp 1644511149
transform 1 0 41952 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_71_449
timestamp 1644511149
transform 1 0 42412 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_455
timestamp 1644511149
transform 1 0 42964 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_462
timestamp 1644511149
transform 1 0 43608 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_469
timestamp 1644511149
transform 1 0 44252 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_24
timestamp 1644511149
transform 1 0 3312 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_32
timestamp 1644511149
transform 1 0 4048 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_38
timestamp 1644511149
transform 1 0 4600 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_60
timestamp 1644511149
transform 1 0 6624 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_72
timestamp 1644511149
transform 1 0 7728 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_85
timestamp 1644511149
transform 1 0 8924 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_93
timestamp 1644511149
transform 1 0 9660 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_72_99
timestamp 1644511149
transform 1 0 10212 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_105
timestamp 1644511149
transform 1 0 10764 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_115
timestamp 1644511149
transform 1 0 11684 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_131
timestamp 1644511149
transform 1 0 13156 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1644511149
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_141
timestamp 1644511149
transform 1 0 14076 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_148
timestamp 1644511149
transform 1 0 14720 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_155
timestamp 1644511149
transform 1 0 15364 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_167
timestamp 1644511149
transform 1 0 16468 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_179
timestamp 1644511149
transform 1 0 17572 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_191
timestamp 1644511149
transform 1 0 18676 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1644511149
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_197
timestamp 1644511149
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_209
timestamp 1644511149
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_221
timestamp 1644511149
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_233
timestamp 1644511149
transform 1 0 22540 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_237
timestamp 1644511149
transform 1 0 22908 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_244
timestamp 1644511149
transform 1 0 23552 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_256
timestamp 1644511149
transform 1 0 24656 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_268
timestamp 1644511149
transform 1 0 25760 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_280
timestamp 1644511149
transform 1 0 26864 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_295
timestamp 1644511149
transform 1 0 28244 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1644511149
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_309
timestamp 1644511149
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_321
timestamp 1644511149
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_333
timestamp 1644511149
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_345
timestamp 1644511149
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1644511149
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1644511149
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_368
timestamp 1644511149
transform 1 0 34960 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_372
timestamp 1644511149
transform 1 0 35328 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_394
timestamp 1644511149
transform 1 0 37352 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_401
timestamp 1644511149
transform 1 0 37996 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_408
timestamp 1644511149
transform 1 0 38640 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_424
timestamp 1644511149
transform 1 0 40112 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_436
timestamp 1644511149
transform 1 0 41216 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_469
timestamp 1644511149
transform 1 0 44252 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_3
timestamp 1644511149
transform 1 0 1380 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_7
timestamp 1644511149
transform 1 0 1748 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_29
timestamp 1644511149
transform 1 0 3772 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_37
timestamp 1644511149
transform 1 0 4508 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_42
timestamp 1644511149
transform 1 0 4968 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_49
timestamp 1644511149
transform 1 0 5612 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1644511149
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_78
timestamp 1644511149
transform 1 0 8280 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_90
timestamp 1644511149
transform 1 0 9384 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_94
timestamp 1644511149
transform 1 0 9752 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_98
timestamp 1644511149
transform 1 0 10120 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_104
timestamp 1644511149
transform 1 0 10672 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_108
timestamp 1644511149
transform 1 0 11040 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_113
timestamp 1644511149
transform 1 0 11500 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_117
timestamp 1644511149
transform 1 0 11868 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_139
timestamp 1644511149
transform 1 0 13892 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_164
timestamp 1644511149
transform 1 0 16192 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_169
timestamp 1644511149
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_181
timestamp 1644511149
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_193
timestamp 1644511149
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_205
timestamp 1644511149
transform 1 0 19964 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_213
timestamp 1644511149
transform 1 0 20700 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1644511149
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1644511149
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_225
timestamp 1644511149
transform 1 0 21804 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_233
timestamp 1644511149
transform 1 0 22540 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_255
timestamp 1644511149
transform 1 0 24564 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_267
timestamp 1644511149
transform 1 0 25668 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_73_276
timestamp 1644511149
transform 1 0 26496 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_284
timestamp 1644511149
transform 1 0 27232 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_73_311
timestamp 1644511149
transform 1 0 29716 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_319
timestamp 1644511149
transform 1 0 30452 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_323
timestamp 1644511149
transform 1 0 30820 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1644511149
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_337
timestamp 1644511149
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_352
timestamp 1644511149
transform 1 0 33488 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_356
timestamp 1644511149
transform 1 0 33856 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_378
timestamp 1644511149
transform 1 0 35880 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1644511149
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1644511149
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_393
timestamp 1644511149
transform 1 0 37260 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_397
timestamp 1644511149
transform 1 0 37628 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_401
timestamp 1644511149
transform 1 0 37996 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_423
timestamp 1644511149
transform 1 0 40020 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_435
timestamp 1644511149
transform 1 0 41124 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1644511149
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_449
timestamp 1644511149
transform 1 0 42412 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_454
timestamp 1644511149
transform 1 0 42872 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_461
timestamp 1644511149
transform 1 0 43516 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_468
timestamp 1644511149
transform 1 0 44160 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_472
timestamp 1644511149
transform 1 0 44528 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_24
timestamp 1644511149
transform 1 0 3312 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_29
timestamp 1644511149
transform 1 0 3772 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_36
timestamp 1644511149
transform 1 0 4416 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_61
timestamp 1644511149
transform 1 0 6716 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_68
timestamp 1644511149
transform 1 0 7360 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_80
timestamp 1644511149
transform 1 0 8464 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_85
timestamp 1644511149
transform 1 0 8924 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_110
timestamp 1644511149
transform 1 0 11224 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_135
timestamp 1644511149
transform 1 0 13524 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1644511149
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_74_141
timestamp 1644511149
transform 1 0 14076 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_74_165
timestamp 1644511149
transform 1 0 16284 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_172
timestamp 1644511149
transform 1 0 16928 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_184
timestamp 1644511149
transform 1 0 18032 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_197
timestamp 1644511149
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_209
timestamp 1644511149
transform 1 0 20332 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_213
timestamp 1644511149
transform 1 0 20700 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_235
timestamp 1644511149
transform 1 0 22724 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_243
timestamp 1644511149
transform 1 0 23460 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_248
timestamp 1644511149
transform 1 0 23920 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_274
timestamp 1644511149
transform 1 0 26312 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_299
timestamp 1644511149
transform 1 0 28612 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1644511149
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_309
timestamp 1644511149
transform 1 0 29532 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_317
timestamp 1644511149
transform 1 0 30268 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_340
timestamp 1644511149
transform 1 0 32384 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_74_351
timestamp 1644511149
transform 1 0 33396 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_360
timestamp 1644511149
transform 1 0 34224 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_365
timestamp 1644511149
transform 1 0 34684 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_74_376
timestamp 1644511149
transform 1 0 35696 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_383
timestamp 1644511149
transform 1 0 36340 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_408
timestamp 1644511149
transform 1 0 38640 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_421
timestamp 1644511149
transform 1 0 39836 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_443
timestamp 1644511149
transform 1 0 41860 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_447
timestamp 1644511149
transform 1 0 42228 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_469
timestamp 1644511149
transform 1 0 44252 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_3
timestamp 1644511149
transform 1 0 1380 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_13
timestamp 1644511149
transform 1 0 2300 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_20
timestamp 1644511149
transform 1 0 2944 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_75_50
timestamp 1644511149
transform 1 0 5704 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_60
timestamp 1644511149
transform 1 0 6624 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_72
timestamp 1644511149
transform 1 0 7728 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_77
timestamp 1644511149
transform 1 0 8188 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_83
timestamp 1644511149
transform 1 0 8740 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_85
timestamp 1644511149
transform 1 0 8924 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_97
timestamp 1644511149
transform 1 0 10028 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_75_108
timestamp 1644511149
transform 1 0 11040 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_113
timestamp 1644511149
transform 1 0 11500 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_118
timestamp 1644511149
transform 1 0 11960 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_125
timestamp 1644511149
transform 1 0 12604 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_129
timestamp 1644511149
transform 1 0 12972 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_133
timestamp 1644511149
transform 1 0 13340 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_139
timestamp 1644511149
transform 1 0 13892 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_162
timestamp 1644511149
transform 1 0 16008 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_169
timestamp 1644511149
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_181
timestamp 1644511149
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_193
timestamp 1644511149
transform 1 0 18860 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_197
timestamp 1644511149
transform 1 0 19228 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_209
timestamp 1644511149
transform 1 0 20332 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_213
timestamp 1644511149
transform 1 0 20700 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1644511149
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1644511149
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_225
timestamp 1644511149
transform 1 0 21804 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_233
timestamp 1644511149
transform 1 0 22540 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_237
timestamp 1644511149
transform 1 0 22908 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_244
timestamp 1644511149
transform 1 0 23552 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_75_274
timestamp 1644511149
transform 1 0 26312 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_75_281
timestamp 1644511149
transform 1 0 26956 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_289
timestamp 1644511149
transform 1 0 27692 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_296
timestamp 1644511149
transform 1 0 28336 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_309
timestamp 1644511149
transform 1 0 29532 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_317
timestamp 1644511149
transform 1 0 30268 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_75_322
timestamp 1644511149
transform 1 0 30728 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_334
timestamp 1644511149
transform 1 0 31832 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_337
timestamp 1644511149
transform 1 0 32108 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_360
timestamp 1644511149
transform 1 0 34224 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_365
timestamp 1644511149
transform 1 0 34684 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_377
timestamp 1644511149
transform 1 0 35788 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_389
timestamp 1644511149
transform 1 0 36892 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_393
timestamp 1644511149
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_405
timestamp 1644511149
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_417
timestamp 1644511149
transform 1 0 39468 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_75_421
timestamp 1644511149
transform 1 0 39836 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_75_426
timestamp 1644511149
transform 1 0 40296 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_438
timestamp 1644511149
transform 1 0 41400 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_446
timestamp 1644511149
transform 1 0 42136 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_449
timestamp 1644511149
transform 1 0 42412 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_453
timestamp 1644511149
transform 1 0 42780 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_457
timestamp 1644511149
transform 1 0 43148 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_461
timestamp 1644511149
transform 1 0 43516 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_465
timestamp 1644511149
transform 1 0 43884 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 44896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 44896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 44896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 44896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 44896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 44896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 44896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 44896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 44896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 44896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 44896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 44896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 44896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 44896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 44896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 44896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 44896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 44896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 44896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 44896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 44896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 44896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 44896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 44896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 44896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 44896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 44896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 44896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 44896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 44896 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 44896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 44896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 44896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 44896 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 44896 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 44896 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 44896 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 44896 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 44896 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 44896 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 44896 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 44896 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 44896 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 44896 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 44896 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 44896 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 44896 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 44896 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 44896 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 44896 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 44896 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 44896 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 44896 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 44896 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 44896 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 44896 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 44896 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 44896 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 44896 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 44896 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 44896 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 44896 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 44896 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 44896 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 44896 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 44896 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 44896 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 44896 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 44896 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 44896 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 44896 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 44896 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1644511149
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1644511149
transform -1 0 44896 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1644511149
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1644511149
transform -1 0 44896 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1644511149
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1644511149
transform -1 0 44896 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1644511149
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1644511149
transform -1 0 44896 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 3680 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1644511149
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1644511149
transform 1 0 8832 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1644511149
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1644511149
transform 1 0 13984 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1644511149
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1644511149
transform 1 0 19136 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1644511149
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1644511149
transform 1 0 24288 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1644511149
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1644511149
transform 1 0 29440 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1644511149
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1644511149
transform 1 0 34592 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1644511149
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1644511149
transform 1 0 39744 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1644511149
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0951_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11316 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  _0952_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12052 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_8  _0953_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9292 0 1 40256
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _0954_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 43516 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0955_
timestamp 1644511149
transform 1 0 20792 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0956_
timestamp 1644511149
transform 1 0 43424 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0957_
timestamp 1644511149
transform -1 0 3036 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0958_
timestamp 1644511149
transform 1 0 43424 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0959_
timestamp 1644511149
transform 1 0 8832 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0960_
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0961_
timestamp 1644511149
transform -1 0 4600 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0962_
timestamp 1644511149
transform 1 0 30544 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0963_
timestamp 1644511149
transform 1 0 43884 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0964_
timestamp 1644511149
transform 1 0 43332 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0965_
timestamp 1644511149
transform 1 0 10672 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  _0966_
timestamp 1644511149
transform 1 0 11776 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0967_
timestamp 1644511149
transform 1 0 5336 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0968_
timestamp 1644511149
transform -1 0 40940 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0969_
timestamp 1644511149
transform -1 0 2484 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0970_
timestamp 1644511149
transform 1 0 42780 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp 1644511149
transform -1 0 2392 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0972_
timestamp 1644511149
transform 1 0 12052 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0973_
timestamp 1644511149
transform 1 0 43332 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0974_
timestamp 1644511149
transform 1 0 41676 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0975_
timestamp 1644511149
transform -1 0 12328 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0976_
timestamp 1644511149
transform -1 0 28244 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0977_
timestamp 1644511149
transform 1 0 43332 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0978_
timestamp 1644511149
transform 1 0 11776 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0979_
timestamp 1644511149
transform -1 0 2668 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0980_
timestamp 1644511149
transform 1 0 43332 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0981_
timestamp 1644511149
transform 1 0 4692 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0982_
timestamp 1644511149
transform -1 0 43056 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0983_
timestamp 1644511149
transform -1 0 2668 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0984_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 11684 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0985_
timestamp 1644511149
transform -1 0 2208 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0986_
timestamp 1644511149
transform -1 0 4048 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0987_
timestamp 1644511149
transform -1 0 10212 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0988_
timestamp 1644511149
transform 1 0 42780 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0989_
timestamp 1644511149
transform -1 0 2208 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _0990_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11868 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _0991_
timestamp 1644511149
transform 1 0 36524 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0992_
timestamp 1644511149
transform -1 0 3128 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0993_
timestamp 1644511149
transform 1 0 43240 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0994_
timestamp 1644511149
transform -1 0 43056 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0995_
timestamp 1644511149
transform 1 0 23276 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0996_
timestamp 1644511149
transform 1 0 3864 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  _0997_
timestamp 1644511149
transform 1 0 4508 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0998_
timestamp 1644511149
transform 1 0 22632 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0999_
timestamp 1644511149
transform -1 0 4508 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1000_
timestamp 1644511149
transform -1 0 4048 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1001_
timestamp 1644511149
transform 1 0 42872 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1002_
timestamp 1644511149
transform 1 0 13064 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1003_
timestamp 1644511149
transform -1 0 5612 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1004_
timestamp 1644511149
transform -1 0 33488 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1005_
timestamp 1644511149
transform 1 0 11776 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1006_
timestamp 1644511149
transform 1 0 38180 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1007_
timestamp 1644511149
transform -1 0 12604 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1008_
timestamp 1644511149
transform -1 0 3312 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1009_
timestamp 1644511149
transform 1 0 6808 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1010_
timestamp 1644511149
transform 1 0 34868 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1011_
timestamp 1644511149
transform -1 0 5612 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1012_
timestamp 1644511149
transform 1 0 43332 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1013_
timestamp 1644511149
transform 1 0 43332 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1014_
timestamp 1644511149
transform 1 0 14444 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1015_
timestamp 1644511149
transform -1 0 5704 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1016_
timestamp 1644511149
transform 1 0 43516 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1017_
timestamp 1644511149
transform 1 0 43516 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1018_
timestamp 1644511149
transform 1 0 43516 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1019_
timestamp 1644511149
transform -1 0 3128 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1020_
timestamp 1644511149
transform -1 0 2392 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _1021_
timestamp 1644511149
transform 1 0 4600 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _1022_
timestamp 1644511149
transform -1 0 2300 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1023_
timestamp 1644511149
transform 1 0 43332 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1024_
timestamp 1644511149
transform -1 0 2116 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1025_
timestamp 1644511149
transform 1 0 43976 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1026_
timestamp 1644511149
transform 1 0 24380 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1027_
timestamp 1644511149
transform 1 0 5336 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _1028_
timestamp 1644511149
transform -1 0 5888 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1029_
timestamp 1644511149
transform -1 0 6624 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1030_
timestamp 1644511149
transform -1 0 15916 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1031_
timestamp 1644511149
transform 1 0 37352 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1032_
timestamp 1644511149
transform -1 0 21068 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1033_
timestamp 1644511149
transform -1 0 36524 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1034_
timestamp 1644511149
transform 1 0 6072 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1035_
timestamp 1644511149
transform 1 0 43332 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1036_
timestamp 1644511149
transform -1 0 42872 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1037_
timestamp 1644511149
transform -1 0 27232 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1038_
timestamp 1644511149
transform -1 0 3036 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1039_
timestamp 1644511149
transform 1 0 43332 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1040_
timestamp 1644511149
transform 1 0 6072 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1041_
timestamp 1644511149
transform 1 0 36524 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1042_
timestamp 1644511149
transform -1 0 2484 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1043_
timestamp 1644511149
transform -1 0 34960 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1044_
timestamp 1644511149
transform -1 0 19504 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1045_
timestamp 1644511149
transform -1 0 2944 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _1046_
timestamp 1644511149
transform 1 0 6716 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _1047_
timestamp 1644511149
transform -1 0 24840 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1048_
timestamp 1644511149
transform 1 0 42964 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1049_
timestamp 1644511149
transform -1 0 29808 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1050_
timestamp 1644511149
transform -1 0 2852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1051_
timestamp 1644511149
transform -1 0 37996 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1052_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1053_
timestamp 1644511149
transform -1 0 3036 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1054_
timestamp 1644511149
transform 1 0 42412 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1055_
timestamp 1644511149
transform 1 0 42412 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1056_
timestamp 1644511149
transform 1 0 41676 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1057_
timestamp 1644511149
transform -1 0 4048 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1058_
timestamp 1644511149
transform 1 0 13248 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1059_
timestamp 1644511149
transform -1 0 43332 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1060_
timestamp 1644511149
transform 1 0 38272 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1061_
timestamp 1644511149
transform -1 0 13340 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1062_
timestamp 1644511149
transform 1 0 13340 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1063_
timestamp 1644511149
transform 1 0 43240 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1064_
timestamp 1644511149
transform 1 0 12052 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1065_
timestamp 1644511149
transform -1 0 3128 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1066_
timestamp 1644511149
transform -1 0 43700 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1067_
timestamp 1644511149
transform -1 0 43700 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1068_
timestamp 1644511149
transform 1 0 43884 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1069_
timestamp 1644511149
transform 1 0 9200 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1070_
timestamp 1644511149
transform 1 0 12236 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1071_
timestamp 1644511149
transform 1 0 10764 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1072_
timestamp 1644511149
transform -1 0 2392 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1073_
timestamp 1644511149
transform 1 0 3404 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1074_
timestamp 1644511149
transform 1 0 14076 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1075_
timestamp 1644511149
transform -1 0 2392 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1076_
timestamp 1644511149
transform -1 0 12880 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1077_
timestamp 1644511149
transform -1 0 23092 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1078_
timestamp 1644511149
transform 1 0 43332 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1079_
timestamp 1644511149
transform 1 0 43332 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1080_
timestamp 1644511149
transform 1 0 16928 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1081_
timestamp 1644511149
transform -1 0 3036 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1082_
timestamp 1644511149
transform 1 0 23644 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1083_
timestamp 1644511149
transform 1 0 39836 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1084_
timestamp 1644511149
transform -1 0 8372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1085_
timestamp 1644511149
transform 1 0 26864 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1086_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28428 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1087_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27600 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__nor4_1  _1088_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 26220 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1089_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 27232 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1090_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26864 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_2  _1091_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29164 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1092_
timestamp 1644511149
transform -1 0 37536 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1093_
timestamp 1644511149
transform 1 0 27692 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1094_
timestamp 1644511149
transform 1 0 27508 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1095_
timestamp 1644511149
transform -1 0 28428 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__nor2b_1  _1096_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 30452 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1097_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29992 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1098_
timestamp 1644511149
transform 1 0 30820 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1099_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 30452 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1100_
timestamp 1644511149
transform 1 0 32844 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1101_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 28704 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1102_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28336 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1103_
timestamp 1644511149
transform 1 0 29348 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1104_
timestamp 1644511149
transform -1 0 30636 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1105_
timestamp 1644511149
transform -1 0 31648 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1106_
timestamp 1644511149
transform 1 0 29808 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _1107_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 29440 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1108_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 27048 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _1109_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 28060 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1110_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26036 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1111_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 25944 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1112_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28428 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1113_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30820 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__o22ai_1  _1114_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31832 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1115_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30544 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1116_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31280 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1117_
timestamp 1644511149
transform 1 0 30360 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1118_
timestamp 1644511149
transform 1 0 34592 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1119_
timestamp 1644511149
transform 1 0 29532 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _1120_
timestamp 1644511149
transform 1 0 31004 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1121_
timestamp 1644511149
transform 1 0 28520 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1122_
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _1123_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 27692 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1124_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1125_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 29256 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _1126_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 31372 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1127_
timestamp 1644511149
transform 1 0 32384 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1128_
timestamp 1644511149
transform -1 0 32844 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1129_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 32568 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1130_
timestamp 1644511149
transform -1 0 32384 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1131_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 27968 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1132_
timestamp 1644511149
transform -1 0 29072 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1133_
timestamp 1644511149
transform 1 0 30820 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1134_
timestamp 1644511149
transform -1 0 28888 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1135_
timestamp 1644511149
transform 1 0 25024 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1136_
timestamp 1644511149
transform 1 0 24656 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1137_
timestamp 1644511149
transform -1 0 25300 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o22ai_1  _1138_
timestamp 1644511149
transform -1 0 29992 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1139_
timestamp 1644511149
transform 1 0 33304 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1140_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30360 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1141_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 31832 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1142_
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1143_
timestamp 1644511149
transform -1 0 32384 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1144_
timestamp 1644511149
transform 1 0 32384 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1145_
timestamp 1644511149
transform -1 0 32108 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _1146_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30544 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1147_
timestamp 1644511149
transform 1 0 29808 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _1148_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30728 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1149_
timestamp 1644511149
transform 1 0 30820 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1150_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 31648 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _1151_
timestamp 1644511149
transform 1 0 25668 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1152_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 26404 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1153_
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1154_
timestamp 1644511149
transform 1 0 28244 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or3_2  _1155_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26772 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _1156_
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _1157_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32844 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _1158_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26680 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1159_
timestamp 1644511149
transform -1 0 37076 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _1160_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32752 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1161_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_2  _1162_
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1163_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1164_
timestamp 1644511149
transform 1 0 32844 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1165_
timestamp 1644511149
transform 1 0 32844 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1166_
timestamp 1644511149
transform 1 0 33672 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1167_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1168_
timestamp 1644511149
transform 1 0 35696 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1169_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 36248 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1170_
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1171_
timestamp 1644511149
transform 1 0 35788 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1172_
timestamp 1644511149
transform 1 0 35788 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1173_
timestamp 1644511149
transform 1 0 37444 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1174_
timestamp 1644511149
transform -1 0 37536 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1175_
timestamp 1644511149
transform 1 0 36708 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1176_
timestamp 1644511149
transform -1 0 37260 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1177_
timestamp 1644511149
transform 1 0 37628 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__xor2_1  _1178_
timestamp 1644511149
transform 1 0 36800 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1179_
timestamp 1644511149
transform 1 0 38548 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1180_
timestamp 1644511149
transform 1 0 37628 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1181_
timestamp 1644511149
transform -1 0 38732 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1182_
timestamp 1644511149
transform -1 0 37720 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1183_
timestamp 1644511149
transform -1 0 28152 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1184_
timestamp 1644511149
transform -1 0 27232 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1185_
timestamp 1644511149
transform -1 0 26496 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1186_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1187_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 28336 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1188_
timestamp 1644511149
transform 1 0 32200 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1189_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33396 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1190_
timestamp 1644511149
transform 1 0 32752 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _1191_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 32752 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1192_
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1193_
timestamp 1644511149
transform 1 0 31096 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1194_
timestamp 1644511149
transform 1 0 32384 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1195_
timestamp 1644511149
transform 1 0 37536 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1196_
timestamp 1644511149
transform -1 0 36800 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1197_
timestamp 1644511149
transform -1 0 38640 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1198_
timestamp 1644511149
transform 1 0 39008 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _1199_
timestamp 1644511149
transform 1 0 35512 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1200_
timestamp 1644511149
transform -1 0 39836 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1201_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 37628 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1202_
timestamp 1644511149
transform 1 0 38088 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _1203_
timestamp 1644511149
transform -1 0 36892 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1204_
timestamp 1644511149
transform -1 0 36156 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1205_
timestamp 1644511149
transform 1 0 33580 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1206_
timestamp 1644511149
transform 1 0 33120 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _1207_
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1208_
timestamp 1644511149
transform 1 0 33764 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1209_
timestamp 1644511149
transform -1 0 38180 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1210_
timestamp 1644511149
transform 1 0 36064 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1211_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 36064 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1212_
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1213_
timestamp 1644511149
transform 1 0 38916 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1214_
timestamp 1644511149
transform 1 0 37352 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1215_
timestamp 1644511149
transform -1 0 34224 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1216_
timestamp 1644511149
transform 1 0 34960 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1217_
timestamp 1644511149
transform 1 0 36156 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1218_
timestamp 1644511149
transform -1 0 36800 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1219_
timestamp 1644511149
transform 1 0 38824 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1220_
timestamp 1644511149
transform 1 0 34868 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1221_
timestamp 1644511149
transform 1 0 33948 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1222_
timestamp 1644511149
transform -1 0 32752 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1223_
timestamp 1644511149
transform 1 0 35236 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1224_
timestamp 1644511149
transform 1 0 38548 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1225_
timestamp 1644511149
transform -1 0 38180 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1226_
timestamp 1644511149
transform 1 0 37996 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1227_
timestamp 1644511149
transform -1 0 39192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1228_
timestamp 1644511149
transform 1 0 37352 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1229_
timestamp 1644511149
transform 1 0 35880 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1230_
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1231_
timestamp 1644511149
transform 1 0 33120 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1232_
timestamp 1644511149
transform 1 0 35512 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1233_
timestamp 1644511149
transform -1 0 36800 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1234_
timestamp 1644511149
transform 1 0 35880 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1235_
timestamp 1644511149
transform 1 0 35604 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1236_
timestamp 1644511149
transform 1 0 35328 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1237_
timestamp 1644511149
transform 1 0 36156 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1238_
timestamp 1644511149
transform -1 0 39008 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1239_
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1240_
timestamp 1644511149
transform 1 0 36984 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1241_
timestamp 1644511149
transform -1 0 36616 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1242_
timestamp 1644511149
transform 1 0 37812 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1243_
timestamp 1644511149
transform 1 0 37628 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1244_
timestamp 1644511149
transform -1 0 38364 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1245_
timestamp 1644511149
transform -1 0 39468 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1246_
timestamp 1644511149
transform -1 0 39376 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1247_
timestamp 1644511149
transform -1 0 17664 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1248_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17572 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1249_
timestamp 1644511149
transform -1 0 20608 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1250_
timestamp 1644511149
transform 1 0 20516 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1251_
timestamp 1644511149
transform 1 0 22448 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1252_
timestamp 1644511149
transform 1 0 22172 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1253_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22908 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1254_
timestamp 1644511149
transform 1 0 40112 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1255_
timestamp 1644511149
transform -1 0 39376 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1256_
timestamp 1644511149
transform 1 0 38732 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1257_
timestamp 1644511149
transform 1 0 42412 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1258_
timestamp 1644511149
transform 1 0 42412 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1259_
timestamp 1644511149
transform -1 0 39376 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1260_
timestamp 1644511149
transform 1 0 39192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1261_
timestamp 1644511149
transform -1 0 41952 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1262_
timestamp 1644511149
transform -1 0 41124 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1263_
timestamp 1644511149
transform 1 0 40664 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1264_
timestamp 1644511149
transform 1 0 42412 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1265_
timestamp 1644511149
transform 1 0 40388 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1266_
timestamp 1644511149
transform -1 0 41584 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1267_
timestamp 1644511149
transform -1 0 19412 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1268_
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1269_
timestamp 1644511149
transform 1 0 18768 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _1270_
timestamp 1644511149
transform -1 0 18492 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1271_
timestamp 1644511149
transform -1 0 23736 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1272_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 18584 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1273_
timestamp 1644511149
transform -1 0 14076 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1274_
timestamp 1644511149
transform 1 0 15824 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1275_
timestamp 1644511149
transform 1 0 17112 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1276_
timestamp 1644511149
transform 1 0 18492 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1277_
timestamp 1644511149
transform 1 0 20424 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1278_
timestamp 1644511149
transform 1 0 17480 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1279_
timestamp 1644511149
transform -1 0 20976 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1280_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19320 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1281_
timestamp 1644511149
transform 1 0 17388 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__or3_1  _1282_
timestamp 1644511149
transform 1 0 17572 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1283_
timestamp 1644511149
transform -1 0 18676 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1284_
timestamp 1644511149
transform 1 0 13248 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1285_
timestamp 1644511149
transform 1 0 28520 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1286_
timestamp 1644511149
transform 1 0 38732 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1287_
timestamp 1644511149
transform -1 0 40204 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_1  _1288_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 38456 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1289_
timestamp 1644511149
transform -1 0 39376 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nor3b_1  _1290_
timestamp 1644511149
transform 1 0 37996 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1291_
timestamp 1644511149
transform 1 0 27784 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1292_
timestamp 1644511149
transform -1 0 28888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1293_
timestamp 1644511149
transform 1 0 28060 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1294_
timestamp 1644511149
transform -1 0 28428 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1295_
timestamp 1644511149
transform 1 0 22356 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1296_
timestamp 1644511149
transform -1 0 23368 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1297_
timestamp 1644511149
transform -1 0 18768 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1298_
timestamp 1644511149
transform 1 0 18308 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1299_
timestamp 1644511149
transform -1 0 18768 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_2  _1300_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 18400 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1301_
timestamp 1644511149
transform -1 0 18768 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1302_
timestamp 1644511149
transform 1 0 19688 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _1303_
timestamp 1644511149
transform 1 0 20516 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1304_
timestamp 1644511149
transform -1 0 21252 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1305_
timestamp 1644511149
transform -1 0 17664 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1306_
timestamp 1644511149
transform -1 0 19964 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1307_
timestamp 1644511149
transform 1 0 19596 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1308_
timestamp 1644511149
transform 1 0 22724 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1309_
timestamp 1644511149
transform 1 0 21896 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1310_
timestamp 1644511149
transform -1 0 23920 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1311_
timestamp 1644511149
transform -1 0 18584 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1312_
timestamp 1644511149
transform 1 0 17572 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1313_
timestamp 1644511149
transform -1 0 17940 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1314_
timestamp 1644511149
transform 1 0 17480 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1315_
timestamp 1644511149
transform 1 0 19872 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1316_
timestamp 1644511149
transform 1 0 20424 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1317_
timestamp 1644511149
transform -1 0 20700 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1318_
timestamp 1644511149
transform -1 0 19872 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1319_
timestamp 1644511149
transform 1 0 22724 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1320_
timestamp 1644511149
transform -1 0 22172 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1321_
timestamp 1644511149
transform -1 0 21436 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1322_
timestamp 1644511149
transform -1 0 23460 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1323_
timestamp 1644511149
transform 1 0 20792 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1324_
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1325_
timestamp 1644511149
transform 1 0 20884 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1326_
timestamp 1644511149
transform 1 0 22724 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1327_
timestamp 1644511149
transform -1 0 22080 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1328_
timestamp 1644511149
transform -1 0 19964 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1329_
timestamp 1644511149
transform 1 0 20792 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1330_
timestamp 1644511149
transform 1 0 19780 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1331_
timestamp 1644511149
transform -1 0 16928 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1332_
timestamp 1644511149
transform -1 0 19964 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1333_
timestamp 1644511149
transform -1 0 19780 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1334_
timestamp 1644511149
transform -1 0 32384 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1335_
timestamp 1644511149
transform -1 0 26404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1336_
timestamp 1644511149
transform 1 0 33948 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1337_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 41952 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _1338_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 38180 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _1339_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 38548 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1340_
timestamp 1644511149
transform -1 0 40296 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1341_
timestamp 1644511149
transform -1 0 34316 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1342_
timestamp 1644511149
transform -1 0 30360 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1343_
timestamp 1644511149
transform -1 0 33948 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _1344_
timestamp 1644511149
transform 1 0 32844 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _1345_
timestamp 1644511149
transform -1 0 36064 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1346_
timestamp 1644511149
transform 1 0 33396 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _1347_
timestamp 1644511149
transform 1 0 34316 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1348_
timestamp 1644511149
transform 1 0 30360 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1349_
timestamp 1644511149
transform 1 0 31280 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1350_
timestamp 1644511149
transform 1 0 30636 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1351_
timestamp 1644511149
transform 1 0 30912 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1352_
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1353_
timestamp 1644511149
transform -1 0 30820 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1354_
timestamp 1644511149
transform -1 0 31556 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1355_
timestamp 1644511149
transform 1 0 29808 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1356_
timestamp 1644511149
transform 1 0 29900 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1357_
timestamp 1644511149
transform 1 0 32108 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1358_
timestamp 1644511149
transform -1 0 33028 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1359_
timestamp 1644511149
transform 1 0 33028 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _1360_
timestamp 1644511149
transform 1 0 32936 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1361_
timestamp 1644511149
transform -1 0 33672 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1362_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32660 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1363_
timestamp 1644511149
transform 1 0 33304 0 1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1364_
timestamp 1644511149
transform 1 0 33764 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1365_
timestamp 1644511149
transform 1 0 34684 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1366_
timestamp 1644511149
transform -1 0 35328 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1367_
timestamp 1644511149
transform 1 0 35052 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1368_
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1369_
timestamp 1644511149
transform -1 0 35052 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1370_
timestamp 1644511149
transform -1 0 34224 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1371_
timestamp 1644511149
transform -1 0 35420 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1372_
timestamp 1644511149
transform 1 0 33856 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1373_
timestamp 1644511149
transform -1 0 35512 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1374_
timestamp 1644511149
transform 1 0 30912 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1375_
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1376_
timestamp 1644511149
transform -1 0 33856 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1377_
timestamp 1644511149
transform 1 0 32476 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1378_
timestamp 1644511149
transform -1 0 32660 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1379_
timestamp 1644511149
transform -1 0 33120 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1380_
timestamp 1644511149
transform 1 0 31280 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1381_
timestamp 1644511149
transform -1 0 32844 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1382_
timestamp 1644511149
transform 1 0 33212 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1383_
timestamp 1644511149
transform 1 0 31924 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1384_
timestamp 1644511149
transform 1 0 31372 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1385_
timestamp 1644511149
transform 1 0 32660 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1386_
timestamp 1644511149
transform -1 0 32660 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1387_
timestamp 1644511149
transform 1 0 32660 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1388_
timestamp 1644511149
transform 1 0 33488 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1389_
timestamp 1644511149
transform -1 0 35696 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1390_
timestamp 1644511149
transform 1 0 33948 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1391_
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1392_
timestamp 1644511149
transform -1 0 36248 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1393_
timestamp 1644511149
transform -1 0 35696 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1394_
timestamp 1644511149
transform 1 0 35236 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1395_
timestamp 1644511149
transform -1 0 36892 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1396_
timestamp 1644511149
transform -1 0 37812 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1397_
timestamp 1644511149
transform 1 0 36064 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1398_
timestamp 1644511149
transform 1 0 36616 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1399_
timestamp 1644511149
transform 1 0 36064 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1400_
timestamp 1644511149
transform 1 0 37352 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1401_
timestamp 1644511149
transform 1 0 37076 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1402_
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1403_
timestamp 1644511149
transform -1 0 38916 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1404_
timestamp 1644511149
transform -1 0 37628 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1405_
timestamp 1644511149
transform -1 0 36800 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1406_
timestamp 1644511149
transform 1 0 38180 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1407_
timestamp 1644511149
transform -1 0 39192 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1408_
timestamp 1644511149
transform 1 0 38364 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1409_
timestamp 1644511149
transform -1 0 39376 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1410_
timestamp 1644511149
transform 1 0 39468 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1411_
timestamp 1644511149
transform -1 0 40388 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1412_
timestamp 1644511149
transform -1 0 41124 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1413_
timestamp 1644511149
transform 1 0 38456 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1414_
timestamp 1644511149
transform 1 0 40296 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1415_
timestamp 1644511149
transform -1 0 39928 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1416_
timestamp 1644511149
transform 1 0 39100 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1417_
timestamp 1644511149
transform 1 0 41492 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1418_
timestamp 1644511149
transform -1 0 41584 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1419_
timestamp 1644511149
transform 1 0 41492 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1420_
timestamp 1644511149
transform -1 0 42872 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1421_
timestamp 1644511149
transform -1 0 43608 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1422_
timestamp 1644511149
transform -1 0 41952 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1423_
timestamp 1644511149
transform -1 0 41952 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1424_
timestamp 1644511149
transform 1 0 40756 0 -1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1425_
timestamp 1644511149
transform 1 0 42412 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1426_
timestamp 1644511149
transform -1 0 41308 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1427_
timestamp 1644511149
transform 1 0 41492 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1428_
timestamp 1644511149
transform -1 0 41124 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1429_
timestamp 1644511149
transform -1 0 40848 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1430_
timestamp 1644511149
transform -1 0 39376 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1431_
timestamp 1644511149
transform 1 0 39836 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1432_
timestamp 1644511149
transform 1 0 39100 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1433_
timestamp 1644511149
transform 1 0 39836 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1434_
timestamp 1644511149
transform 1 0 39560 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1435_
timestamp 1644511149
transform 1 0 38824 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1436_
timestamp 1644511149
transform 1 0 39836 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1437_
timestamp 1644511149
transform -1 0 37628 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1438_
timestamp 1644511149
transform -1 0 37352 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1439_
timestamp 1644511149
transform 1 0 37260 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1440_
timestamp 1644511149
transform 1 0 36984 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1441_
timestamp 1644511149
transform -1 0 37720 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1442_
timestamp 1644511149
transform 1 0 36524 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1443_
timestamp 1644511149
transform 1 0 25300 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1444_
timestamp 1644511149
transform -1 0 24012 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1445_
timestamp 1644511149
transform 1 0 23276 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1446_
timestamp 1644511149
transform -1 0 24656 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1447_
timestamp 1644511149
transform 1 0 23276 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1448_
timestamp 1644511149
transform -1 0 23920 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1449_
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1450_
timestamp 1644511149
transform -1 0 25024 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1451_
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1452_
timestamp 1644511149
transform -1 0 25300 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1453_
timestamp 1644511149
transform 1 0 24104 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1454_
timestamp 1644511149
transform -1 0 25668 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1455_
timestamp 1644511149
transform 1 0 23644 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1456_
timestamp 1644511149
transform 1 0 24564 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1457_
timestamp 1644511149
transform 1 0 25668 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1458_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 25760 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1459_
timestamp 1644511149
transform -1 0 22540 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1460_
timestamp 1644511149
transform 1 0 23000 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1461_
timestamp 1644511149
transform -1 0 24656 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1462_
timestamp 1644511149
transform 1 0 30820 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _1463_
timestamp 1644511149
transform 1 0 22724 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1464_
timestamp 1644511149
transform -1 0 26312 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1465_
timestamp 1644511149
transform -1 0 22080 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1466_
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1467_
timestamp 1644511149
transform -1 0 21988 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _1468_
timestamp 1644511149
transform -1 0 22356 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1469_
timestamp 1644511149
transform 1 0 23000 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1470_
timestamp 1644511149
transform -1 0 23644 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a21boi_1  _1471_
timestamp 1644511149
transform -1 0 24932 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1472_
timestamp 1644511149
transform -1 0 17388 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1473_
timestamp 1644511149
transform 1 0 20148 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1474_
timestamp 1644511149
transform 1 0 19964 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1475_
timestamp 1644511149
transform -1 0 21068 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1476_
timestamp 1644511149
transform 1 0 20700 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1477_
timestamp 1644511149
transform -1 0 21160 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1478_
timestamp 1644511149
transform 1 0 20700 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1479_
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1480_
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1481_
timestamp 1644511149
transform -1 0 23092 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1482_
timestamp 1644511149
transform 1 0 17204 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1483_
timestamp 1644511149
transform -1 0 20884 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1484_
timestamp 1644511149
transform 1 0 19872 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1485_
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1486_
timestamp 1644511149
transform -1 0 23276 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1487_
timestamp 1644511149
transform -1 0 16192 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1488_
timestamp 1644511149
transform -1 0 20516 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1489_
timestamp 1644511149
transform 1 0 20884 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1490_
timestamp 1644511149
transform -1 0 22356 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1491_
timestamp 1644511149
transform 1 0 15916 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1492_
timestamp 1644511149
transform -1 0 19688 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a21boi_1  _1493_
timestamp 1644511149
transform -1 0 19780 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1494_
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1495_
timestamp 1644511149
transform 1 0 20240 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1496_
timestamp 1644511149
transform -1 0 20700 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1497_
timestamp 1644511149
transform -1 0 19872 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1498_
timestamp 1644511149
transform -1 0 21620 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1499_
timestamp 1644511149
transform -1 0 17204 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1500_
timestamp 1644511149
transform 1 0 16652 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1501_
timestamp 1644511149
transform 1 0 17572 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1502_
timestamp 1644511149
transform -1 0 18216 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1503_
timestamp 1644511149
transform -1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1504_
timestamp 1644511149
transform -1 0 17940 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1505_
timestamp 1644511149
transform -1 0 16192 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1506_
timestamp 1644511149
transform 1 0 20424 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1507_
timestamp 1644511149
transform 1 0 15456 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1508_
timestamp 1644511149
transform -1 0 18584 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1509_
timestamp 1644511149
transform 1 0 17940 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1510_
timestamp 1644511149
transform 1 0 17480 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _1511_
timestamp 1644511149
transform -1 0 19412 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1512_
timestamp 1644511149
transform -1 0 19504 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1513_
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1514_
timestamp 1644511149
transform 1 0 18124 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_2  _1515_
timestamp 1644511149
transform -1 0 18768 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1516_
timestamp 1644511149
transform 1 0 18124 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1517_
timestamp 1644511149
transform 1 0 29900 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _1518_
timestamp 1644511149
transform -1 0 25944 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1519_
timestamp 1644511149
transform 1 0 19136 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1520_
timestamp 1644511149
transform 1 0 20056 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1521_
timestamp 1644511149
transform -1 0 19320 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1522_
timestamp 1644511149
transform 1 0 17848 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1523_
timestamp 1644511149
transform 1 0 15732 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1524_
timestamp 1644511149
transform -1 0 15456 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1525_
timestamp 1644511149
transform 1 0 14536 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1526_
timestamp 1644511149
transform 1 0 15180 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1527_
timestamp 1644511149
transform 1 0 15916 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1528_
timestamp 1644511149
transform -1 0 14904 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1529_
timestamp 1644511149
transform -1 0 14076 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1530_
timestamp 1644511149
transform 1 0 14996 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1531_
timestamp 1644511149
transform 1 0 14628 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1532_
timestamp 1644511149
transform -1 0 17296 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1533_
timestamp 1644511149
transform 1 0 15272 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1534_
timestamp 1644511149
transform -1 0 17112 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _1535_
timestamp 1644511149
transform -1 0 18216 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1536_
timestamp 1644511149
transform -1 0 17388 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1537_
timestamp 1644511149
transform -1 0 15824 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1538_
timestamp 1644511149
transform -1 0 20332 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1539_
timestamp 1644511149
transform -1 0 16928 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1540_
timestamp 1644511149
transform -1 0 16192 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1541_
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1542_
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1543_
timestamp 1644511149
transform -1 0 19596 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1544_
timestamp 1644511149
transform 1 0 17204 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_2  _1545_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17020 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__o31a_1  _1546_
timestamp 1644511149
transform -1 0 18032 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1547_
timestamp 1644511149
transform -1 0 27784 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1548_
timestamp 1644511149
transform -1 0 27692 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1549_
timestamp 1644511149
transform 1 0 25668 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1550_
timestamp 1644511149
transform 1 0 23276 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1551_
timestamp 1644511149
transform 1 0 25852 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_2  _1552_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 26220 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1553_
timestamp 1644511149
transform 1 0 25116 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1554_
timestamp 1644511149
transform 1 0 18400 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1555_
timestamp 1644511149
transform 1 0 18032 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1556_
timestamp 1644511149
transform -1 0 18400 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_1  _1557_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17848 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1558_
timestamp 1644511149
transform 1 0 22816 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1559_
timestamp 1644511149
transform -1 0 17112 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1560_
timestamp 1644511149
transform 1 0 17204 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1561_
timestamp 1644511149
transform 1 0 17112 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1562_
timestamp 1644511149
transform -1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1563_
timestamp 1644511149
transform -1 0 16836 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1564_
timestamp 1644511149
transform -1 0 18492 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1565_
timestamp 1644511149
transform -1 0 16192 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _1566_
timestamp 1644511149
transform -1 0 18400 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1567_
timestamp 1644511149
transform -1 0 17848 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1568_
timestamp 1644511149
transform -1 0 15640 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1569_
timestamp 1644511149
transform -1 0 17664 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1570_
timestamp 1644511149
transform 1 0 16836 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1571_
timestamp 1644511149
transform 1 0 16284 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1572_
timestamp 1644511149
transform 1 0 16100 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1573_
timestamp 1644511149
transform -1 0 15272 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1574_
timestamp 1644511149
transform 1 0 14260 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1575_
timestamp 1644511149
transform 1 0 16928 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1576_
timestamp 1644511149
transform -1 0 16836 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1577_
timestamp 1644511149
transform 1 0 17480 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _1578_
timestamp 1644511149
transform -1 0 18216 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1579_
timestamp 1644511149
transform -1 0 19320 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1580_
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1581_
timestamp 1644511149
transform 1 0 17848 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1582_
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1583_
timestamp 1644511149
transform 1 0 15732 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1584_
timestamp 1644511149
transform 1 0 16376 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1585_
timestamp 1644511149
transform -1 0 19872 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1586_
timestamp 1644511149
transform -1 0 18584 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1587_
timestamp 1644511149
transform -1 0 17388 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1588_
timestamp 1644511149
transform -1 0 19136 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1589_
timestamp 1644511149
transform 1 0 17664 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1590_
timestamp 1644511149
transform -1 0 15824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1591_
timestamp 1644511149
transform 1 0 26312 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1592_
timestamp 1644511149
transform 1 0 15916 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1593_
timestamp 1644511149
transform 1 0 16192 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _1594_
timestamp 1644511149
transform -1 0 26404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1595_
timestamp 1644511149
transform -1 0 26128 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1596_
timestamp 1644511149
transform 1 0 17848 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1597_
timestamp 1644511149
transform -1 0 19504 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1598_
timestamp 1644511149
transform 1 0 18216 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1599_
timestamp 1644511149
transform -1 0 18952 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1600_
timestamp 1644511149
transform -1 0 16192 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1601_
timestamp 1644511149
transform -1 0 18768 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1602_
timestamp 1644511149
transform -1 0 26128 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _1603_
timestamp 1644511149
transform -1 0 18584 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1604_
timestamp 1644511149
transform -1 0 19688 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1605_
timestamp 1644511149
transform -1 0 17112 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1606_
timestamp 1644511149
transform 1 0 15824 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1607_
timestamp 1644511149
transform -1 0 16192 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1608_
timestamp 1644511149
transform 1 0 15916 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _1609_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15456 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1610_
timestamp 1644511149
transform 1 0 23552 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1611_
timestamp 1644511149
transform -1 0 19688 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1612_
timestamp 1644511149
transform -1 0 21344 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1613_
timestamp 1644511149
transform 1 0 22080 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1614_
timestamp 1644511149
transform -1 0 23736 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _1615_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20884 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__o31a_1  _1616_
timestamp 1644511149
transform 1 0 19780 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1617_
timestamp 1644511149
transform 1 0 18400 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1618_
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1619_
timestamp 1644511149
transform -1 0 17940 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_1  _1620_
timestamp 1644511149
transform -1 0 17204 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1621_
timestamp 1644511149
transform 1 0 17020 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1622_
timestamp 1644511149
transform 1 0 18124 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1623_
timestamp 1644511149
transform 1 0 18400 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1624_
timestamp 1644511149
transform -1 0 17204 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1625_
timestamp 1644511149
transform 1 0 20976 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1626_
timestamp 1644511149
transform 1 0 19320 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _1627_
timestamp 1644511149
transform 1 0 18584 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1628_
timestamp 1644511149
transform 1 0 20976 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1629_
timestamp 1644511149
transform 1 0 20148 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1630_
timestamp 1644511149
transform 1 0 19320 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1631_
timestamp 1644511149
transform -1 0 19596 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1632_
timestamp 1644511149
transform -1 0 19964 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1633_
timestamp 1644511149
transform 1 0 19964 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1634_
timestamp 1644511149
transform -1 0 20792 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1635_
timestamp 1644511149
transform 1 0 17756 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1636_
timestamp 1644511149
transform 1 0 20148 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1637_
timestamp 1644511149
transform 1 0 20976 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1638_
timestamp 1644511149
transform 1 0 18492 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o221ai_1  _1639_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20424 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1640_
timestamp 1644511149
transform -1 0 22816 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1641_
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1642_
timestamp 1644511149
transform 1 0 22080 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1643_
timestamp 1644511149
transform -1 0 21344 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1644_
timestamp 1644511149
transform 1 0 20240 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1645_
timestamp 1644511149
transform -1 0 21344 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1646_
timestamp 1644511149
transform 1 0 19780 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1647_
timestamp 1644511149
transform 1 0 19504 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1648_
timestamp 1644511149
transform 1 0 19780 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1649_
timestamp 1644511149
transform -1 0 22448 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1650_
timestamp 1644511149
transform 1 0 22816 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1651_
timestamp 1644511149
transform -1 0 23460 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1652_
timestamp 1644511149
transform -1 0 24104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1653_
timestamp 1644511149
transform 1 0 22724 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1654_
timestamp 1644511149
transform -1 0 23736 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1655_
timestamp 1644511149
transform -1 0 22724 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1656_
timestamp 1644511149
transform -1 0 24840 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1657_
timestamp 1644511149
transform 1 0 23276 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1658_
timestamp 1644511149
transform -1 0 23552 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1659_
timestamp 1644511149
transform 1 0 22356 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1660_
timestamp 1644511149
transform 1 0 22448 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1661_
timestamp 1644511149
transform 1 0 22172 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1662_
timestamp 1644511149
transform -1 0 22908 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1663_
timestamp 1644511149
transform 1 0 25668 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _1664_
timestamp 1644511149
transform 1 0 27508 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _1665_
timestamp 1644511149
transform 1 0 27324 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1666_
timestamp 1644511149
transform -1 0 26496 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1667_
timestamp 1644511149
transform 1 0 26128 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1668_
timestamp 1644511149
transform 1 0 25576 0 -1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1669_
timestamp 1644511149
transform -1 0 25760 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1670_
timestamp 1644511149
transform -1 0 25116 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_1  _1671_
timestamp 1644511149
transform -1 0 23920 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1672_
timestamp 1644511149
transform 1 0 24380 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1673_
timestamp 1644511149
transform 1 0 25116 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1674_
timestamp 1644511149
transform 1 0 25392 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1675_
timestamp 1644511149
transform -1 0 24748 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1676_
timestamp 1644511149
transform 1 0 28060 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1677_
timestamp 1644511149
transform 1 0 25852 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1678_
timestamp 1644511149
transform -1 0 25484 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1679_
timestamp 1644511149
transform -1 0 22356 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1680_
timestamp 1644511149
transform 1 0 25944 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1681_
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1682_
timestamp 1644511149
transform -1 0 26036 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1683_
timestamp 1644511149
transform 1 0 26404 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1684_
timestamp 1644511149
transform 1 0 27416 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1685_
timestamp 1644511149
transform 1 0 27876 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1686_
timestamp 1644511149
transform 1 0 26496 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1687_
timestamp 1644511149
transform -1 0 28980 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1688_
timestamp 1644511149
transform -1 0 27968 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1689_
timestamp 1644511149
transform 1 0 28244 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1690_
timestamp 1644511149
transform 1 0 28244 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1691_
timestamp 1644511149
transform 1 0 24840 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__o221ai_1  _1692_
timestamp 1644511149
transform 1 0 28612 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1693_
timestamp 1644511149
transform -1 0 28244 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1694_
timestamp 1644511149
transform -1 0 27876 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1695_
timestamp 1644511149
transform 1 0 27324 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1696_
timestamp 1644511149
transform -1 0 27232 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1697_
timestamp 1644511149
transform 1 0 24932 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1698_
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1699_
timestamp 1644511149
transform 1 0 26496 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1700_
timestamp 1644511149
transform -1 0 25300 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1701_
timestamp 1644511149
transform -1 0 25024 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1702_
timestamp 1644511149
transform 1 0 27600 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1703_
timestamp 1644511149
transform 1 0 27784 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1704_
timestamp 1644511149
transform 1 0 28612 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1705_
timestamp 1644511149
transform -1 0 29900 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1706_
timestamp 1644511149
transform 1 0 28520 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1707_
timestamp 1644511149
transform -1 0 29808 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1708_
timestamp 1644511149
transform -1 0 27324 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1709_
timestamp 1644511149
transform 1 0 27876 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1710_
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1711_
timestamp 1644511149
transform -1 0 27508 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1712_
timestamp 1644511149
transform -1 0 26496 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1713_
timestamp 1644511149
transform 1 0 27692 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1714_
timestamp 1644511149
transform -1 0 28428 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1715_
timestamp 1644511149
transform 1 0 25208 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1716_
timestamp 1644511149
transform -1 0 32384 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _1717_
timestamp 1644511149
transform -1 0 34224 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__o21bai_1  _1718_
timestamp 1644511149
transform 1 0 31556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1719_
timestamp 1644511149
transform 1 0 33488 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1720_
timestamp 1644511149
transform -1 0 35144 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1721_
timestamp 1644511149
transform -1 0 31648 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1722_
timestamp 1644511149
transform 1 0 31188 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1723_
timestamp 1644511149
transform -1 0 29716 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1724_
timestamp 1644511149
transform 1 0 30084 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _1725_
timestamp 1644511149
transform 1 0 29992 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1726_
timestamp 1644511149
transform -1 0 32292 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1727_
timestamp 1644511149
transform -1 0 31188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1728_
timestamp 1644511149
transform -1 0 32476 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1729_
timestamp 1644511149
transform 1 0 30452 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1730_
timestamp 1644511149
transform 1 0 31188 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1731_
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1732_
timestamp 1644511149
transform 1 0 30176 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1733_
timestamp 1644511149
transform -1 0 32568 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1734_
timestamp 1644511149
transform 1 0 29992 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _1735_
timestamp 1644511149
transform 1 0 30912 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1736_
timestamp 1644511149
transform -1 0 32752 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1737_
timestamp 1644511149
transform -1 0 31648 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1738_
timestamp 1644511149
transform -1 0 32384 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1739_
timestamp 1644511149
transform -1 0 31648 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1740_
timestamp 1644511149
transform 1 0 35144 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1741_
timestamp 1644511149
transform 1 0 28428 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1742_
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1743_
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1744_
timestamp 1644511149
transform -1 0 33856 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1745_
timestamp 1644511149
transform -1 0 34960 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1746_
timestamp 1644511149
transform 1 0 32752 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1747_
timestamp 1644511149
transform -1 0 34776 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1748_
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1749_
timestamp 1644511149
transform -1 0 36064 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1750_
timestamp 1644511149
transform -1 0 33856 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1751_
timestamp 1644511149
transform -1 0 34132 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1752_
timestamp 1644511149
transform 1 0 24196 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1753_
timestamp 1644511149
transform -1 0 24748 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1754_
timestamp 1644511149
transform -1 0 28796 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1755_
timestamp 1644511149
transform 1 0 27692 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1756_
timestamp 1644511149
transform -1 0 29624 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1757_
timestamp 1644511149
transform -1 0 27232 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1758_
timestamp 1644511149
transform -1 0 25024 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _1759_
timestamp 1644511149
transform -1 0 26496 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1760_
timestamp 1644511149
transform -1 0 25392 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1761_
timestamp 1644511149
transform -1 0 28152 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1762_
timestamp 1644511149
transform -1 0 27324 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1763_
timestamp 1644511149
transform -1 0 27968 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1764_
timestamp 1644511149
transform 1 0 28520 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1765_
timestamp 1644511149
transform 1 0 27876 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1766_
timestamp 1644511149
transform 1 0 28704 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1767_
timestamp 1644511149
transform 1 0 28060 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1768_
timestamp 1644511149
transform 1 0 28060 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1769_
timestamp 1644511149
transform -1 0 27692 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1770_
timestamp 1644511149
transform 1 0 25944 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1771_
timestamp 1644511149
transform 1 0 26128 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1772_
timestamp 1644511149
transform -1 0 26588 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1773_
timestamp 1644511149
transform -1 0 25300 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_1  _1774_
timestamp 1644511149
transform -1 0 24656 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1775_
timestamp 1644511149
transform -1 0 23644 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1776_
timestamp 1644511149
transform -1 0 23552 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1777_
timestamp 1644511149
transform -1 0 26220 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1778_
timestamp 1644511149
transform -1 0 23552 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1779_
timestamp 1644511149
transform -1 0 22908 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1780_
timestamp 1644511149
transform 1 0 22172 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1781_
timestamp 1644511149
transform -1 0 22356 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1782_
timestamp 1644511149
transform -1 0 21896 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1783_
timestamp 1644511149
transform 1 0 20792 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1784_
timestamp 1644511149
transform 1 0 20700 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_4  _1785_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25392 0 1 34816
box -38 -48 1602 592
use sky130_fd_sc_hd__xor2_1  _1786_
timestamp 1644511149
transform 1 0 24472 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1787_
timestamp 1644511149
transform 1 0 25484 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1788_
timestamp 1644511149
transform 1 0 26312 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1789_
timestamp 1644511149
transform -1 0 23920 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1790_
timestamp 1644511149
transform -1 0 23828 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1791_
timestamp 1644511149
transform 1 0 23460 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1792_
timestamp 1644511149
transform 1 0 22080 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1793_
timestamp 1644511149
transform 1 0 22908 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1794_
timestamp 1644511149
transform 1 0 22816 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1795_
timestamp 1644511149
transform 1 0 21804 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1796_
timestamp 1644511149
transform 1 0 20792 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1797_
timestamp 1644511149
transform -1 0 21436 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1798_
timestamp 1644511149
transform 1 0 19964 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1799_
timestamp 1644511149
transform 1 0 20148 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1800_
timestamp 1644511149
transform -1 0 33672 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1801_
timestamp 1644511149
transform 1 0 33580 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1802_
timestamp 1644511149
transform -1 0 34224 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1803_
timestamp 1644511149
transform 1 0 34132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1804_
timestamp 1644511149
transform 1 0 33120 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1805_
timestamp 1644511149
transform -1 0 34960 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1806_
timestamp 1644511149
transform 1 0 33580 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1807_
timestamp 1644511149
transform 1 0 32660 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1808_
timestamp 1644511149
transform 1 0 34224 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1809_
timestamp 1644511149
transform -1 0 36064 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1810_
timestamp 1644511149
transform -1 0 36708 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1811_
timestamp 1644511149
transform 1 0 35512 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1812_
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1813_
timestamp 1644511149
transform 1 0 36064 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1814_
timestamp 1644511149
transform -1 0 36800 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1815_
timestamp 1644511149
transform 1 0 29716 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1816_
timestamp 1644511149
transform 1 0 30176 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1817_
timestamp 1644511149
transform 1 0 31740 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1818_
timestamp 1644511149
transform -1 0 32384 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1819_
timestamp 1644511149
transform 1 0 30820 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _1820_
timestamp 1644511149
transform -1 0 31188 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1821_
timestamp 1644511149
transform 1 0 27600 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1822_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 40388 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1823_
timestamp 1644511149
transform 1 0 38272 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1824_
timestamp 1644511149
transform 1 0 39928 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1825_
timestamp 1644511149
transform 1 0 35420 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1826_
timestamp 1644511149
transform 1 0 31188 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1827_
timestamp 1644511149
transform 1 0 33304 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1828_
timestamp 1644511149
transform 1 0 31004 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1829_
timestamp 1644511149
transform 1 0 30912 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1830_
timestamp 1644511149
transform 1 0 37812 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1831_
timestamp 1644511149
transform -1 0 34224 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1832_
timestamp 1644511149
transform -1 0 33580 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1833_
timestamp 1644511149
transform -1 0 33580 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1834_
timestamp 1644511149
transform 1 0 28428 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1835_
timestamp 1644511149
transform 1 0 40112 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1836_
timestamp 1644511149
transform 1 0 39652 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1837_
timestamp 1644511149
transform 1 0 28796 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1838_
timestamp 1644511149
transform 1 0 30176 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1839_
timestamp 1644511149
transform 1 0 20884 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1840_
timestamp 1644511149
transform 1 0 19320 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1841_
timestamp 1644511149
transform -1 0 24196 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1842_
timestamp 1644511149
transform 1 0 17296 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1843_
timestamp 1644511149
transform 1 0 16928 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1844_
timestamp 1644511149
transform 1 0 20240 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1845_
timestamp 1644511149
transform 1 0 22172 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1846_
timestamp 1644511149
transform -1 0 23000 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1847_
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1848_
timestamp 1644511149
transform 1 0 19596 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1849_
timestamp 1644511149
transform 1 0 30728 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1850_
timestamp 1644511149
transform 1 0 29440 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1851_
timestamp 1644511149
transform -1 0 34224 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1852_
timestamp 1644511149
transform -1 0 35972 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1853_
timestamp 1644511149
transform -1 0 35696 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1854_
timestamp 1644511149
transform -1 0 36248 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1855_
timestamp 1644511149
transform -1 0 31280 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1856_
timestamp 1644511149
transform 1 0 30636 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1857_
timestamp 1644511149
transform 1 0 30544 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1858_
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1859_
timestamp 1644511149
transform -1 0 34868 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1860_
timestamp 1644511149
transform 1 0 34776 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1861_
timestamp 1644511149
transform 1 0 35972 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1862_
timestamp 1644511149
transform -1 0 38732 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1863_
timestamp 1644511149
transform 1 0 36616 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1864_
timestamp 1644511149
transform -1 0 40296 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1865_
timestamp 1644511149
transform 1 0 39928 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1866_
timestamp 1644511149
transform 1 0 38640 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1867_
timestamp 1644511149
transform 1 0 40480 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1868_
timestamp 1644511149
transform 1 0 42412 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1869_
timestamp 1644511149
transform 1 0 40480 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1870_
timestamp 1644511149
transform 1 0 40480 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1871_
timestamp 1644511149
transform -1 0 39376 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1872_
timestamp 1644511149
transform -1 0 39928 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1873_
timestamp 1644511149
transform 1 0 37260 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1874_
timestamp 1644511149
transform 1 0 36064 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1875_
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1876_
timestamp 1644511149
transform 1 0 24380 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1877_
timestamp 1644511149
transform 1 0 25024 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1878_
timestamp 1644511149
transform 1 0 25300 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1879_
timestamp 1644511149
transform 1 0 25208 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1880_
timestamp 1644511149
transform 1 0 25392 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1881_
timestamp 1644511149
transform 1 0 24288 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1882_
timestamp 1644511149
transform 1 0 26036 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1883_
timestamp 1644511149
transform 1 0 22448 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1884_
timestamp 1644511149
transform 1 0 25024 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1885_
timestamp 1644511149
transform 1 0 20976 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1886_
timestamp 1644511149
transform 1 0 21528 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1887_
timestamp 1644511149
transform 1 0 21436 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1888_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23460 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1889_
timestamp 1644511149
transform 1 0 23000 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1890_
timestamp 1644511149
transform 1 0 24840 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1891_
timestamp 1644511149
transform 1 0 23460 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1892_
timestamp 1644511149
transform 1 0 20792 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1893_
timestamp 1644511149
transform 1 0 23920 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1894_
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1895_
timestamp 1644511149
transform 1 0 15364 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1896_
timestamp 1644511149
transform 1 0 15548 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1897_
timestamp 1644511149
transform 1 0 18676 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1898_
timestamp 1644511149
transform 1 0 19596 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1899_
timestamp 1644511149
transform 1 0 14720 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1900_
timestamp 1644511149
transform 1 0 13984 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1901_
timestamp 1644511149
transform -1 0 15548 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1902_
timestamp 1644511149
transform -1 0 15548 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1903_
timestamp 1644511149
transform 1 0 17296 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1904_
timestamp 1644511149
transform -1 0 16744 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1905_
timestamp 1644511149
transform 1 0 17848 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1906_
timestamp 1644511149
transform 1 0 15548 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1907_
timestamp 1644511149
transform 1 0 14720 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1908_
timestamp 1644511149
transform 1 0 14260 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1909_
timestamp 1644511149
transform 1 0 13616 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1910_
timestamp 1644511149
transform 1 0 15364 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1911_
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1912_
timestamp 1644511149
transform -1 0 20700 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1913_
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1914_
timestamp 1644511149
transform 1 0 13892 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1915_
timestamp 1644511149
transform 1 0 15916 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1916_
timestamp 1644511149
transform 1 0 16284 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1917_
timestamp 1644511149
transform -1 0 21712 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1918_
timestamp 1644511149
transform 1 0 18676 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1919_
timestamp 1644511149
transform 1 0 20424 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1920_
timestamp 1644511149
transform 1 0 19872 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1921_
timestamp 1644511149
transform 1 0 19228 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1922_
timestamp 1644511149
transform -1 0 24196 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1923_
timestamp 1644511149
transform 1 0 21988 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1924_
timestamp 1644511149
transform 1 0 22448 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1925_
timestamp 1644511149
transform 1 0 22908 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1926_
timestamp 1644511149
transform 1 0 24012 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1927_
timestamp 1644511149
transform 1 0 21896 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1928_
timestamp 1644511149
transform 1 0 26956 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1929_
timestamp 1644511149
transform 1 0 27508 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1930_
timestamp 1644511149
transform 1 0 24656 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1931_
timestamp 1644511149
transform 1 0 24656 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1932_
timestamp 1644511149
transform -1 0 31004 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1933_
timestamp 1644511149
transform 1 0 27232 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1934_
timestamp 1644511149
transform -1 0 30084 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1935_
timestamp 1644511149
transform 1 0 32752 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1936_
timestamp 1644511149
transform -1 0 31740 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1937_
timestamp 1644511149
transform 1 0 32384 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1938_
timestamp 1644511149
transform 1 0 32752 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1939_
timestamp 1644511149
transform -1 0 36800 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1940_
timestamp 1644511149
transform -1 0 37260 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1941_
timestamp 1644511149
transform -1 0 34224 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1942_
timestamp 1644511149
transform 1 0 25668 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1943_
timestamp 1644511149
transform 1 0 27600 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1944_
timestamp 1644511149
transform 1 0 27784 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1945_
timestamp 1644511149
transform 1 0 25668 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1946_
timestamp 1644511149
transform 1 0 23092 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1947_
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1948_
timestamp 1644511149
transform 1 0 19872 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1949_
timestamp 1644511149
transform 1 0 25024 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1950_
timestamp 1644511149
transform 1 0 23644 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1951_
timestamp 1644511149
transform 1 0 21896 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1952_
timestamp 1644511149
transform 1 0 19688 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1953_
timestamp 1644511149
transform 1 0 34040 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1954_
timestamp 1644511149
transform -1 0 35144 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1955_
timestamp 1644511149
transform 1 0 33856 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1956_
timestamp 1644511149
transform 1 0 30268 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1957_
timestamp 1644511149
transform 1 0 29624 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1958_
timestamp 1644511149
transform 1 0 28336 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1959_
timestamp 1644511149
transform 1 0 28520 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1960_
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1961_
timestamp 1644511149
transform 1 0 28520 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1962_
timestamp 1644511149
transform 1 0 28704 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1963_
timestamp 1644511149
transform 1 0 28244 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1964_
timestamp 1644511149
transform 1 0 27416 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1965_
timestamp 1644511149
transform 1 0 27232 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1966_
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1967_
timestamp 1644511149
transform 1 0 35880 0 1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1968_
timestamp 1644511149
transform -1 0 29716 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1969_
timestamp 1644511149
transform -1 0 31556 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1970_
timestamp 1644511149
transform -1 0 36984 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1971_
timestamp 1644511149
transform 1 0 36432 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1972_
timestamp 1644511149
transform -1 0 27968 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1973__6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 7636 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1974__7
timestamp 1644511149
transform 1 0 1564 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1975__8
timestamp 1644511149
transform 1 0 18492 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1976__9
timestamp 1644511149
transform 1 0 1748 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1977__10
timestamp 1644511149
transform -1 0 42688 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1978__11
timestamp 1644511149
transform 1 0 2392 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1979__12
timestamp 1644511149
transform 1 0 43608 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1980__13
timestamp 1644511149
transform -1 0 4048 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1981__14
timestamp 1644511149
transform -1 0 43148 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1982__15
timestamp 1644511149
transform -1 0 43148 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1983__16
timestamp 1644511149
transform 1 0 43976 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1984__17
timestamp 1644511149
transform 1 0 19964 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1985__18
timestamp 1644511149
transform -1 0 38640 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1986__19
timestamp 1644511149
transform 1 0 4140 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1987__20
timestamp 1644511149
transform 1 0 23644 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1988__21
timestamp 1644511149
transform -1 0 1748 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1989__22
timestamp 1644511149
transform 1 0 43976 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1990__23
timestamp 1644511149
transform -1 0 43884 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1991__24
timestamp 1644511149
transform 1 0 6348 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1992__25
timestamp 1644511149
transform 1 0 43700 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1993__26
timestamp 1644511149
transform 1 0 1748 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1994__27
timestamp 1644511149
transform 1 0 43608 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1995__28
timestamp 1644511149
transform -1 0 28336 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1996__29
timestamp 1644511149
transform 1 0 12696 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1997__30
timestamp 1644511149
transform 1 0 43976 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1998__31
timestamp 1644511149
transform 1 0 1748 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1999__32
timestamp 1644511149
transform -1 0 43884 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2000__33
timestamp 1644511149
transform -1 0 3772 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2001__34
timestamp 1644511149
transform -1 0 40296 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2002__35
timestamp 1644511149
transform -1 0 6624 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2003__36
timestamp 1644511149
transform 1 0 43976 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2004__37
timestamp 1644511149
transform 1 0 43608 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2005__38
timestamp 1644511149
transform -1 0 40296 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2006__39
timestamp 1644511149
transform -1 0 30728 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2007__40
timestamp 1644511149
transform -1 0 6624 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2008__41
timestamp 1644511149
transform -1 0 2300 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2009__42
timestamp 1644511149
transform 1 0 43608 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2010__43
timestamp 1644511149
transform -1 0 21068 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2011__44
timestamp 1644511149
transform 1 0 43976 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2012__45
timestamp 1644511149
transform -1 0 2300 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2013__46
timestamp 1644511149
transform -1 0 18032 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2014__47
timestamp 1644511149
transform -1 0 2392 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2015__48
timestamp 1644511149
transform 1 0 43608 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2016__49
timestamp 1644511149
transform -1 0 2300 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2017__50
timestamp 1644511149
transform 1 0 36064 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2018__51
timestamp 1644511149
transform 1 0 1932 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2019__52
timestamp 1644511149
transform 1 0 28796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2020__53
timestamp 1644511149
transform -1 0 43884 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2021__54
timestamp 1644511149
transform -1 0 25484 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2022__55
timestamp 1644511149
transform -1 0 34224 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2023__56
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2024__57
timestamp 1644511149
transform -1 0 35696 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2025__58
timestamp 1644511149
transform -1 0 15824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2026__59
timestamp 1644511149
transform 1 0 43608 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2027__60
timestamp 1644511149
transform -1 0 2024 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2028__61
timestamp 1644511149
transform -1 0 2024 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2029__62
timestamp 1644511149
transform 1 0 2668 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2030__63
timestamp 1644511149
transform 1 0 43608 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2031__64
timestamp 1644511149
transform 1 0 43976 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2032__65
timestamp 1644511149
transform 1 0 43884 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2033__66
timestamp 1644511149
transform -1 0 15364 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2034__67
timestamp 1644511149
transform -1 0 42964 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2035__68
timestamp 1644511149
transform 1 0 24012 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2036__69
timestamp 1644511149
transform -1 0 35972 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2037__70
timestamp 1644511149
transform -1 0 16928 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2038__71
timestamp 1644511149
transform -1 0 23184 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2039__72
timestamp 1644511149
transform -1 0 44252 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2040__73
timestamp 1644511149
transform -1 0 2024 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2041__74
timestamp 1644511149
transform -1 0 42964 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2042__75
timestamp 1644511149
transform -1 0 11960 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2043__76
timestamp 1644511149
transform -1 0 4324 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2044__77
timestamp 1644511149
transform -1 0 9568 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2045__78
timestamp 1644511149
transform 1 0 1564 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2046__79
timestamp 1644511149
transform -1 0 44160 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2047__80
timestamp 1644511149
transform -1 0 43056 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2048__81
timestamp 1644511149
transform -1 0 43056 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2049__82
timestamp 1644511149
transform -1 0 5152 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2050__83
timestamp 1644511149
transform 1 0 10764 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2051__84
timestamp 1644511149
transform -1 0 39100 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2052__85
timestamp 1644511149
transform -1 0 12696 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2053__86
timestamp 1644511149
transform -1 0 33396 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2054__87
timestamp 1644511149
transform 1 0 13248 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2055__88
timestamp 1644511149
transform -1 0 43884 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2056__89
timestamp 1644511149
transform -1 0 4048 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2057__90
timestamp 1644511149
transform -1 0 4692 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2058__91
timestamp 1644511149
transform -1 0 22908 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2059__92
timestamp 1644511149
transform 1 0 23276 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2060__93
timestamp 1644511149
transform -1 0 43240 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2061__94
timestamp 1644511149
transform 1 0 43976 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2062__95
timestamp 1644511149
transform 1 0 26220 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2063__96
timestamp 1644511149
transform -1 0 37536 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2064__97
timestamp 1644511149
transform 1 0 43976 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2065__98
timestamp 1644511149
transform -1 0 7360 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2066__99
timestamp 1644511149
transform -1 0 38180 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2067__100
timestamp 1644511149
transform 1 0 2576 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2068__101
timestamp 1644511149
transform -1 0 43884 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2069__102
timestamp 1644511149
transform -1 0 10120 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2070__103
timestamp 1644511149
transform -1 0 2024 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2071__104
timestamp 1644511149
transform 1 0 1840 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2072__105
timestamp 1644511149
transform -1 0 2116 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2073_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7268 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2074_
timestamp 1644511149
transform 1 0 1840 0 -1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2075_
timestamp 1644511149
transform 1 0 18768 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2076_
timestamp 1644511149
transform 1 0 1932 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2077_
timestamp 1644511149
transform 1 0 41676 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2078_
timestamp 1644511149
transform 1 0 3496 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2079_
timestamp 1644511149
transform -1 0 44252 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2080_
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2081_
timestamp 1644511149
transform 1 0 42320 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2082_
timestamp 1644511149
transform 1 0 42320 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2083_
timestamp 1644511149
transform -1 0 44252 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2084_
timestamp 1644511149
transform 1 0 20608 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2085_
timestamp 1644511149
transform 1 0 38088 0 -1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2086_
timestamp 1644511149
transform -1 0 6716 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2087_
timestamp 1644511149
transform 1 0 24380 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2088_
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2089_
timestamp 1644511149
transform -1 0 44252 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2090_
timestamp 1644511149
transform 1 0 42320 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2091_
timestamp 1644511149
transform -1 0 6624 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2092_
timestamp 1644511149
transform -1 0 44252 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2093_
timestamp 1644511149
transform 1 0 1932 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2094_
timestamp 1644511149
transform -1 0 44252 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2095_
timestamp 1644511149
transform 1 0 27784 0 -1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2096_
timestamp 1644511149
transform -1 0 13432 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2097_
timestamp 1644511149
transform -1 0 44252 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2098_
timestamp 1644511149
transform -1 0 3312 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2099_
timestamp 1644511149
transform 1 0 42320 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2100_
timestamp 1644511149
transform -1 0 3312 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2101_
timestamp 1644511149
transform 1 0 40020 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2102_
timestamp 1644511149
transform 1 0 5336 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2103_
timestamp 1644511149
transform -1 0 44252 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2104_
timestamp 1644511149
transform -1 0 44252 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2105_
timestamp 1644511149
transform 1 0 39928 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2106_
timestamp 1644511149
transform 1 0 30452 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2107_
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2108_
timestamp 1644511149
transform 1 0 1932 0 -1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2109_
timestamp 1644511149
transform -1 0 44252 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2110_
timestamp 1644511149
transform 1 0 20792 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2111_
timestamp 1644511149
transform -1 0 44252 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2112_
timestamp 1644511149
transform 1 0 2024 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2113_
timestamp 1644511149
transform 1 0 16836 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2114_
timestamp 1644511149
transform 1 0 2024 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2115_
timestamp 1644511149
transform -1 0 44252 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2116_
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2117_
timestamp 1644511149
transform 1 0 12880 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2118_
timestamp 1644511149
transform 1 0 38180 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2119_
timestamp 1644511149
transform 1 0 42320 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2120_
timestamp 1644511149
transform -1 0 5244 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2121_
timestamp 1644511149
transform 1 0 42320 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2122_
timestamp 1644511149
transform 1 0 41584 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2123_
timestamp 1644511149
transform 1 0 41860 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2124_
timestamp 1644511149
transform 1 0 1932 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2125_
timestamp 1644511149
transform 1 0 36708 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2126_
timestamp 1644511149
transform -1 0 3312 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2127_
timestamp 1644511149
transform 1 0 29164 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2128_
timestamp 1644511149
transform 1 0 42320 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2129_
timestamp 1644511149
transform 1 0 24380 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2130_
timestamp 1644511149
transform 1 0 33948 0 -1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2131_
timestamp 1644511149
transform 1 0 1932 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2132_
timestamp 1644511149
transform 1 0 35420 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2133_
timestamp 1644511149
transform 1 0 15456 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2134_
timestamp 1644511149
transform -1 0 44252 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2135_
timestamp 1644511149
transform 1 0 1656 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2136_
timestamp 1644511149
transform 1 0 1656 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2137_
timestamp 1644511149
transform -1 0 3312 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2138_
timestamp 1644511149
transform -1 0 44252 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2139_
timestamp 1644511149
transform -1 0 44252 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2140_
timestamp 1644511149
transform -1 0 44252 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2141_
timestamp 1644511149
transform 1 0 14352 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2142_
timestamp 1644511149
transform -1 0 41952 0 -1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2143_
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2144_
timestamp 1644511149
transform 1 0 35604 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2145_
timestamp 1644511149
transform 1 0 14260 0 -1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2146_
timestamp 1644511149
transform 1 0 22080 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2147_
timestamp 1644511149
transform -1 0 41952 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2148_
timestamp 1644511149
transform 1 0 1748 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2149_
timestamp 1644511149
transform 1 0 42320 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2150_
timestamp 1644511149
transform 1 0 11592 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2151_
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2152_
timestamp 1644511149
transform 1 0 9200 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2153_
timestamp 1644511149
transform 1 0 1656 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2154_
timestamp 1644511149
transform -1 0 41952 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2155_
timestamp 1644511149
transform 1 0 42320 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2156_
timestamp 1644511149
transform -1 0 41952 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2157_
timestamp 1644511149
transform -1 0 4416 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2158_
timestamp 1644511149
transform 1 0 11960 0 -1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2159_
timestamp 1644511149
transform 1 0 38824 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2160_
timestamp 1644511149
transform 1 0 11684 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2161_
timestamp 1644511149
transform 1 0 32292 0 -1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2162_
timestamp 1644511149
transform 1 0 14076 0 -1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2163_
timestamp 1644511149
transform 1 0 42320 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2164_
timestamp 1644511149
transform 1 0 3772 0 -1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2165_
timestamp 1644511149
transform 1 0 4048 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2166_
timestamp 1644511149
transform 1 0 22632 0 -1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2167_
timestamp 1644511149
transform 1 0 24380 0 -1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2168_
timestamp 1644511149
transform -1 0 39652 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2169_
timestamp 1644511149
transform -1 0 44252 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2170_
timestamp 1644511149
transform 1 0 26680 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2171_
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2172_
timestamp 1644511149
transform -1 0 44252 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2173_
timestamp 1644511149
transform 1 0 6348 0 -1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2174_
timestamp 1644511149
transform 1 0 37352 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2175_
timestamp 1644511149
transform -1 0 3312 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2176_
timestamp 1644511149
transform 1 0 42320 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2177_
timestamp 1644511149
transform 1 0 9292 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2178_
timestamp 1644511149
transform 1 0 1656 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2179_
timestamp 1644511149
transform -1 0 3312 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _2180_
timestamp 1644511149
transform 1 0 1748 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i
timestamp 1644511149
transform -1 0 29164 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_wb_clk_i
timestamp 1644511149
transform -1 0 25668 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 29348 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_wb_clk_i
timestamp 1644511149
transform -1 0 21712 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_wb_clk_i
timestamp 1644511149
transform -1 0 24840 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 33856 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_0_0_wb_clk_i
timestamp 1644511149
transform -1 0 21804 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 22080 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_2_0_wb_clk_i
timestamp 1644511149
transform -1 0 27876 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 30360 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_4_0_wb_clk_i
timestamp 1644511149
transform -1 0 24564 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_5_0_wb_clk_i
timestamp 1644511149
transform -1 0 23920 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_6_0_wb_clk_i
timestamp 1644511149
transform -1 0 35328 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_7_0_wb_clk_i
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_0_0_wb_clk_i
timestamp 1644511149
transform -1 0 19688 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 23828 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_2_0_wb_clk_i
timestamp 1644511149
transform -1 0 20056 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 22356 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_4_0_wb_clk_i
timestamp 1644511149
transform -1 0 27416 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_5_0_wb_clk_i
timestamp 1644511149
transform 1 0 30912 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_6_0_wb_clk_i
timestamp 1644511149
transform -1 0 30268 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_7_0_wb_clk_i
timestamp 1644511149
transform 1 0 31924 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_8_0_wb_clk_i
timestamp 1644511149
transform -1 0 21528 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_9_0_wb_clk_i
timestamp 1644511149
transform 1 0 24472 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_10_0_wb_clk_i
timestamp 1644511149
transform -1 0 22356 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_11_0_wb_clk_i
timestamp 1644511149
transform 1 0 24104 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_12_0_wb_clk_i
timestamp 1644511149
transform -1 0 32936 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_13_0_wb_clk_i
timestamp 1644511149
transform 1 0 36064 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_14_0_wb_clk_i
timestamp 1644511149
transform -1 0 33488 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_15_0_wb_clk_i
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29808 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2
timestamp 1644511149
transform 1 0 30176 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  input1
timestamp 1644511149
transform 1 0 1748 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1644511149
transform -1 0 27692 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input3
timestamp 1644511149
transform -1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input4
timestamp 1644511149
transform 1 0 7820 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 1644511149
transform -1 0 44252 0 1 7616
box -38 -48 406 592
<< labels >>
rlabel metal3 s 0 42788 800 43028 6 active
port 0 nsew signal input
rlabel metal2 s 14158 0 14270 800 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 25750 45200 25862 46000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s -10 45200 102 46000 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 45200 38708 46000 38948 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 21886 0 21998 800 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 17378 45200 17490 46000 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 45200 40748 46000 40988 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 45200 3348 46000 3588 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 9650 45200 9762 46000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 10938 45200 11050 46000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 39918 0 40030 800 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 0 14908 800 15148 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 0 26468 800 26708 6 io_in[20]
port 13 nsew signal input
rlabel metal3 s 0 17628 800 17868 6 io_in[21]
port 14 nsew signal input
rlabel metal3 s 45200 14228 46000 14468 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 8362 45200 8474 46000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 5786 45200 5898 46000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 34766 0 34878 800 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 33478 0 33590 800 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 45200 10148 46000 10388 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 30258 0 30370 800 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 45714 45200 45826 46000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 14802 0 14914 800 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 45200 18308 46000 18548 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 40748 800 40988 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 28326 0 28438 800 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 23748 800 23988 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 34766 45200 34878 46000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 39918 45200 40030 46000 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 45200 28508 46000 28748 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 41206 45200 41318 46000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 26394 45200 26506 46000 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 45200 27828 46000 28068 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 45200 44148 46000 44388 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 0 28508 800 28748 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 0 19668 800 19908 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 45200 30548 46000 30788 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 7718 45200 7830 46000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 24462 0 24574 800 6 io_oeb[0]
port 39 nsew signal tristate
rlabel metal3 s 0 15588 800 15828 6 io_oeb[10]
port 40 nsew signal tristate
rlabel metal3 s 45200 25788 46000 26028 6 io_oeb[11]
port 41 nsew signal tristate
rlabel metal3 s 45200 13548 46000 13788 6 io_oeb[12]
port 42 nsew signal tristate
rlabel metal3 s 45200 12868 46000 13108 6 io_oeb[13]
port 43 nsew signal tristate
rlabel metal3 s 0 4028 800 4268 6 io_oeb[14]
port 44 nsew signal tristate
rlabel metal2 s 12870 45200 12982 46000 6 io_oeb[15]
port 45 nsew signal tristate
rlabel metal3 s 45200 1988 46000 2228 6 io_oeb[16]
port 46 nsew signal tristate
rlabel metal2 s 12226 0 12338 800 6 io_oeb[17]
port 47 nsew signal tristate
rlabel metal2 s 33478 45200 33590 46000 6 io_oeb[18]
port 48 nsew signal tristate
rlabel metal2 s 13514 45200 13626 46000 6 io_oeb[19]
port 49 nsew signal tristate
rlabel metal2 s 36054 0 36166 800 6 io_oeb[1]
port 50 nsew signal tristate
rlabel metal3 s 45200 19668 46000 19908 6 io_oeb[20]
port 51 nsew signal tristate
rlabel metal2 s 1922 45200 2034 46000 6 io_oeb[21]
port 52 nsew signal tristate
rlabel metal2 s 4498 0 4610 800 6 io_oeb[22]
port 53 nsew signal tristate
rlabel metal2 s 23174 45200 23286 46000 6 io_oeb[23]
port 54 nsew signal tristate
rlabel metal2 s 23818 45200 23930 46000 6 io_oeb[24]
port 55 nsew signal tristate
rlabel metal2 s 43782 0 43894 800 6 io_oeb[25]
port 56 nsew signal tristate
rlabel metal3 s 45200 35988 46000 36228 6 io_oeb[26]
port 57 nsew signal tristate
rlabel metal2 s 27038 45200 27150 46000 6 io_oeb[27]
port 58 nsew signal tristate
rlabel metal2 s 38630 0 38742 800 6 io_oeb[28]
port 59 nsew signal tristate
rlabel metal3 s 45200 29868 46000 30108 6 io_oeb[29]
port 60 nsew signal tristate
rlabel metal2 s 38630 45200 38742 46000 6 io_oeb[2]
port 61 nsew signal tristate
rlabel metal2 s 2566 45200 2678 46000 6 io_oeb[30]
port 62 nsew signal tristate
rlabel metal2 s 37986 0 38098 800 6 io_oeb[31]
port 63 nsew signal tristate
rlabel metal3 s 0 23068 800 23308 6 io_oeb[32]
port 64 nsew signal tristate
rlabel metal2 s 45070 0 45182 800 6 io_oeb[33]
port 65 nsew signal tristate
rlabel metal2 s 10294 45200 10406 46000 6 io_oeb[34]
port 66 nsew signal tristate
rlabel metal3 s 0 20348 800 20588 6 io_oeb[35]
port 67 nsew signal tristate
rlabel metal3 s 0 10148 800 10388 6 io_oeb[36]
port 68 nsew signal tristate
rlabel metal3 s 0 16948 800 17188 6 io_oeb[37]
port 69 nsew signal tristate
rlabel metal2 s 23174 0 23286 800 6 io_oeb[3]
port 70 nsew signal tristate
rlabel metal3 s 45200 -52 46000 188 6 io_oeb[4]
port 71 nsew signal tristate
rlabel metal3 s 0 29868 800 30108 6 io_oeb[5]
port 72 nsew signal tristate
rlabel metal3 s 45200 16268 46000 16508 6 io_oeb[6]
port 73 nsew signal tristate
rlabel metal2 s 12226 45200 12338 46000 6 io_oeb[7]
port 74 nsew signal tristate
rlabel metal2 s 3854 0 3966 800 6 io_oeb[8]
port 75 nsew signal tristate
rlabel metal2 s 9650 0 9762 800 6 io_oeb[9]
port 76 nsew signal tristate
rlabel metal3 s 45200 43468 46000 43708 6 io_out[0]
port 77 nsew signal tristate
rlabel metal3 s 45200 25108 46000 25348 6 io_out[10]
port 78 nsew signal tristate
rlabel metal3 s 0 1988 800 2228 6 io_out[11]
port 79 nsew signal tristate
rlabel metal3 s 0 6748 800 6988 6 io_out[12]
port 80 nsew signal tristate
rlabel metal2 s 37342 0 37454 800 6 io_out[13]
port 81 nsew signal tristate
rlabel metal3 s 45200 36668 46000 36908 6 io_out[14]
port 82 nsew signal tristate
rlabel metal3 s 0 38028 800 38268 6 io_out[15]
port 83 nsew signal tristate
rlabel metal3 s 45200 24428 46000 24668 6 io_out[16]
port 84 nsew signal tristate
rlabel metal2 s 42494 45200 42606 46000 6 io_out[17]
port 85 nsew signal tristate
rlabel metal2 s 43138 0 43250 800 6 io_out[18]
port 86 nsew signal tristate
rlabel metal3 s 0 22388 800 22628 6 io_out[19]
port 87 nsew signal tristate
rlabel metal2 s 30902 45200 31014 46000 6 io_out[1]
port 88 nsew signal tristate
rlabel metal2 s 37342 45200 37454 46000 6 io_out[20]
port 89 nsew signal tristate
rlabel metal3 s 0 37348 800 37588 6 io_out[21]
port 90 nsew signal tristate
rlabel metal2 s 29614 0 29726 800 6 io_out[22]
port 91 nsew signal tristate
rlabel metal3 s 45200 21028 46000 21268 6 io_out[23]
port 92 nsew signal tristate
rlabel metal2 s 25106 0 25218 800 6 io_out[24]
port 93 nsew signal tristate
rlabel metal2 s 34122 45200 34234 46000 6 io_out[25]
port 94 nsew signal tristate
rlabel metal3 s 0 4708 800 4948 6 io_out[26]
port 95 nsew signal tristate
rlabel metal2 s 36054 45200 36166 46000 6 io_out[27]
port 96 nsew signal tristate
rlabel metal2 s 16090 0 16202 800 6 io_out[28]
port 97 nsew signal tristate
rlabel metal3 s 45200 628 46000 868 6 io_out[29]
port 98 nsew signal tristate
rlabel metal2 s 6430 0 6542 800 6 io_out[2]
port 99 nsew signal tristate
rlabel metal3 s 0 6068 800 6308 6 io_out[30]
port 100 nsew signal tristate
rlabel metal3 s 0 12868 800 13108 6 io_out[31]
port 101 nsew signal tristate
rlabel metal3 s 0 43468 800 43708 6 io_out[32]
port 102 nsew signal tristate
rlabel metal3 s 45200 6068 46000 6308 6 io_out[33]
port 103 nsew signal tristate
rlabel metal3 s 45200 38028 46000 38268 6 io_out[34]
port 104 nsew signal tristate
rlabel metal3 s 45200 35308 46000 35548 6 io_out[35]
port 105 nsew signal tristate
rlabel metal2 s 14802 45200 14914 46000 6 io_out[36]
port 106 nsew signal tristate
rlabel metal3 s 45200 41428 46000 41668 6 io_out[37]
port 107 nsew signal tristate
rlabel metal3 s 0 40068 800 40308 6 io_out[3]
port 108 nsew signal tristate
rlabel metal3 s 45200 27148 46000 27388 6 io_out[4]
port 109 nsew signal tristate
rlabel metal2 s 21242 45200 21354 46000 6 io_out[5]
port 110 nsew signal tristate
rlabel metal2 s 44426 45200 44538 46000 6 io_out[6]
port 111 nsew signal tristate
rlabel metal3 s 0 18308 800 18548 6 io_out[7]
port 112 nsew signal tristate
rlabel metal2 s 17378 0 17490 800 6 io_out[8]
port 113 nsew signal tristate
rlabel metal3 s 0 14228 800 14468 6 io_out[9]
port 114 nsew signal tristate
rlabel metal3 s 45200 7428 46000 7668 6 la1_data_in[0]
port 115 nsew signal input
rlabel metal2 s 19954 0 20066 800 6 la1_data_in[10]
port 116 nsew signal input
rlabel metal3 s 45200 5388 46000 5628 6 la1_data_in[11]
port 117 nsew signal input
rlabel metal3 s 0 34628 800 34868 6 la1_data_in[12]
port 118 nsew signal input
rlabel metal2 s 30902 0 31014 800 6 la1_data_in[13]
port 119 nsew signal input
rlabel metal3 s 0 12188 800 12428 6 la1_data_in[14]
port 120 nsew signal input
rlabel metal2 s 15446 45200 15558 46000 6 la1_data_in[15]
port 121 nsew signal input
rlabel metal2 s 28970 45200 29082 46000 6 la1_data_in[16]
port 122 nsew signal input
rlabel metal2 s 22530 45200 22642 46000 6 la1_data_in[17]
port 123 nsew signal input
rlabel metal2 s 40562 0 40674 800 6 la1_data_in[18]
port 124 nsew signal input
rlabel metal2 s 16090 45200 16202 46000 6 la1_data_in[19]
port 125 nsew signal input
rlabel metal2 s 18666 0 18778 800 6 la1_data_in[1]
port 126 nsew signal input
rlabel metal3 s 0 33948 800 34188 6 la1_data_in[20]
port 127 nsew signal input
rlabel metal2 s 45070 45200 45182 46000 6 la1_data_in[21]
port 128 nsew signal input
rlabel metal3 s 45200 8108 46000 8348 6 la1_data_in[22]
port 129 nsew signal input
rlabel metal3 s 0 628 800 868 6 la1_data_in[23]
port 130 nsew signal input
rlabel metal2 s 13514 0 13626 800 6 la1_data_in[24]
port 131 nsew signal input
rlabel metal3 s 0 35308 800 35548 6 la1_data_in[25]
port 132 nsew signal input
rlabel metal3 s 45200 2668 46000 2908 6 la1_data_in[26]
port 133 nsew signal input
rlabel metal2 s 27038 0 27150 800 6 la1_data_in[27]
port 134 nsew signal input
rlabel metal3 s 0 31228 800 31468 6 la1_data_in[28]
port 135 nsew signal input
rlabel metal2 s 634 45200 746 46000 6 la1_data_in[29]
port 136 nsew signal input
rlabel metal2 s 10938 0 11050 800 6 la1_data_in[2]
port 137 nsew signal input
rlabel metal2 s 1278 0 1390 800 6 la1_data_in[30]
port 138 nsew signal input
rlabel metal2 s 35410 0 35522 800 6 la1_data_in[31]
port 139 nsew signal input
rlabel metal3 s 0 29188 800 29428 6 la1_data_in[3]
port 140 nsew signal input
rlabel metal2 s 39274 45200 39386 46000 6 la1_data_in[4]
port 141 nsew signal input
rlabel metal3 s 45200 22388 46000 22628 6 la1_data_in[5]
port 142 nsew signal input
rlabel metal2 s 18022 45200 18134 46000 6 la1_data_in[6]
port 143 nsew signal input
rlabel metal3 s 0 21028 800 21268 6 la1_data_in[7]
port 144 nsew signal input
rlabel metal2 s 18666 45200 18778 46000 6 la1_data_in[8]
port 145 nsew signal input
rlabel metal3 s 0 31908 800 32148 6 la1_data_in[9]
port 146 nsew signal input
rlabel metal2 s 7074 0 7186 800 6 la1_data_out[0]
port 147 nsew signal tristate
rlabel metal3 s 45200 10828 46000 11068 6 la1_data_out[10]
port 148 nsew signal tristate
rlabel metal2 s 21242 0 21354 800 6 la1_data_out[11]
port 149 nsew signal tristate
rlabel metal3 s 45200 42108 46000 42348 6 la1_data_out[12]
port 150 nsew signal tristate
rlabel metal2 s 4498 45200 4610 46000 6 la1_data_out[13]
port 151 nsew signal tristate
rlabel metal2 s 24462 45200 24574 46000 6 la1_data_out[14]
port 152 nsew signal tristate
rlabel metal3 s 0 1308 800 1548 6 la1_data_out[15]
port 153 nsew signal tristate
rlabel metal3 s 45200 15588 46000 15828 6 la1_data_out[16]
port 154 nsew signal tristate
rlabel metal3 s 45200 33268 46000 33508 6 la1_data_out[17]
port 155 nsew signal tristate
rlabel metal2 s 5142 45200 5254 46000 6 la1_data_out[18]
port 156 nsew signal tristate
rlabel metal3 s 45200 23068 46000 23308 6 la1_data_out[19]
port 157 nsew signal tristate
rlabel metal3 s 0 42108 800 42348 6 la1_data_out[1]
port 158 nsew signal tristate
rlabel metal3 s 0 9468 800 9708 6 la1_data_out[20]
port 159 nsew signal tristate
rlabel metal3 s 45200 39388 46000 39628 6 la1_data_out[21]
port 160 nsew signal tristate
rlabel metal2 s 28326 45200 28438 46000 6 la1_data_out[22]
port 161 nsew signal tristate
rlabel metal2 s 11582 0 11694 800 6 la1_data_out[23]
port 162 nsew signal tristate
rlabel metal3 s 45200 16948 46000 17188 6 la1_data_out[24]
port 163 nsew signal tristate
rlabel metal3 s 0 3348 800 3588 6 la1_data_out[25]
port 164 nsew signal tristate
rlabel metal3 s 45200 4708 46000 4948 6 la1_data_out[26]
port 165 nsew signal tristate
rlabel metal3 s 0 44828 800 45068 6 la1_data_out[27]
port 166 nsew signal tristate
rlabel metal2 s 41206 0 41318 800 6 la1_data_out[28]
port 167 nsew signal tristate
rlabel metal2 s 5786 0 5898 800 6 la1_data_out[29]
port 168 nsew signal tristate
rlabel metal2 s 19310 0 19422 800 6 la1_data_out[2]
port 169 nsew signal tristate
rlabel metal3 s 45200 11508 46000 11748 6 la1_data_out[30]
port 170 nsew signal tristate
rlabel metal3 s 45200 44828 46000 45068 6 la1_data_out[31]
port 171 nsew signal tristate
rlabel metal3 s 0 8788 800 9028 6 la1_data_out[3]
port 172 nsew signal tristate
rlabel metal2 s 42494 0 42606 800 6 la1_data_out[4]
port 173 nsew signal tristate
rlabel metal2 s 3210 0 3322 800 6 la1_data_out[5]
port 174 nsew signal tristate
rlabel metal3 s 45200 18988 46000 19228 6 la1_data_out[6]
port 175 nsew signal tristate
rlabel metal2 s 634 0 746 800 6 la1_data_out[7]
port 176 nsew signal tristate
rlabel metal3 s 45200 33948 46000 34188 6 la1_data_out[8]
port 177 nsew signal tristate
rlabel metal2 s 43782 45200 43894 46000 6 la1_data_out[9]
port 178 nsew signal tristate
rlabel metal2 s 45714 0 45826 800 6 la1_oenb[0]
port 179 nsew signal input
rlabel metal2 s 41850 45200 41962 46000 6 la1_oenb[10]
port 180 nsew signal input
rlabel metal3 s 0 25788 800 26028 6 la1_oenb[11]
port 181 nsew signal input
rlabel metal3 s 0 27148 800 27388 6 la1_oenb[12]
port 182 nsew signal input
rlabel metal2 s 27682 0 27794 800 6 la1_oenb[13]
port 183 nsew signal input
rlabel metal2 s -10 0 102 800 6 la1_oenb[14]
port 184 nsew signal input
rlabel metal2 s 32834 0 32946 800 6 la1_oenb[15]
port 185 nsew signal input
rlabel metal3 s 0 32588 800 32828 6 la1_oenb[16]
port 186 nsew signal input
rlabel metal2 s 3210 45200 3322 46000 6 la1_oenb[17]
port 187 nsew signal input
rlabel metal2 s 20598 45200 20710 46000 6 la1_oenb[18]
port 188 nsew signal input
rlabel metal3 s 0 24428 800 24668 6 la1_oenb[19]
port 189 nsew signal input
rlabel metal2 s 8362 0 8474 800 6 la1_oenb[1]
port 190 nsew signal input
rlabel metal2 s 1922 0 2034 800 6 la1_oenb[20]
port 191 nsew signal input
rlabel metal2 s 29614 45200 29726 46000 6 la1_oenb[21]
port 192 nsew signal input
rlabel metal2 s 19954 45200 20066 46000 6 la1_oenb[22]
port 193 nsew signal input
rlabel metal2 s 22530 0 22642 800 6 la1_oenb[23]
port 194 nsew signal input
rlabel metal2 s 36698 45200 36810 46000 6 la1_oenb[24]
port 195 nsew signal input
rlabel metal3 s 45200 8788 46000 9028 6 la1_oenb[25]
port 196 nsew signal input
rlabel metal3 s 0 36668 800 36908 6 la1_oenb[26]
port 197 nsew signal input
rlabel metal3 s 45200 32588 46000 32828 6 la1_oenb[27]
port 198 nsew signal input
rlabel metal2 s 9006 0 9118 800 6 la1_oenb[28]
port 199 nsew signal input
rlabel metal2 s 16734 0 16846 800 6 la1_oenb[29]
port 200 nsew signal input
rlabel metal3 s 0 7428 800 7668 6 la1_oenb[2]
port 201 nsew signal input
rlabel metal3 s 45200 31228 46000 31468 6 la1_oenb[30]
port 202 nsew signal input
rlabel metal2 s 25750 0 25862 800 6 la1_oenb[31]
port 203 nsew signal input
rlabel metal2 s 32190 45200 32302 46000 6 la1_oenb[3]
port 204 nsew signal input
rlabel metal2 s 31546 45200 31658 46000 6 la1_oenb[4]
port 205 nsew signal input
rlabel metal3 s 0 45508 800 45748 6 la1_oenb[5]
port 206 nsew signal input
rlabel metal2 s 7074 45200 7186 46000 6 la1_oenb[6]
port 207 nsew signal input
rlabel metal2 s 32190 0 32302 800 6 la1_oenb[7]
port 208 nsew signal input
rlabel metal3 s 0 11508 800 11748 6 la1_oenb[8]
port 209 nsew signal input
rlabel metal3 s 0 39388 800 39628 6 la1_oenb[9]
port 210 nsew signal input
rlabel metal4 s 4208 2128 4528 43568 6 vccd1
port 211 nsew power input
rlabel metal4 s 34928 2128 35248 43568 6 vccd1
port 211 nsew power input
rlabel metal4 s 19568 2128 19888 43568 6 vssd1
port 212 nsew ground input
rlabel metal3 s 45200 21708 46000 21948 6 wb_clk_i
port 213 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 46000 46000
<< end >>
