magic
tech sky130A
magscale 1 2
timestamp 1647448291
<< obsli1 >>
rect 1104 2159 42872 41361
<< obsm1 >>
rect 658 2048 43226 41392
<< metal2 >>
rect 18 43200 74 44000
rect 662 43200 718 44000
rect 1950 43200 2006 44000
rect 2594 43200 2650 44000
rect 3238 43200 3294 44000
rect 4526 43200 4582 44000
rect 5170 43200 5226 44000
rect 5814 43200 5870 44000
rect 6458 43200 6514 44000
rect 7746 43200 7802 44000
rect 8390 43200 8446 44000
rect 9034 43200 9090 44000
rect 9678 43200 9734 44000
rect 10966 43200 11022 44000
rect 11610 43200 11666 44000
rect 12254 43200 12310 44000
rect 12898 43200 12954 44000
rect 14186 43200 14242 44000
rect 14830 43200 14886 44000
rect 15474 43200 15530 44000
rect 16762 43200 16818 44000
rect 17406 43200 17462 44000
rect 18050 43200 18106 44000
rect 18694 43200 18750 44000
rect 19982 43200 20038 44000
rect 20626 43200 20682 44000
rect 21270 43200 21326 44000
rect 21914 43200 21970 44000
rect 23202 43200 23258 44000
rect 23846 43200 23902 44000
rect 24490 43200 24546 44000
rect 25134 43200 25190 44000
rect 26422 43200 26478 44000
rect 27066 43200 27122 44000
rect 27710 43200 27766 44000
rect 28354 43200 28410 44000
rect 29642 43200 29698 44000
rect 30286 43200 30342 44000
rect 30930 43200 30986 44000
rect 32218 43200 32274 44000
rect 32862 43200 32918 44000
rect 33506 43200 33562 44000
rect 34150 43200 34206 44000
rect 35438 43200 35494 44000
rect 36082 43200 36138 44000
rect 36726 43200 36782 44000
rect 37370 43200 37426 44000
rect 38658 43200 38714 44000
rect 39302 43200 39358 44000
rect 39946 43200 40002 44000
rect 40590 43200 40646 44000
rect 41878 43200 41934 44000
rect 42522 43200 42578 44000
rect 43166 43200 43222 44000
rect 43810 43200 43866 44000
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 1950 0 2006 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 23846 0 23902 800
rect 25134 0 25190 800
rect 25778 0 25834 800
rect 26422 0 26478 800
rect 27066 0 27122 800
rect 28354 0 28410 800
rect 28998 0 29054 800
rect 29642 0 29698 800
rect 30930 0 30986 800
rect 31574 0 31630 800
rect 32218 0 32274 800
rect 32862 0 32918 800
rect 34150 0 34206 800
rect 34794 0 34850 800
rect 35438 0 35494 800
rect 36082 0 36138 800
rect 37370 0 37426 800
rect 38014 0 38070 800
rect 38658 0 38714 800
rect 39302 0 39358 800
rect 40590 0 40646 800
rect 41234 0 41290 800
rect 41878 0 41934 800
rect 43166 0 43222 800
rect 43810 0 43866 800
<< obsm2 >>
rect 774 43144 1894 43330
rect 2062 43144 2538 43330
rect 2706 43144 3182 43330
rect 3350 43144 4470 43330
rect 4638 43144 5114 43330
rect 5282 43144 5758 43330
rect 5926 43144 6402 43330
rect 6570 43144 7690 43330
rect 7858 43144 8334 43330
rect 8502 43144 8978 43330
rect 9146 43144 9622 43330
rect 9790 43144 10910 43330
rect 11078 43144 11554 43330
rect 11722 43144 12198 43330
rect 12366 43144 12842 43330
rect 13010 43144 14130 43330
rect 14298 43144 14774 43330
rect 14942 43144 15418 43330
rect 15586 43144 16706 43330
rect 16874 43144 17350 43330
rect 17518 43144 17994 43330
rect 18162 43144 18638 43330
rect 18806 43144 19926 43330
rect 20094 43144 20570 43330
rect 20738 43144 21214 43330
rect 21382 43144 21858 43330
rect 22026 43144 23146 43330
rect 23314 43144 23790 43330
rect 23958 43144 24434 43330
rect 24602 43144 25078 43330
rect 25246 43144 26366 43330
rect 26534 43144 27010 43330
rect 27178 43144 27654 43330
rect 27822 43144 28298 43330
rect 28466 43144 29586 43330
rect 29754 43144 30230 43330
rect 30398 43144 30874 43330
rect 31042 43144 32162 43330
rect 32330 43144 32806 43330
rect 32974 43144 33450 43330
rect 33618 43144 34094 43330
rect 34262 43144 35382 43330
rect 35550 43144 36026 43330
rect 36194 43144 36670 43330
rect 36838 43144 37314 43330
rect 37482 43144 38602 43330
rect 38770 43144 39246 43330
rect 39414 43144 39890 43330
rect 40058 43144 40534 43330
rect 40702 43144 41822 43330
rect 41990 43144 42466 43330
rect 42634 43144 43110 43330
rect 664 856 43220 43144
rect 774 31 1250 856
rect 1418 31 1894 856
rect 2062 31 3182 856
rect 3350 31 3826 856
rect 3994 31 4470 856
rect 4638 31 5114 856
rect 5282 31 6402 856
rect 6570 31 7046 856
rect 7214 31 7690 856
rect 7858 31 8334 856
rect 8502 31 9622 856
rect 9790 31 10266 856
rect 10434 31 10910 856
rect 11078 31 11554 856
rect 11722 31 12842 856
rect 13010 31 13486 856
rect 13654 31 14130 856
rect 14298 31 15418 856
rect 15586 31 16062 856
rect 16230 31 16706 856
rect 16874 31 17350 856
rect 17518 31 18638 856
rect 18806 31 19282 856
rect 19450 31 19926 856
rect 20094 31 20570 856
rect 20738 31 21858 856
rect 22026 31 22502 856
rect 22670 31 23146 856
rect 23314 31 23790 856
rect 23958 31 25078 856
rect 25246 31 25722 856
rect 25890 31 26366 856
rect 26534 31 27010 856
rect 27178 31 28298 856
rect 28466 31 28942 856
rect 29110 31 29586 856
rect 29754 31 30874 856
rect 31042 31 31518 856
rect 31686 31 32162 856
rect 32330 31 32806 856
rect 32974 31 34094 856
rect 34262 31 34738 856
rect 34906 31 35382 856
rect 35550 31 36026 856
rect 36194 31 37314 856
rect 37482 31 37958 856
rect 38126 31 38602 856
rect 38770 31 39246 856
rect 39414 31 40534 856
rect 40702 31 41178 856
rect 41346 31 41822 856
rect 41990 31 43110 856
<< metal3 >>
rect 0 43528 800 43648
rect 0 42848 800 42968
rect 43200 42848 44000 42968
rect 43200 42168 44000 42288
rect 0 41488 800 41608
rect 43200 41488 44000 41608
rect 0 40808 800 40928
rect 0 40128 800 40248
rect 43200 40128 44000 40248
rect 0 39448 800 39568
rect 43200 39448 44000 39568
rect 43200 38768 44000 38888
rect 0 38088 800 38208
rect 43200 38088 44000 38208
rect 0 37408 800 37528
rect 0 36728 800 36848
rect 43200 36728 44000 36848
rect 0 36048 800 36168
rect 43200 36048 44000 36168
rect 43200 35368 44000 35488
rect 0 34688 800 34808
rect 43200 34688 44000 34808
rect 0 34008 800 34128
rect 0 33328 800 33448
rect 43200 33328 44000 33448
rect 0 32648 800 32768
rect 43200 32648 44000 32768
rect 43200 31968 44000 32088
rect 0 31288 800 31408
rect 43200 31288 44000 31408
rect 0 30608 800 30728
rect 0 29928 800 30048
rect 43200 29928 44000 30048
rect 43200 29248 44000 29368
rect 0 28568 800 28688
rect 43200 28568 44000 28688
rect 0 27888 800 28008
rect 0 27208 800 27328
rect 43200 27208 44000 27328
rect 0 26528 800 26648
rect 43200 26528 44000 26648
rect 43200 25848 44000 25968
rect 0 25168 800 25288
rect 43200 25168 44000 25288
rect 0 24488 800 24608
rect 0 23808 800 23928
rect 43200 23808 44000 23928
rect 0 23128 800 23248
rect 43200 23128 44000 23248
rect 43200 22448 44000 22568
rect 0 21768 800 21888
rect 43200 21768 44000 21888
rect 0 21088 800 21208
rect 0 20408 800 20528
rect 43200 20408 44000 20528
rect 0 19728 800 19848
rect 43200 19728 44000 19848
rect 43200 19048 44000 19168
rect 0 18368 800 18488
rect 43200 18368 44000 18488
rect 0 17688 800 17808
rect 0 17008 800 17128
rect 43200 17008 44000 17128
rect 0 16328 800 16448
rect 43200 16328 44000 16448
rect 43200 15648 44000 15768
rect 0 14968 800 15088
rect 43200 14968 44000 15088
rect 0 14288 800 14408
rect 0 13608 800 13728
rect 43200 13608 44000 13728
rect 43200 12928 44000 13048
rect 0 12248 800 12368
rect 43200 12248 44000 12368
rect 0 11568 800 11688
rect 0 10888 800 11008
rect 43200 10888 44000 11008
rect 0 10208 800 10328
rect 43200 10208 44000 10328
rect 43200 9528 44000 9648
rect 0 8848 800 8968
rect 43200 8848 44000 8968
rect 0 8168 800 8288
rect 0 7488 800 7608
rect 43200 7488 44000 7608
rect 0 6808 800 6928
rect 43200 6808 44000 6928
rect 43200 6128 44000 6248
rect 0 5448 800 5568
rect 43200 5448 44000 5568
rect 0 4768 800 4888
rect 0 4088 800 4208
rect 43200 4088 44000 4208
rect 0 3408 800 3528
rect 43200 3408 44000 3528
rect 43200 2728 44000 2848
rect 0 2048 800 2168
rect 43200 2048 44000 2168
rect 0 1368 800 1488
rect 0 688 800 808
rect 43200 688 44000 808
rect 43200 8 44000 128
<< obsm3 >>
rect 880 42768 43120 42941
rect 800 42368 43200 42768
rect 800 42088 43120 42368
rect 800 41688 43200 42088
rect 880 41408 43120 41688
rect 800 41008 43200 41408
rect 880 40728 43200 41008
rect 800 40328 43200 40728
rect 880 40048 43120 40328
rect 800 39648 43200 40048
rect 880 39368 43120 39648
rect 800 38968 43200 39368
rect 800 38688 43120 38968
rect 800 38288 43200 38688
rect 880 38008 43120 38288
rect 800 37608 43200 38008
rect 880 37328 43200 37608
rect 800 36928 43200 37328
rect 880 36648 43120 36928
rect 800 36248 43200 36648
rect 880 35968 43120 36248
rect 800 35568 43200 35968
rect 800 35288 43120 35568
rect 800 34888 43200 35288
rect 880 34608 43120 34888
rect 800 34208 43200 34608
rect 880 33928 43200 34208
rect 800 33528 43200 33928
rect 880 33248 43120 33528
rect 800 32848 43200 33248
rect 880 32568 43120 32848
rect 800 32168 43200 32568
rect 800 31888 43120 32168
rect 800 31488 43200 31888
rect 880 31208 43120 31488
rect 800 30808 43200 31208
rect 880 30528 43200 30808
rect 800 30128 43200 30528
rect 880 29848 43120 30128
rect 800 29448 43200 29848
rect 800 29168 43120 29448
rect 800 28768 43200 29168
rect 880 28488 43120 28768
rect 800 28088 43200 28488
rect 880 27808 43200 28088
rect 800 27408 43200 27808
rect 880 27128 43120 27408
rect 800 26728 43200 27128
rect 880 26448 43120 26728
rect 800 26048 43200 26448
rect 800 25768 43120 26048
rect 800 25368 43200 25768
rect 880 25088 43120 25368
rect 800 24688 43200 25088
rect 880 24408 43200 24688
rect 800 24008 43200 24408
rect 880 23728 43120 24008
rect 800 23328 43200 23728
rect 880 23048 43120 23328
rect 800 22648 43200 23048
rect 800 22368 43120 22648
rect 800 21968 43200 22368
rect 880 21688 43120 21968
rect 800 21288 43200 21688
rect 880 21008 43200 21288
rect 800 20608 43200 21008
rect 880 20328 43120 20608
rect 800 19928 43200 20328
rect 880 19648 43120 19928
rect 800 19248 43200 19648
rect 800 18968 43120 19248
rect 800 18568 43200 18968
rect 880 18288 43120 18568
rect 800 17888 43200 18288
rect 880 17608 43200 17888
rect 800 17208 43200 17608
rect 880 16928 43120 17208
rect 800 16528 43200 16928
rect 880 16248 43120 16528
rect 800 15848 43200 16248
rect 800 15568 43120 15848
rect 800 15168 43200 15568
rect 880 14888 43120 15168
rect 800 14488 43200 14888
rect 880 14208 43200 14488
rect 800 13808 43200 14208
rect 880 13528 43120 13808
rect 800 13128 43200 13528
rect 800 12848 43120 13128
rect 800 12448 43200 12848
rect 880 12168 43120 12448
rect 800 11768 43200 12168
rect 880 11488 43200 11768
rect 800 11088 43200 11488
rect 880 10808 43120 11088
rect 800 10408 43200 10808
rect 880 10128 43120 10408
rect 800 9728 43200 10128
rect 800 9448 43120 9728
rect 800 9048 43200 9448
rect 880 8768 43120 9048
rect 800 8368 43200 8768
rect 880 8088 43200 8368
rect 800 7688 43200 8088
rect 880 7408 43120 7688
rect 800 7008 43200 7408
rect 880 6728 43120 7008
rect 800 6328 43200 6728
rect 800 6048 43120 6328
rect 800 5648 43200 6048
rect 880 5368 43120 5648
rect 800 4968 43200 5368
rect 880 4688 43200 4968
rect 800 4288 43200 4688
rect 880 4008 43120 4288
rect 800 3608 43200 4008
rect 880 3328 43120 3608
rect 800 2928 43200 3328
rect 800 2648 43120 2928
rect 800 2248 43200 2648
rect 880 1968 43120 2248
rect 800 1568 43200 1968
rect 880 1288 43200 1568
rect 800 888 43200 1288
rect 880 608 43120 888
rect 800 208 43200 608
rect 800 35 43120 208
<< metal4 >>
rect 4208 2128 4528 41392
rect 19568 2128 19888 41392
rect 34928 2128 35248 41392
<< labels >>
rlabel metal3 s 0 40808 800 40928 6 active
port 1 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 24490 43200 24546 44000 6 io_in[10]
port 3 nsew signal input
rlabel metal2 s 18 43200 74 44000 6 io_in[11]
port 4 nsew signal input
rlabel metal3 s 43200 36728 44000 36848 6 io_in[12]
port 5 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 io_in[13]
port 6 nsew signal input
rlabel metal2 s 16762 43200 16818 44000 6 io_in[14]
port 7 nsew signal input
rlabel metal3 s 43200 38768 44000 38888 6 io_in[15]
port 8 nsew signal input
rlabel metal3 s 43200 3408 44000 3528 6 io_in[16]
port 9 nsew signal input
rlabel metal2 s 9034 43200 9090 44000 6 io_in[17]
port 10 nsew signal input
rlabel metal2 s 10966 43200 11022 44000 6 io_in[18]
port 11 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 io_in[19]
port 12 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 io_in[1]
port 13 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 io_in[20]
port 14 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 io_in[21]
port 15 nsew signal input
rlabel metal3 s 43200 13608 44000 13728 6 io_in[22]
port 16 nsew signal input
rlabel metal2 s 8390 43200 8446 44000 6 io_in[23]
port 17 nsew signal input
rlabel metal2 s 5814 43200 5870 44000 6 io_in[24]
port 18 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 io_in[25]
port 19 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 io_in[26]
port 20 nsew signal input
rlabel metal3 s 43200 9528 44000 9648 6 io_in[27]
port 21 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 io_in[28]
port 22 nsew signal input
rlabel metal2 s 43810 43200 43866 44000 6 io_in[29]
port 23 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 io_in[2]
port 24 nsew signal input
rlabel metal3 s 43200 17008 44000 17128 6 io_in[30]
port 25 nsew signal input
rlabel metal3 s 0 39448 800 39568 6 io_in[31]
port 26 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 io_in[32]
port 27 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 io_in[33]
port 28 nsew signal input
rlabel metal2 s 33506 43200 33562 44000 6 io_in[34]
port 29 nsew signal input
rlabel metal2 s 38658 43200 38714 44000 6 io_in[35]
port 30 nsew signal input
rlabel metal3 s 43200 27208 44000 27328 6 io_in[36]
port 31 nsew signal input
rlabel metal2 s 39302 43200 39358 44000 6 io_in[37]
port 32 nsew signal input
rlabel metal2 s 25134 43200 25190 44000 6 io_in[3]
port 33 nsew signal input
rlabel metal3 s 43200 26528 44000 26648 6 io_in[4]
port 34 nsew signal input
rlabel metal3 s 43200 42168 44000 42288 6 io_in[5]
port 35 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 io_in[6]
port 36 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 io_in[7]
port 37 nsew signal input
rlabel metal3 s 43200 29248 44000 29368 6 io_in[8]
port 38 nsew signal input
rlabel metal2 s 7746 43200 7802 44000 6 io_in[9]
port 39 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 io_oeb[0]
port 40 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 io_oeb[10]
port 41 nsew signal output
rlabel metal3 s 43200 25168 44000 25288 6 io_oeb[11]
port 42 nsew signal output
rlabel metal3 s 43200 12928 44000 13048 6 io_oeb[12]
port 43 nsew signal output
rlabel metal3 s 43200 12248 44000 12368 6 io_oeb[13]
port 44 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 io_oeb[14]
port 45 nsew signal output
rlabel metal2 s 12254 43200 12310 44000 6 io_oeb[15]
port 46 nsew signal output
rlabel metal3 s 43200 2048 44000 2168 6 io_oeb[16]
port 47 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 io_oeb[17]
port 48 nsew signal output
rlabel metal2 s 32218 43200 32274 44000 6 io_oeb[18]
port 49 nsew signal output
rlabel metal2 s 12898 43200 12954 44000 6 io_oeb[19]
port 50 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 io_oeb[1]
port 51 nsew signal output
rlabel metal3 s 43200 19048 44000 19168 6 io_oeb[20]
port 52 nsew signal output
rlabel metal2 s 1950 43200 2006 44000 6 io_oeb[21]
port 53 nsew signal output
rlabel metal2 s 4526 0 4582 800 6 io_oeb[22]
port 54 nsew signal output
rlabel metal2 s 21914 43200 21970 44000 6 io_oeb[23]
port 55 nsew signal output
rlabel metal2 s 23202 43200 23258 44000 6 io_oeb[24]
port 56 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 io_oeb[25]
port 57 nsew signal output
rlabel metal3 s 43200 34688 44000 34808 6 io_oeb[26]
port 58 nsew signal output
rlabel metal2 s 26422 43200 26478 44000 6 io_oeb[27]
port 59 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 io_oeb[28]
port 60 nsew signal output
rlabel metal3 s 43200 28568 44000 28688 6 io_oeb[29]
port 61 nsew signal output
rlabel metal2 s 36726 43200 36782 44000 6 io_oeb[2]
port 62 nsew signal output
rlabel metal2 s 2594 43200 2650 44000 6 io_oeb[30]
port 63 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 io_oeb[31]
port 64 nsew signal output
rlabel metal3 s 0 21768 800 21888 6 io_oeb[32]
port 65 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 io_oeb[33]
port 66 nsew signal output
rlabel metal2 s 9678 43200 9734 44000 6 io_oeb[34]
port 67 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 io_oeb[35]
port 68 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 io_oeb[36]
port 69 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 io_oeb[37]
port 70 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 io_oeb[3]
port 71 nsew signal output
rlabel metal3 s 43200 8 44000 128 6 io_oeb[4]
port 72 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 io_oeb[5]
port 73 nsew signal output
rlabel metal3 s 43200 15648 44000 15768 6 io_oeb[6]
port 74 nsew signal output
rlabel metal2 s 11610 43200 11666 44000 6 io_oeb[7]
port 75 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 io_oeb[8]
port 76 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 io_oeb[9]
port 77 nsew signal output
rlabel metal3 s 43200 41488 44000 41608 6 io_out[0]
port 78 nsew signal output
rlabel metal3 s 43200 23808 44000 23928 6 io_out[10]
port 79 nsew signal output
rlabel metal3 s 0 2048 800 2168 6 io_out[11]
port 80 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 io_out[12]
port 81 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 io_out[13]
port 82 nsew signal output
rlabel metal3 s 43200 35368 44000 35488 6 io_out[14]
port 83 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 io_out[15]
port 84 nsew signal output
rlabel metal3 s 43200 23128 44000 23248 6 io_out[16]
port 85 nsew signal output
rlabel metal2 s 40590 43200 40646 44000 6 io_out[17]
port 86 nsew signal output
rlabel metal2 s 41234 0 41290 800 6 io_out[18]
port 87 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 io_out[19]
port 88 nsew signal output
rlabel metal2 s 29642 43200 29698 44000 6 io_out[1]
port 89 nsew signal output
rlabel metal2 s 36082 43200 36138 44000 6 io_out[20]
port 90 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 io_out[21]
port 91 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 io_out[22]
port 92 nsew signal output
rlabel metal3 s 43200 19728 44000 19848 6 io_out[23]
port 93 nsew signal output
rlabel metal2 s 23846 0 23902 800 6 io_out[24]
port 94 nsew signal output
rlabel metal2 s 32862 43200 32918 44000 6 io_out[25]
port 95 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 io_out[26]
port 96 nsew signal output
rlabel metal2 s 34150 43200 34206 44000 6 io_out[27]
port 97 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 io_out[28]
port 98 nsew signal output
rlabel metal3 s 43200 688 44000 808 6 io_out[29]
port 99 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 io_out[2]
port 100 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 io_out[30]
port 101 nsew signal output
rlabel metal3 s 0 12248 800 12368 6 io_out[31]
port 102 nsew signal output
rlabel metal3 s 0 41488 800 41608 6 io_out[32]
port 103 nsew signal output
rlabel metal3 s 43200 6128 44000 6248 6 io_out[33]
port 104 nsew signal output
rlabel metal3 s 43200 36048 44000 36168 6 io_out[34]
port 105 nsew signal output
rlabel metal3 s 43200 33328 44000 33448 6 io_out[35]
port 106 nsew signal output
rlabel metal2 s 14186 43200 14242 44000 6 io_out[36]
port 107 nsew signal output
rlabel metal3 s 43200 39448 44000 39568 6 io_out[37]
port 108 nsew signal output
rlabel metal3 s 0 38088 800 38208 6 io_out[3]
port 109 nsew signal output
rlabel metal3 s 43200 25848 44000 25968 6 io_out[4]
port 110 nsew signal output
rlabel metal2 s 20626 43200 20682 44000 6 io_out[5]
port 111 nsew signal output
rlabel metal2 s 42522 43200 42578 44000 6 io_out[6]
port 112 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 io_out[7]
port 113 nsew signal output
rlabel metal2 s 16762 0 16818 800 6 io_out[8]
port 114 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 io_out[9]
port 115 nsew signal output
rlabel metal3 s 43200 6808 44000 6928 6 la1_data_in[0]
port 116 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 la1_data_in[10]
port 117 nsew signal input
rlabel metal3 s 43200 5448 44000 5568 6 la1_data_in[11]
port 118 nsew signal input
rlabel metal3 s 0 33328 800 33448 6 la1_data_in[12]
port 119 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 la1_data_in[13]
port 120 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 la1_data_in[14]
port 121 nsew signal input
rlabel metal2 s 14830 43200 14886 44000 6 la1_data_in[15]
port 122 nsew signal input
rlabel metal2 s 27710 43200 27766 44000 6 la1_data_in[16]
port 123 nsew signal input
rlabel metal2 s 21270 43200 21326 44000 6 la1_data_in[17]
port 124 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 la1_data_in[18]
port 125 nsew signal input
rlabel metal2 s 15474 43200 15530 44000 6 la1_data_in[19]
port 126 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 la1_data_in[1]
port 127 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 la1_data_in[20]
port 128 nsew signal input
rlabel metal2 s 43166 43200 43222 44000 6 la1_data_in[21]
port 129 nsew signal input
rlabel metal3 s 43200 7488 44000 7608 6 la1_data_in[22]
port 130 nsew signal input
rlabel metal3 s 0 688 800 808 6 la1_data_in[23]
port 131 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 la1_data_in[24]
port 132 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 la1_data_in[25]
port 133 nsew signal input
rlabel metal3 s 43200 2728 44000 2848 6 la1_data_in[26]
port 134 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 la1_data_in[27]
port 135 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 la1_data_in[28]
port 136 nsew signal input
rlabel metal2 s 662 43200 718 44000 6 la1_data_in[29]
port 137 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 la1_data_in[2]
port 138 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 la1_data_in[30]
port 139 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 la1_data_in[31]
port 140 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 la1_data_in[3]
port 141 nsew signal input
rlabel metal2 s 37370 43200 37426 44000 6 la1_data_in[4]
port 142 nsew signal input
rlabel metal3 s 43200 21768 44000 21888 6 la1_data_in[5]
port 143 nsew signal input
rlabel metal2 s 17406 43200 17462 44000 6 la1_data_in[6]
port 144 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 la1_data_in[7]
port 145 nsew signal input
rlabel metal2 s 18050 43200 18106 44000 6 la1_data_in[8]
port 146 nsew signal input
rlabel metal3 s 0 30608 800 30728 6 la1_data_in[9]
port 147 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 la1_data_out[0]
port 148 nsew signal output
rlabel metal3 s 43200 10208 44000 10328 6 la1_data_out[10]
port 149 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 la1_data_out[11]
port 150 nsew signal output
rlabel metal3 s 43200 40128 44000 40248 6 la1_data_out[12]
port 151 nsew signal output
rlabel metal2 s 4526 43200 4582 44000 6 la1_data_out[13]
port 152 nsew signal output
rlabel metal2 s 23846 43200 23902 44000 6 la1_data_out[14]
port 153 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 la1_data_out[15]
port 154 nsew signal output
rlabel metal3 s 43200 14968 44000 15088 6 la1_data_out[16]
port 155 nsew signal output
rlabel metal3 s 43200 31968 44000 32088 6 la1_data_out[17]
port 156 nsew signal output
rlabel metal2 s 5170 43200 5226 44000 6 la1_data_out[18]
port 157 nsew signal output
rlabel metal3 s 43200 22448 44000 22568 6 la1_data_out[19]
port 158 nsew signal output
rlabel metal3 s 0 40128 800 40248 6 la1_data_out[1]
port 159 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 la1_data_out[20]
port 160 nsew signal output
rlabel metal3 s 43200 38088 44000 38208 6 la1_data_out[21]
port 161 nsew signal output
rlabel metal2 s 27066 43200 27122 44000 6 la1_data_out[22]
port 162 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 la1_data_out[23]
port 163 nsew signal output
rlabel metal3 s 43200 16328 44000 16448 6 la1_data_out[24]
port 164 nsew signal output
rlabel metal3 s 0 3408 800 3528 6 la1_data_out[25]
port 165 nsew signal output
rlabel metal3 s 43200 4088 44000 4208 6 la1_data_out[26]
port 166 nsew signal output
rlabel metal3 s 0 42848 800 42968 6 la1_data_out[27]
port 167 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 la1_data_out[28]
port 168 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 la1_data_out[29]
port 169 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 la1_data_out[2]
port 170 nsew signal output
rlabel metal3 s 43200 10888 44000 11008 6 la1_data_out[30]
port 171 nsew signal output
rlabel metal3 s 43200 42848 44000 42968 6 la1_data_out[31]
port 172 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 la1_data_out[3]
port 173 nsew signal output
rlabel metal2 s 40590 0 40646 800 6 la1_data_out[4]
port 174 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 la1_data_out[5]
port 175 nsew signal output
rlabel metal3 s 43200 18368 44000 18488 6 la1_data_out[6]
port 176 nsew signal output
rlabel metal2 s 662 0 718 800 6 la1_data_out[7]
port 177 nsew signal output
rlabel metal3 s 43200 32648 44000 32768 6 la1_data_out[8]
port 178 nsew signal output
rlabel metal2 s 41878 43200 41934 44000 6 la1_data_out[9]
port 179 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 la1_oenb[0]
port 180 nsew signal input
rlabel metal2 s 39946 43200 40002 44000 6 la1_oenb[10]
port 181 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 la1_oenb[11]
port 182 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 la1_oenb[12]
port 183 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 la1_oenb[13]
port 184 nsew signal input
rlabel metal2 s 18 0 74 800 6 la1_oenb[14]
port 185 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 la1_oenb[15]
port 186 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 la1_oenb[16]
port 187 nsew signal input
rlabel metal2 s 3238 43200 3294 44000 6 la1_oenb[17]
port 188 nsew signal input
rlabel metal2 s 19982 43200 20038 44000 6 la1_oenb[18]
port 189 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 la1_oenb[19]
port 190 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 la1_oenb[1]
port 191 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 la1_oenb[20]
port 192 nsew signal input
rlabel metal2 s 28354 43200 28410 44000 6 la1_oenb[21]
port 193 nsew signal input
rlabel metal2 s 18694 43200 18750 44000 6 la1_oenb[22]
port 194 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 la1_oenb[23]
port 195 nsew signal input
rlabel metal2 s 35438 43200 35494 44000 6 la1_oenb[24]
port 196 nsew signal input
rlabel metal3 s 43200 8848 44000 8968 6 la1_oenb[25]
port 197 nsew signal input
rlabel metal3 s 0 34688 800 34808 6 la1_oenb[26]
port 198 nsew signal input
rlabel metal3 s 43200 31288 44000 31408 6 la1_oenb[27]
port 199 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 la1_oenb[28]
port 200 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 la1_oenb[29]
port 201 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 la1_oenb[2]
port 202 nsew signal input
rlabel metal3 s 43200 29928 44000 30048 6 la1_oenb[30]
port 203 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 la1_oenb[31]
port 204 nsew signal input
rlabel metal2 s 30930 43200 30986 44000 6 la1_oenb[3]
port 205 nsew signal input
rlabel metal2 s 30286 43200 30342 44000 6 la1_oenb[4]
port 206 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 la1_oenb[5]
port 207 nsew signal input
rlabel metal2 s 6458 43200 6514 44000 6 la1_oenb[6]
port 208 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 la1_oenb[7]
port 209 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 la1_oenb[8]
port 210 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 la1_oenb[9]
port 211 nsew signal input
rlabel metal4 s 4208 2128 4528 41392 6 vccd1
port 212 nsew power input
rlabel metal4 s 34928 2128 35248 41392 6 vccd1
port 212 nsew power input
rlabel metal4 s 19568 2128 19888 41392 6 vssd1
port 213 nsew ground input
rlabel metal3 s 43200 20408 44000 20528 6 wb_clk_i
port 214 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 44000 44000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3284258
string GDS_FILE /openlane/designs/wrapped_vga_clock/runs/RUN_2022.03.16_16.30.12/results/finishing/wrapped_vga_clock.magic.gds
string GDS_START 518106
<< end >>

